magic
tech sky130A
magscale 1 2
timestamp 1669319831
<< nwell >>
rect 14932 41259 42638 41492
rect 14932 39846 42639 41259
rect 15029 39845 42639 39846
rect 14050 33739 41756 33972
rect 14050 32326 41757 33739
rect 14147 32325 41757 32326
rect 5916 29979 33622 30212
rect 33944 29979 36918 30212
rect 5916 28566 33623 29979
rect 33944 28566 36919 29979
rect 6013 28565 33623 28566
rect 34041 28565 36919 28566
rect 9444 26219 15166 26452
rect 9444 24806 15167 26219
rect 9541 24805 15167 24806
rect 7582 22459 13304 22692
rect 7582 21046 13305 22459
rect 7679 21045 13305 21046
rect 23850 18699 26824 18932
rect 23850 17286 26825 18699
rect 23947 17285 26825 17286
<< pwell >>
rect 5958 40126 6526 40978
rect 5898 39606 5990 39778
rect 30024 37249 39404 37402
rect 28302 36366 28870 37218
rect 30024 36215 30177 37249
rect 31211 36215 31517 37249
rect 32551 36215 32857 37249
rect 33891 36215 34197 37249
rect 35231 36215 35537 37249
rect 36571 36215 36877 37249
rect 37911 36215 38217 37249
rect 39251 36215 39404 37249
rect 40632 36556 41300 36788
rect 30024 36062 39404 36215
rect 28242 35846 28334 36018
rect 38280 29036 38948 29268
rect 41024 29036 41692 29268
rect 7606 25276 8274 25508
rect 28260 25969 38980 26122
rect 22942 25086 27174 25938
rect 28260 24935 28413 25969
rect 29447 24935 29753 25969
rect 30787 24935 31093 25969
rect 32127 24935 32433 25969
rect 33467 24935 33773 25969
rect 34807 24935 35113 25969
rect 36147 24935 36453 25969
rect 37487 24935 37793 25969
rect 38827 24935 38980 25969
rect 40632 25276 41300 25508
rect 28260 24782 38980 24935
rect 22882 24566 22974 24738
rect 23942 24566 24114 24668
rect 25242 24566 25414 24668
rect 21008 22209 22348 22362
rect 21008 21175 21161 22209
rect 22195 21175 22348 22209
rect 28260 22209 38980 22362
rect 22942 21326 27174 22178
rect 21008 21022 22348 21175
rect 28260 21175 28413 22209
rect 29447 21175 29753 22209
rect 30787 21175 31093 22209
rect 32127 21175 32433 22209
rect 33467 21175 33773 22209
rect 34807 21175 35113 22209
rect 36147 21175 36453 22209
rect 37487 21175 37793 22209
rect 38827 21175 38980 22209
rect 40632 21516 41300 21748
rect 28260 21022 38980 21175
rect 22882 20806 22974 20978
rect 23942 20806 24114 20908
rect 25242 20806 25414 20908
rect 5988 17566 10220 18418
rect 11526 17756 12194 17988
rect 14270 17756 14938 17988
rect 28260 18449 38980 18602
rect 28260 17415 28413 18449
rect 29447 17415 29753 18449
rect 30787 17415 31093 18449
rect 32127 17415 32433 18449
rect 33467 17415 33773 18449
rect 34807 17415 35113 18449
rect 36147 17415 36453 18449
rect 37487 17415 37793 18449
rect 38827 17415 38980 18449
rect 40142 17756 40810 17988
rect 28260 17262 38980 17415
rect 5928 17046 6020 17218
rect 6988 17046 7160 17148
rect 8288 17046 8460 17148
rect 28260 14689 38980 14842
rect 8782 13996 9450 14228
rect 11526 13996 12194 14228
rect 14270 13996 14938 14228
rect 24462 13996 25130 14228
rect 28260 13655 28413 14689
rect 29447 13655 29753 14689
rect 30787 13655 31093 14689
rect 32127 13655 32433 14689
rect 33467 13655 33773 14689
rect 34807 13655 35113 14689
rect 36147 13655 36453 14689
rect 37487 13655 37793 14689
rect 38827 13655 38980 14689
rect 40142 13996 40810 14228
rect 28260 13502 38980 13655
rect 8782 10236 9450 10468
rect 11526 10236 12194 10468
rect 14270 10236 14938 10468
rect 24750 10236 25418 10468
rect 27794 10236 28462 10468
rect 30538 10236 31206 10468
rect 33282 10236 33950 10468
rect 36026 10236 36694 10468
rect 38770 10236 39438 10468
rect 8782 6476 9450 6708
rect 15440 6476 16108 6708
rect 18484 6476 19152 6708
rect 21228 6476 21896 6708
rect 23972 6476 24640 6708
rect 26716 6476 27384 6708
rect 29460 6476 30128 6708
rect 32204 6476 32872 6708
rect 36026 6476 36694 6708
rect 38770 6476 39438 6708
<< nbase >>
rect 30177 36215 31211 37249
rect 31517 36215 32551 37249
rect 32857 36215 33891 37249
rect 34197 36215 35231 37249
rect 35537 36215 36571 37249
rect 36877 36215 37911 37249
rect 38217 36215 39251 37249
rect 28413 24935 29447 25969
rect 29753 24935 30787 25969
rect 31093 24935 32127 25969
rect 32433 24935 33467 25969
rect 33773 24935 34807 25969
rect 35113 24935 36147 25969
rect 36453 24935 37487 25969
rect 37793 24935 38827 25969
rect 21161 21175 22195 22209
rect 28413 21175 29447 22209
rect 29753 21175 30787 22209
rect 31093 21175 32127 22209
rect 32433 21175 33467 22209
rect 33773 21175 34807 22209
rect 35113 21175 36147 22209
rect 36453 21175 37487 22209
rect 37793 21175 38827 22209
rect 28413 17415 29447 18449
rect 29753 17415 30787 18449
rect 31093 17415 32127 18449
rect 32433 17415 33467 18449
rect 33773 17415 34807 18449
rect 35113 17415 36147 18449
rect 36453 17415 37487 18449
rect 37793 17415 38827 18449
rect 28413 13655 29447 14689
rect 29753 13655 30787 14689
rect 31093 13655 32127 14689
rect 32433 13655 33467 14689
rect 33773 13655 34807 14689
rect 35113 13655 36147 14689
rect 36453 13655 37487 14689
rect 37793 13655 38827 14689
<< pmoslvt >>
rect 15123 39907 15523 41197
rect 15581 39907 15981 41197
rect 16039 39907 16439 41197
rect 16497 39907 16897 41197
rect 16955 39907 17355 41197
rect 17413 39907 17813 41197
rect 17871 39907 18271 41197
rect 18329 39907 18729 41197
rect 18787 39907 19187 41197
rect 19245 39907 19645 41197
rect 19703 39907 20103 41197
rect 20161 39907 20561 41197
rect 20619 39907 21019 41197
rect 21077 39907 21477 41197
rect 21535 39907 21935 41197
rect 21993 39907 22393 41197
rect 22451 39907 22851 41197
rect 22909 39907 23309 41197
rect 23367 39907 23767 41197
rect 23825 39907 24225 41197
rect 24283 39907 24683 41197
rect 24741 39907 25141 41197
rect 25199 39907 25599 41197
rect 25657 39907 26057 41197
rect 26115 39907 26515 41197
rect 26573 39907 26973 41197
rect 27031 39907 27431 41197
rect 27489 39907 27889 41197
rect 27947 39907 28347 41197
rect 28405 39907 28805 41197
rect 28863 39907 29263 41197
rect 29321 39907 29721 41197
rect 29779 39907 30179 41197
rect 30237 39907 30637 41197
rect 30695 39907 31095 41197
rect 31153 39907 31553 41197
rect 31611 39907 32011 41197
rect 32069 39907 32469 41197
rect 32527 39907 32927 41197
rect 32985 39907 33385 41197
rect 33443 39907 33843 41197
rect 33901 39907 34301 41197
rect 34359 39907 34759 41197
rect 34817 39907 35217 41197
rect 35275 39907 35675 41197
rect 35733 39907 36133 41197
rect 36191 39907 36591 41197
rect 36649 39907 37049 41197
rect 37107 39907 37507 41197
rect 37565 39907 37965 41197
rect 38023 39907 38423 41197
rect 38481 39907 38881 41197
rect 38939 39907 39339 41197
rect 39397 39907 39797 41197
rect 39855 39907 40255 41197
rect 40313 39907 40713 41197
rect 40771 39907 41171 41197
rect 41229 39907 41629 41197
rect 41687 39907 42087 41197
rect 42145 39907 42545 41197
rect 14241 32387 14641 33677
rect 14699 32387 15099 33677
rect 15157 32387 15557 33677
rect 15615 32387 16015 33677
rect 16073 32387 16473 33677
rect 16531 32387 16931 33677
rect 16989 32387 17389 33677
rect 17447 32387 17847 33677
rect 17905 32387 18305 33677
rect 18363 32387 18763 33677
rect 18821 32387 19221 33677
rect 19279 32387 19679 33677
rect 19737 32387 20137 33677
rect 20195 32387 20595 33677
rect 20653 32387 21053 33677
rect 21111 32387 21511 33677
rect 21569 32387 21969 33677
rect 22027 32387 22427 33677
rect 22485 32387 22885 33677
rect 22943 32387 23343 33677
rect 23401 32387 23801 33677
rect 23859 32387 24259 33677
rect 24317 32387 24717 33677
rect 24775 32387 25175 33677
rect 25233 32387 25633 33677
rect 25691 32387 26091 33677
rect 26149 32387 26549 33677
rect 26607 32387 27007 33677
rect 27065 32387 27465 33677
rect 27523 32387 27923 33677
rect 27981 32387 28381 33677
rect 28439 32387 28839 33677
rect 28897 32387 29297 33677
rect 29355 32387 29755 33677
rect 29813 32387 30213 33677
rect 30271 32387 30671 33677
rect 30729 32387 31129 33677
rect 31187 32387 31587 33677
rect 31645 32387 32045 33677
rect 32103 32387 32503 33677
rect 32561 32387 32961 33677
rect 33019 32387 33419 33677
rect 33477 32387 33877 33677
rect 33935 32387 34335 33677
rect 34393 32387 34793 33677
rect 34851 32387 35251 33677
rect 35309 32387 35709 33677
rect 35767 32387 36167 33677
rect 36225 32387 36625 33677
rect 36683 32387 37083 33677
rect 37141 32387 37541 33677
rect 37599 32387 37999 33677
rect 38057 32387 38457 33677
rect 38515 32387 38915 33677
rect 38973 32387 39373 33677
rect 39431 32387 39831 33677
rect 39889 32387 40289 33677
rect 40347 32387 40747 33677
rect 40805 32387 41205 33677
rect 41263 32387 41663 33677
rect 6107 28627 6507 29917
rect 6565 28627 6965 29917
rect 7023 28627 7423 29917
rect 7481 28627 7881 29917
rect 7939 28627 8339 29917
rect 8397 28627 8797 29917
rect 8855 28627 9255 29917
rect 9313 28627 9713 29917
rect 9771 28627 10171 29917
rect 10229 28627 10629 29917
rect 10687 28627 11087 29917
rect 11145 28627 11545 29917
rect 11603 28627 12003 29917
rect 12061 28627 12461 29917
rect 12519 28627 12919 29917
rect 12977 28627 13377 29917
rect 13435 28627 13835 29917
rect 13893 28627 14293 29917
rect 14351 28627 14751 29917
rect 14809 28627 15209 29917
rect 15267 28627 15667 29917
rect 15725 28627 16125 29917
rect 16183 28627 16583 29917
rect 16641 28627 17041 29917
rect 17099 28627 17499 29917
rect 17557 28627 17957 29917
rect 18015 28627 18415 29917
rect 18473 28627 18873 29917
rect 18931 28627 19331 29917
rect 19389 28627 19789 29917
rect 19847 28627 20247 29917
rect 20305 28627 20705 29917
rect 20763 28627 21163 29917
rect 21221 28627 21621 29917
rect 21679 28627 22079 29917
rect 22137 28627 22537 29917
rect 22595 28627 22995 29917
rect 23053 28627 23453 29917
rect 23511 28627 23911 29917
rect 23969 28627 24369 29917
rect 24427 28627 24827 29917
rect 24885 28627 25285 29917
rect 25343 28627 25743 29917
rect 25801 28627 26201 29917
rect 26259 28627 26659 29917
rect 26717 28627 27117 29917
rect 27175 28627 27575 29917
rect 27633 28627 28033 29917
rect 28091 28627 28491 29917
rect 28549 28627 28949 29917
rect 29007 28627 29407 29917
rect 29465 28627 29865 29917
rect 29923 28627 30323 29917
rect 30381 28627 30781 29917
rect 30839 28627 31239 29917
rect 31297 28627 31697 29917
rect 31755 28627 32155 29917
rect 32213 28627 32613 29917
rect 32671 28627 33071 29917
rect 33129 28627 33529 29917
rect 34135 28627 34535 29917
rect 34593 28627 34993 29917
rect 35051 28627 35451 29917
rect 35509 28627 35909 29917
rect 35967 28627 36367 29917
rect 36425 28627 36825 29917
rect 9635 24867 10035 26157
rect 10093 24867 10493 26157
rect 10551 24867 10951 26157
rect 11009 24867 11409 26157
rect 11467 24867 11867 26157
rect 11925 24867 12325 26157
rect 12383 24867 12783 26157
rect 12841 24867 13241 26157
rect 13299 24867 13699 26157
rect 13757 24867 14157 26157
rect 14215 24867 14615 26157
rect 14673 24867 15073 26157
rect 7773 21107 8173 22397
rect 8231 21107 8631 22397
rect 8689 21107 9089 22397
rect 9147 21107 9547 22397
rect 9605 21107 10005 22397
rect 10063 21107 10463 22397
rect 10521 21107 10921 22397
rect 10979 21107 11379 22397
rect 11437 21107 11837 22397
rect 11895 21107 12295 22397
rect 12353 21107 12753 22397
rect 12811 21107 13211 22397
rect 24041 17347 24441 18637
rect 24499 17347 24899 18637
rect 24957 17347 25357 18637
rect 25415 17347 25815 18637
rect 25873 17347 26273 18637
rect 26331 17347 26731 18637
<< nmoslvt >>
rect 6042 40152 6442 40952
rect 28386 36392 28786 37192
rect 23026 25112 23426 25912
rect 23484 25112 23884 25912
rect 23942 25112 24342 25912
rect 24400 25112 24800 25912
rect 24858 25112 25258 25912
rect 25316 25112 25716 25912
rect 25774 25112 26174 25912
rect 26232 25112 26632 25912
rect 26690 25112 27090 25912
rect 23026 21352 23426 22152
rect 23484 21352 23884 22152
rect 23942 21352 24342 22152
rect 24400 21352 24800 22152
rect 24858 21352 25258 22152
rect 25316 21352 25716 22152
rect 25774 21352 26174 22152
rect 26232 21352 26632 22152
rect 26690 21352 27090 22152
rect 6072 17592 6472 18392
rect 6530 17592 6930 18392
rect 6988 17592 7388 18392
rect 7446 17592 7846 18392
rect 7904 17592 8304 18392
rect 8362 17592 8762 18392
rect 8820 17592 9220 18392
rect 9278 17592 9678 18392
rect 9736 17592 10136 18392
<< ndiff >>
rect 5984 40909 6042 40952
rect 5984 40875 5996 40909
rect 6030 40875 6042 40909
rect 5984 40841 6042 40875
rect 5984 40807 5996 40841
rect 6030 40807 6042 40841
rect 5984 40773 6042 40807
rect 5984 40739 5996 40773
rect 6030 40739 6042 40773
rect 5984 40705 6042 40739
rect 5984 40671 5996 40705
rect 6030 40671 6042 40705
rect 5984 40637 6042 40671
rect 5984 40603 5996 40637
rect 6030 40603 6042 40637
rect 5984 40569 6042 40603
rect 5984 40535 5996 40569
rect 6030 40535 6042 40569
rect 5984 40501 6042 40535
rect 5984 40467 5996 40501
rect 6030 40467 6042 40501
rect 5984 40433 6042 40467
rect 5984 40399 5996 40433
rect 6030 40399 6042 40433
rect 5984 40365 6042 40399
rect 5984 40331 5996 40365
rect 6030 40331 6042 40365
rect 5984 40297 6042 40331
rect 5984 40263 5996 40297
rect 6030 40263 6042 40297
rect 5984 40229 6042 40263
rect 5984 40195 5996 40229
rect 6030 40195 6042 40229
rect 5984 40152 6042 40195
rect 6442 40909 6500 40952
rect 6442 40875 6454 40909
rect 6488 40875 6500 40909
rect 6442 40841 6500 40875
rect 6442 40807 6454 40841
rect 6488 40807 6500 40841
rect 6442 40773 6500 40807
rect 6442 40739 6454 40773
rect 6488 40739 6500 40773
rect 6442 40705 6500 40739
rect 6442 40671 6454 40705
rect 6488 40671 6500 40705
rect 6442 40637 6500 40671
rect 6442 40603 6454 40637
rect 6488 40603 6500 40637
rect 6442 40569 6500 40603
rect 6442 40535 6454 40569
rect 6488 40535 6500 40569
rect 6442 40501 6500 40535
rect 6442 40467 6454 40501
rect 6488 40467 6500 40501
rect 6442 40433 6500 40467
rect 6442 40399 6454 40433
rect 6488 40399 6500 40433
rect 6442 40365 6500 40399
rect 6442 40331 6454 40365
rect 6488 40331 6500 40365
rect 6442 40297 6500 40331
rect 6442 40263 6454 40297
rect 6488 40263 6500 40297
rect 6442 40229 6500 40263
rect 6442 40195 6454 40229
rect 6488 40195 6500 40229
rect 6442 40152 6500 40195
rect 28328 37149 28386 37192
rect 28328 37115 28340 37149
rect 28374 37115 28386 37149
rect 28328 37081 28386 37115
rect 28328 37047 28340 37081
rect 28374 37047 28386 37081
rect 28328 37013 28386 37047
rect 28328 36979 28340 37013
rect 28374 36979 28386 37013
rect 28328 36945 28386 36979
rect 28328 36911 28340 36945
rect 28374 36911 28386 36945
rect 28328 36877 28386 36911
rect 28328 36843 28340 36877
rect 28374 36843 28386 36877
rect 28328 36809 28386 36843
rect 28328 36775 28340 36809
rect 28374 36775 28386 36809
rect 28328 36741 28386 36775
rect 28328 36707 28340 36741
rect 28374 36707 28386 36741
rect 28328 36673 28386 36707
rect 28328 36639 28340 36673
rect 28374 36639 28386 36673
rect 28328 36605 28386 36639
rect 28328 36571 28340 36605
rect 28374 36571 28386 36605
rect 28328 36537 28386 36571
rect 28328 36503 28340 36537
rect 28374 36503 28386 36537
rect 28328 36469 28386 36503
rect 28328 36435 28340 36469
rect 28374 36435 28386 36469
rect 28328 36392 28386 36435
rect 28786 37149 28844 37192
rect 28786 37115 28798 37149
rect 28832 37115 28844 37149
rect 28786 37081 28844 37115
rect 28786 37047 28798 37081
rect 28832 37047 28844 37081
rect 28786 37013 28844 37047
rect 28786 36979 28798 37013
rect 28832 36979 28844 37013
rect 28786 36945 28844 36979
rect 28786 36911 28798 36945
rect 28832 36911 28844 36945
rect 28786 36877 28844 36911
rect 28786 36843 28798 36877
rect 28832 36843 28844 36877
rect 28786 36809 28844 36843
rect 28786 36775 28798 36809
rect 28832 36775 28844 36809
rect 28786 36741 28844 36775
rect 28786 36707 28798 36741
rect 28832 36707 28844 36741
rect 28786 36673 28844 36707
rect 28786 36639 28798 36673
rect 28832 36639 28844 36673
rect 28786 36605 28844 36639
rect 28786 36571 28798 36605
rect 28832 36571 28844 36605
rect 28786 36537 28844 36571
rect 28786 36503 28798 36537
rect 28832 36503 28844 36537
rect 28786 36469 28844 36503
rect 28786 36435 28798 36469
rect 28832 36435 28844 36469
rect 28786 36392 28844 36435
rect 22968 25869 23026 25912
rect 22968 25835 22980 25869
rect 23014 25835 23026 25869
rect 22968 25801 23026 25835
rect 22968 25767 22980 25801
rect 23014 25767 23026 25801
rect 22968 25733 23026 25767
rect 22968 25699 22980 25733
rect 23014 25699 23026 25733
rect 22968 25665 23026 25699
rect 22968 25631 22980 25665
rect 23014 25631 23026 25665
rect 22968 25597 23026 25631
rect 22968 25563 22980 25597
rect 23014 25563 23026 25597
rect 22968 25529 23026 25563
rect 22968 25495 22980 25529
rect 23014 25495 23026 25529
rect 22968 25461 23026 25495
rect 22968 25427 22980 25461
rect 23014 25427 23026 25461
rect 22968 25393 23026 25427
rect 22968 25359 22980 25393
rect 23014 25359 23026 25393
rect 22968 25325 23026 25359
rect 22968 25291 22980 25325
rect 23014 25291 23026 25325
rect 22968 25257 23026 25291
rect 22968 25223 22980 25257
rect 23014 25223 23026 25257
rect 22968 25189 23026 25223
rect 22968 25155 22980 25189
rect 23014 25155 23026 25189
rect 22968 25112 23026 25155
rect 23426 25869 23484 25912
rect 23426 25835 23438 25869
rect 23472 25835 23484 25869
rect 23426 25801 23484 25835
rect 23426 25767 23438 25801
rect 23472 25767 23484 25801
rect 23426 25733 23484 25767
rect 23426 25699 23438 25733
rect 23472 25699 23484 25733
rect 23426 25665 23484 25699
rect 23426 25631 23438 25665
rect 23472 25631 23484 25665
rect 23426 25597 23484 25631
rect 23426 25563 23438 25597
rect 23472 25563 23484 25597
rect 23426 25529 23484 25563
rect 23426 25495 23438 25529
rect 23472 25495 23484 25529
rect 23426 25461 23484 25495
rect 23426 25427 23438 25461
rect 23472 25427 23484 25461
rect 23426 25393 23484 25427
rect 23426 25359 23438 25393
rect 23472 25359 23484 25393
rect 23426 25325 23484 25359
rect 23426 25291 23438 25325
rect 23472 25291 23484 25325
rect 23426 25257 23484 25291
rect 23426 25223 23438 25257
rect 23472 25223 23484 25257
rect 23426 25189 23484 25223
rect 23426 25155 23438 25189
rect 23472 25155 23484 25189
rect 23426 25112 23484 25155
rect 23884 25869 23942 25912
rect 23884 25835 23896 25869
rect 23930 25835 23942 25869
rect 23884 25801 23942 25835
rect 23884 25767 23896 25801
rect 23930 25767 23942 25801
rect 23884 25733 23942 25767
rect 23884 25699 23896 25733
rect 23930 25699 23942 25733
rect 23884 25665 23942 25699
rect 23884 25631 23896 25665
rect 23930 25631 23942 25665
rect 23884 25597 23942 25631
rect 23884 25563 23896 25597
rect 23930 25563 23942 25597
rect 23884 25529 23942 25563
rect 23884 25495 23896 25529
rect 23930 25495 23942 25529
rect 23884 25461 23942 25495
rect 23884 25427 23896 25461
rect 23930 25427 23942 25461
rect 23884 25393 23942 25427
rect 23884 25359 23896 25393
rect 23930 25359 23942 25393
rect 23884 25325 23942 25359
rect 23884 25291 23896 25325
rect 23930 25291 23942 25325
rect 23884 25257 23942 25291
rect 23884 25223 23896 25257
rect 23930 25223 23942 25257
rect 23884 25189 23942 25223
rect 23884 25155 23896 25189
rect 23930 25155 23942 25189
rect 23884 25112 23942 25155
rect 24342 25869 24400 25912
rect 24342 25835 24354 25869
rect 24388 25835 24400 25869
rect 24342 25801 24400 25835
rect 24342 25767 24354 25801
rect 24388 25767 24400 25801
rect 24342 25733 24400 25767
rect 24342 25699 24354 25733
rect 24388 25699 24400 25733
rect 24342 25665 24400 25699
rect 24342 25631 24354 25665
rect 24388 25631 24400 25665
rect 24342 25597 24400 25631
rect 24342 25563 24354 25597
rect 24388 25563 24400 25597
rect 24342 25529 24400 25563
rect 24342 25495 24354 25529
rect 24388 25495 24400 25529
rect 24342 25461 24400 25495
rect 24342 25427 24354 25461
rect 24388 25427 24400 25461
rect 24342 25393 24400 25427
rect 24342 25359 24354 25393
rect 24388 25359 24400 25393
rect 24342 25325 24400 25359
rect 24342 25291 24354 25325
rect 24388 25291 24400 25325
rect 24342 25257 24400 25291
rect 24342 25223 24354 25257
rect 24388 25223 24400 25257
rect 24342 25189 24400 25223
rect 24342 25155 24354 25189
rect 24388 25155 24400 25189
rect 24342 25112 24400 25155
rect 24800 25869 24858 25912
rect 24800 25835 24812 25869
rect 24846 25835 24858 25869
rect 24800 25801 24858 25835
rect 24800 25767 24812 25801
rect 24846 25767 24858 25801
rect 24800 25733 24858 25767
rect 24800 25699 24812 25733
rect 24846 25699 24858 25733
rect 24800 25665 24858 25699
rect 24800 25631 24812 25665
rect 24846 25631 24858 25665
rect 24800 25597 24858 25631
rect 24800 25563 24812 25597
rect 24846 25563 24858 25597
rect 24800 25529 24858 25563
rect 24800 25495 24812 25529
rect 24846 25495 24858 25529
rect 24800 25461 24858 25495
rect 24800 25427 24812 25461
rect 24846 25427 24858 25461
rect 24800 25393 24858 25427
rect 24800 25359 24812 25393
rect 24846 25359 24858 25393
rect 24800 25325 24858 25359
rect 24800 25291 24812 25325
rect 24846 25291 24858 25325
rect 24800 25257 24858 25291
rect 24800 25223 24812 25257
rect 24846 25223 24858 25257
rect 24800 25189 24858 25223
rect 24800 25155 24812 25189
rect 24846 25155 24858 25189
rect 24800 25112 24858 25155
rect 25258 25869 25316 25912
rect 25258 25835 25270 25869
rect 25304 25835 25316 25869
rect 25258 25801 25316 25835
rect 25258 25767 25270 25801
rect 25304 25767 25316 25801
rect 25258 25733 25316 25767
rect 25258 25699 25270 25733
rect 25304 25699 25316 25733
rect 25258 25665 25316 25699
rect 25258 25631 25270 25665
rect 25304 25631 25316 25665
rect 25258 25597 25316 25631
rect 25258 25563 25270 25597
rect 25304 25563 25316 25597
rect 25258 25529 25316 25563
rect 25258 25495 25270 25529
rect 25304 25495 25316 25529
rect 25258 25461 25316 25495
rect 25258 25427 25270 25461
rect 25304 25427 25316 25461
rect 25258 25393 25316 25427
rect 25258 25359 25270 25393
rect 25304 25359 25316 25393
rect 25258 25325 25316 25359
rect 25258 25291 25270 25325
rect 25304 25291 25316 25325
rect 25258 25257 25316 25291
rect 25258 25223 25270 25257
rect 25304 25223 25316 25257
rect 25258 25189 25316 25223
rect 25258 25155 25270 25189
rect 25304 25155 25316 25189
rect 25258 25112 25316 25155
rect 25716 25869 25774 25912
rect 25716 25835 25728 25869
rect 25762 25835 25774 25869
rect 25716 25801 25774 25835
rect 25716 25767 25728 25801
rect 25762 25767 25774 25801
rect 25716 25733 25774 25767
rect 25716 25699 25728 25733
rect 25762 25699 25774 25733
rect 25716 25665 25774 25699
rect 25716 25631 25728 25665
rect 25762 25631 25774 25665
rect 25716 25597 25774 25631
rect 25716 25563 25728 25597
rect 25762 25563 25774 25597
rect 25716 25529 25774 25563
rect 25716 25495 25728 25529
rect 25762 25495 25774 25529
rect 25716 25461 25774 25495
rect 25716 25427 25728 25461
rect 25762 25427 25774 25461
rect 25716 25393 25774 25427
rect 25716 25359 25728 25393
rect 25762 25359 25774 25393
rect 25716 25325 25774 25359
rect 25716 25291 25728 25325
rect 25762 25291 25774 25325
rect 25716 25257 25774 25291
rect 25716 25223 25728 25257
rect 25762 25223 25774 25257
rect 25716 25189 25774 25223
rect 25716 25155 25728 25189
rect 25762 25155 25774 25189
rect 25716 25112 25774 25155
rect 26174 25869 26232 25912
rect 26174 25835 26186 25869
rect 26220 25835 26232 25869
rect 26174 25801 26232 25835
rect 26174 25767 26186 25801
rect 26220 25767 26232 25801
rect 26174 25733 26232 25767
rect 26174 25699 26186 25733
rect 26220 25699 26232 25733
rect 26174 25665 26232 25699
rect 26174 25631 26186 25665
rect 26220 25631 26232 25665
rect 26174 25597 26232 25631
rect 26174 25563 26186 25597
rect 26220 25563 26232 25597
rect 26174 25529 26232 25563
rect 26174 25495 26186 25529
rect 26220 25495 26232 25529
rect 26174 25461 26232 25495
rect 26174 25427 26186 25461
rect 26220 25427 26232 25461
rect 26174 25393 26232 25427
rect 26174 25359 26186 25393
rect 26220 25359 26232 25393
rect 26174 25325 26232 25359
rect 26174 25291 26186 25325
rect 26220 25291 26232 25325
rect 26174 25257 26232 25291
rect 26174 25223 26186 25257
rect 26220 25223 26232 25257
rect 26174 25189 26232 25223
rect 26174 25155 26186 25189
rect 26220 25155 26232 25189
rect 26174 25112 26232 25155
rect 26632 25869 26690 25912
rect 26632 25835 26644 25869
rect 26678 25835 26690 25869
rect 26632 25801 26690 25835
rect 26632 25767 26644 25801
rect 26678 25767 26690 25801
rect 26632 25733 26690 25767
rect 26632 25699 26644 25733
rect 26678 25699 26690 25733
rect 26632 25665 26690 25699
rect 26632 25631 26644 25665
rect 26678 25631 26690 25665
rect 26632 25597 26690 25631
rect 26632 25563 26644 25597
rect 26678 25563 26690 25597
rect 26632 25529 26690 25563
rect 26632 25495 26644 25529
rect 26678 25495 26690 25529
rect 26632 25461 26690 25495
rect 26632 25427 26644 25461
rect 26678 25427 26690 25461
rect 26632 25393 26690 25427
rect 26632 25359 26644 25393
rect 26678 25359 26690 25393
rect 26632 25325 26690 25359
rect 26632 25291 26644 25325
rect 26678 25291 26690 25325
rect 26632 25257 26690 25291
rect 26632 25223 26644 25257
rect 26678 25223 26690 25257
rect 26632 25189 26690 25223
rect 26632 25155 26644 25189
rect 26678 25155 26690 25189
rect 26632 25112 26690 25155
rect 27090 25869 27148 25912
rect 27090 25835 27102 25869
rect 27136 25835 27148 25869
rect 27090 25801 27148 25835
rect 27090 25767 27102 25801
rect 27136 25767 27148 25801
rect 27090 25733 27148 25767
rect 27090 25699 27102 25733
rect 27136 25699 27148 25733
rect 27090 25665 27148 25699
rect 27090 25631 27102 25665
rect 27136 25631 27148 25665
rect 27090 25597 27148 25631
rect 27090 25563 27102 25597
rect 27136 25563 27148 25597
rect 27090 25529 27148 25563
rect 27090 25495 27102 25529
rect 27136 25495 27148 25529
rect 27090 25461 27148 25495
rect 27090 25427 27102 25461
rect 27136 25427 27148 25461
rect 27090 25393 27148 25427
rect 27090 25359 27102 25393
rect 27136 25359 27148 25393
rect 27090 25325 27148 25359
rect 27090 25291 27102 25325
rect 27136 25291 27148 25325
rect 27090 25257 27148 25291
rect 27090 25223 27102 25257
rect 27136 25223 27148 25257
rect 27090 25189 27148 25223
rect 27090 25155 27102 25189
rect 27136 25155 27148 25189
rect 27090 25112 27148 25155
rect 22968 22109 23026 22152
rect 22968 22075 22980 22109
rect 23014 22075 23026 22109
rect 22968 22041 23026 22075
rect 22968 22007 22980 22041
rect 23014 22007 23026 22041
rect 22968 21973 23026 22007
rect 22968 21939 22980 21973
rect 23014 21939 23026 21973
rect 22968 21905 23026 21939
rect 22968 21871 22980 21905
rect 23014 21871 23026 21905
rect 22968 21837 23026 21871
rect 22968 21803 22980 21837
rect 23014 21803 23026 21837
rect 22968 21769 23026 21803
rect 22968 21735 22980 21769
rect 23014 21735 23026 21769
rect 22968 21701 23026 21735
rect 22968 21667 22980 21701
rect 23014 21667 23026 21701
rect 22968 21633 23026 21667
rect 22968 21599 22980 21633
rect 23014 21599 23026 21633
rect 22968 21565 23026 21599
rect 22968 21531 22980 21565
rect 23014 21531 23026 21565
rect 22968 21497 23026 21531
rect 22968 21463 22980 21497
rect 23014 21463 23026 21497
rect 22968 21429 23026 21463
rect 22968 21395 22980 21429
rect 23014 21395 23026 21429
rect 22968 21352 23026 21395
rect 23426 22109 23484 22152
rect 23426 22075 23438 22109
rect 23472 22075 23484 22109
rect 23426 22041 23484 22075
rect 23426 22007 23438 22041
rect 23472 22007 23484 22041
rect 23426 21973 23484 22007
rect 23426 21939 23438 21973
rect 23472 21939 23484 21973
rect 23426 21905 23484 21939
rect 23426 21871 23438 21905
rect 23472 21871 23484 21905
rect 23426 21837 23484 21871
rect 23426 21803 23438 21837
rect 23472 21803 23484 21837
rect 23426 21769 23484 21803
rect 23426 21735 23438 21769
rect 23472 21735 23484 21769
rect 23426 21701 23484 21735
rect 23426 21667 23438 21701
rect 23472 21667 23484 21701
rect 23426 21633 23484 21667
rect 23426 21599 23438 21633
rect 23472 21599 23484 21633
rect 23426 21565 23484 21599
rect 23426 21531 23438 21565
rect 23472 21531 23484 21565
rect 23426 21497 23484 21531
rect 23426 21463 23438 21497
rect 23472 21463 23484 21497
rect 23426 21429 23484 21463
rect 23426 21395 23438 21429
rect 23472 21395 23484 21429
rect 23426 21352 23484 21395
rect 23884 22109 23942 22152
rect 23884 22075 23896 22109
rect 23930 22075 23942 22109
rect 23884 22041 23942 22075
rect 23884 22007 23896 22041
rect 23930 22007 23942 22041
rect 23884 21973 23942 22007
rect 23884 21939 23896 21973
rect 23930 21939 23942 21973
rect 23884 21905 23942 21939
rect 23884 21871 23896 21905
rect 23930 21871 23942 21905
rect 23884 21837 23942 21871
rect 23884 21803 23896 21837
rect 23930 21803 23942 21837
rect 23884 21769 23942 21803
rect 23884 21735 23896 21769
rect 23930 21735 23942 21769
rect 23884 21701 23942 21735
rect 23884 21667 23896 21701
rect 23930 21667 23942 21701
rect 23884 21633 23942 21667
rect 23884 21599 23896 21633
rect 23930 21599 23942 21633
rect 23884 21565 23942 21599
rect 23884 21531 23896 21565
rect 23930 21531 23942 21565
rect 23884 21497 23942 21531
rect 23884 21463 23896 21497
rect 23930 21463 23942 21497
rect 23884 21429 23942 21463
rect 23884 21395 23896 21429
rect 23930 21395 23942 21429
rect 23884 21352 23942 21395
rect 24342 22109 24400 22152
rect 24342 22075 24354 22109
rect 24388 22075 24400 22109
rect 24342 22041 24400 22075
rect 24342 22007 24354 22041
rect 24388 22007 24400 22041
rect 24342 21973 24400 22007
rect 24342 21939 24354 21973
rect 24388 21939 24400 21973
rect 24342 21905 24400 21939
rect 24342 21871 24354 21905
rect 24388 21871 24400 21905
rect 24342 21837 24400 21871
rect 24342 21803 24354 21837
rect 24388 21803 24400 21837
rect 24342 21769 24400 21803
rect 24342 21735 24354 21769
rect 24388 21735 24400 21769
rect 24342 21701 24400 21735
rect 24342 21667 24354 21701
rect 24388 21667 24400 21701
rect 24342 21633 24400 21667
rect 24342 21599 24354 21633
rect 24388 21599 24400 21633
rect 24342 21565 24400 21599
rect 24342 21531 24354 21565
rect 24388 21531 24400 21565
rect 24342 21497 24400 21531
rect 24342 21463 24354 21497
rect 24388 21463 24400 21497
rect 24342 21429 24400 21463
rect 24342 21395 24354 21429
rect 24388 21395 24400 21429
rect 24342 21352 24400 21395
rect 24800 22109 24858 22152
rect 24800 22075 24812 22109
rect 24846 22075 24858 22109
rect 24800 22041 24858 22075
rect 24800 22007 24812 22041
rect 24846 22007 24858 22041
rect 24800 21973 24858 22007
rect 24800 21939 24812 21973
rect 24846 21939 24858 21973
rect 24800 21905 24858 21939
rect 24800 21871 24812 21905
rect 24846 21871 24858 21905
rect 24800 21837 24858 21871
rect 24800 21803 24812 21837
rect 24846 21803 24858 21837
rect 24800 21769 24858 21803
rect 24800 21735 24812 21769
rect 24846 21735 24858 21769
rect 24800 21701 24858 21735
rect 24800 21667 24812 21701
rect 24846 21667 24858 21701
rect 24800 21633 24858 21667
rect 24800 21599 24812 21633
rect 24846 21599 24858 21633
rect 24800 21565 24858 21599
rect 24800 21531 24812 21565
rect 24846 21531 24858 21565
rect 24800 21497 24858 21531
rect 24800 21463 24812 21497
rect 24846 21463 24858 21497
rect 24800 21429 24858 21463
rect 24800 21395 24812 21429
rect 24846 21395 24858 21429
rect 24800 21352 24858 21395
rect 25258 22109 25316 22152
rect 25258 22075 25270 22109
rect 25304 22075 25316 22109
rect 25258 22041 25316 22075
rect 25258 22007 25270 22041
rect 25304 22007 25316 22041
rect 25258 21973 25316 22007
rect 25258 21939 25270 21973
rect 25304 21939 25316 21973
rect 25258 21905 25316 21939
rect 25258 21871 25270 21905
rect 25304 21871 25316 21905
rect 25258 21837 25316 21871
rect 25258 21803 25270 21837
rect 25304 21803 25316 21837
rect 25258 21769 25316 21803
rect 25258 21735 25270 21769
rect 25304 21735 25316 21769
rect 25258 21701 25316 21735
rect 25258 21667 25270 21701
rect 25304 21667 25316 21701
rect 25258 21633 25316 21667
rect 25258 21599 25270 21633
rect 25304 21599 25316 21633
rect 25258 21565 25316 21599
rect 25258 21531 25270 21565
rect 25304 21531 25316 21565
rect 25258 21497 25316 21531
rect 25258 21463 25270 21497
rect 25304 21463 25316 21497
rect 25258 21429 25316 21463
rect 25258 21395 25270 21429
rect 25304 21395 25316 21429
rect 25258 21352 25316 21395
rect 25716 22109 25774 22152
rect 25716 22075 25728 22109
rect 25762 22075 25774 22109
rect 25716 22041 25774 22075
rect 25716 22007 25728 22041
rect 25762 22007 25774 22041
rect 25716 21973 25774 22007
rect 25716 21939 25728 21973
rect 25762 21939 25774 21973
rect 25716 21905 25774 21939
rect 25716 21871 25728 21905
rect 25762 21871 25774 21905
rect 25716 21837 25774 21871
rect 25716 21803 25728 21837
rect 25762 21803 25774 21837
rect 25716 21769 25774 21803
rect 25716 21735 25728 21769
rect 25762 21735 25774 21769
rect 25716 21701 25774 21735
rect 25716 21667 25728 21701
rect 25762 21667 25774 21701
rect 25716 21633 25774 21667
rect 25716 21599 25728 21633
rect 25762 21599 25774 21633
rect 25716 21565 25774 21599
rect 25716 21531 25728 21565
rect 25762 21531 25774 21565
rect 25716 21497 25774 21531
rect 25716 21463 25728 21497
rect 25762 21463 25774 21497
rect 25716 21429 25774 21463
rect 25716 21395 25728 21429
rect 25762 21395 25774 21429
rect 25716 21352 25774 21395
rect 26174 22109 26232 22152
rect 26174 22075 26186 22109
rect 26220 22075 26232 22109
rect 26174 22041 26232 22075
rect 26174 22007 26186 22041
rect 26220 22007 26232 22041
rect 26174 21973 26232 22007
rect 26174 21939 26186 21973
rect 26220 21939 26232 21973
rect 26174 21905 26232 21939
rect 26174 21871 26186 21905
rect 26220 21871 26232 21905
rect 26174 21837 26232 21871
rect 26174 21803 26186 21837
rect 26220 21803 26232 21837
rect 26174 21769 26232 21803
rect 26174 21735 26186 21769
rect 26220 21735 26232 21769
rect 26174 21701 26232 21735
rect 26174 21667 26186 21701
rect 26220 21667 26232 21701
rect 26174 21633 26232 21667
rect 26174 21599 26186 21633
rect 26220 21599 26232 21633
rect 26174 21565 26232 21599
rect 26174 21531 26186 21565
rect 26220 21531 26232 21565
rect 26174 21497 26232 21531
rect 26174 21463 26186 21497
rect 26220 21463 26232 21497
rect 26174 21429 26232 21463
rect 26174 21395 26186 21429
rect 26220 21395 26232 21429
rect 26174 21352 26232 21395
rect 26632 22109 26690 22152
rect 26632 22075 26644 22109
rect 26678 22075 26690 22109
rect 26632 22041 26690 22075
rect 26632 22007 26644 22041
rect 26678 22007 26690 22041
rect 26632 21973 26690 22007
rect 26632 21939 26644 21973
rect 26678 21939 26690 21973
rect 26632 21905 26690 21939
rect 26632 21871 26644 21905
rect 26678 21871 26690 21905
rect 26632 21837 26690 21871
rect 26632 21803 26644 21837
rect 26678 21803 26690 21837
rect 26632 21769 26690 21803
rect 26632 21735 26644 21769
rect 26678 21735 26690 21769
rect 26632 21701 26690 21735
rect 26632 21667 26644 21701
rect 26678 21667 26690 21701
rect 26632 21633 26690 21667
rect 26632 21599 26644 21633
rect 26678 21599 26690 21633
rect 26632 21565 26690 21599
rect 26632 21531 26644 21565
rect 26678 21531 26690 21565
rect 26632 21497 26690 21531
rect 26632 21463 26644 21497
rect 26678 21463 26690 21497
rect 26632 21429 26690 21463
rect 26632 21395 26644 21429
rect 26678 21395 26690 21429
rect 26632 21352 26690 21395
rect 27090 22109 27148 22152
rect 27090 22075 27102 22109
rect 27136 22075 27148 22109
rect 27090 22041 27148 22075
rect 27090 22007 27102 22041
rect 27136 22007 27148 22041
rect 27090 21973 27148 22007
rect 27090 21939 27102 21973
rect 27136 21939 27148 21973
rect 27090 21905 27148 21939
rect 27090 21871 27102 21905
rect 27136 21871 27148 21905
rect 27090 21837 27148 21871
rect 27090 21803 27102 21837
rect 27136 21803 27148 21837
rect 27090 21769 27148 21803
rect 27090 21735 27102 21769
rect 27136 21735 27148 21769
rect 27090 21701 27148 21735
rect 27090 21667 27102 21701
rect 27136 21667 27148 21701
rect 27090 21633 27148 21667
rect 27090 21599 27102 21633
rect 27136 21599 27148 21633
rect 27090 21565 27148 21599
rect 27090 21531 27102 21565
rect 27136 21531 27148 21565
rect 27090 21497 27148 21531
rect 27090 21463 27102 21497
rect 27136 21463 27148 21497
rect 27090 21429 27148 21463
rect 27090 21395 27102 21429
rect 27136 21395 27148 21429
rect 27090 21352 27148 21395
rect 6014 18349 6072 18392
rect 6014 18315 6026 18349
rect 6060 18315 6072 18349
rect 6014 18281 6072 18315
rect 6014 18247 6026 18281
rect 6060 18247 6072 18281
rect 6014 18213 6072 18247
rect 6014 18179 6026 18213
rect 6060 18179 6072 18213
rect 6014 18145 6072 18179
rect 6014 18111 6026 18145
rect 6060 18111 6072 18145
rect 6014 18077 6072 18111
rect 6014 18043 6026 18077
rect 6060 18043 6072 18077
rect 6014 18009 6072 18043
rect 6014 17975 6026 18009
rect 6060 17975 6072 18009
rect 6014 17941 6072 17975
rect 6014 17907 6026 17941
rect 6060 17907 6072 17941
rect 6014 17873 6072 17907
rect 6014 17839 6026 17873
rect 6060 17839 6072 17873
rect 6014 17805 6072 17839
rect 6014 17771 6026 17805
rect 6060 17771 6072 17805
rect 6014 17737 6072 17771
rect 6014 17703 6026 17737
rect 6060 17703 6072 17737
rect 6014 17669 6072 17703
rect 6014 17635 6026 17669
rect 6060 17635 6072 17669
rect 6014 17592 6072 17635
rect 6472 18349 6530 18392
rect 6472 18315 6484 18349
rect 6518 18315 6530 18349
rect 6472 18281 6530 18315
rect 6472 18247 6484 18281
rect 6518 18247 6530 18281
rect 6472 18213 6530 18247
rect 6472 18179 6484 18213
rect 6518 18179 6530 18213
rect 6472 18145 6530 18179
rect 6472 18111 6484 18145
rect 6518 18111 6530 18145
rect 6472 18077 6530 18111
rect 6472 18043 6484 18077
rect 6518 18043 6530 18077
rect 6472 18009 6530 18043
rect 6472 17975 6484 18009
rect 6518 17975 6530 18009
rect 6472 17941 6530 17975
rect 6472 17907 6484 17941
rect 6518 17907 6530 17941
rect 6472 17873 6530 17907
rect 6472 17839 6484 17873
rect 6518 17839 6530 17873
rect 6472 17805 6530 17839
rect 6472 17771 6484 17805
rect 6518 17771 6530 17805
rect 6472 17737 6530 17771
rect 6472 17703 6484 17737
rect 6518 17703 6530 17737
rect 6472 17669 6530 17703
rect 6472 17635 6484 17669
rect 6518 17635 6530 17669
rect 6472 17592 6530 17635
rect 6930 18349 6988 18392
rect 6930 18315 6942 18349
rect 6976 18315 6988 18349
rect 6930 18281 6988 18315
rect 6930 18247 6942 18281
rect 6976 18247 6988 18281
rect 6930 18213 6988 18247
rect 6930 18179 6942 18213
rect 6976 18179 6988 18213
rect 6930 18145 6988 18179
rect 6930 18111 6942 18145
rect 6976 18111 6988 18145
rect 6930 18077 6988 18111
rect 6930 18043 6942 18077
rect 6976 18043 6988 18077
rect 6930 18009 6988 18043
rect 6930 17975 6942 18009
rect 6976 17975 6988 18009
rect 6930 17941 6988 17975
rect 6930 17907 6942 17941
rect 6976 17907 6988 17941
rect 6930 17873 6988 17907
rect 6930 17839 6942 17873
rect 6976 17839 6988 17873
rect 6930 17805 6988 17839
rect 6930 17771 6942 17805
rect 6976 17771 6988 17805
rect 6930 17737 6988 17771
rect 6930 17703 6942 17737
rect 6976 17703 6988 17737
rect 6930 17669 6988 17703
rect 6930 17635 6942 17669
rect 6976 17635 6988 17669
rect 6930 17592 6988 17635
rect 7388 18349 7446 18392
rect 7388 18315 7400 18349
rect 7434 18315 7446 18349
rect 7388 18281 7446 18315
rect 7388 18247 7400 18281
rect 7434 18247 7446 18281
rect 7388 18213 7446 18247
rect 7388 18179 7400 18213
rect 7434 18179 7446 18213
rect 7388 18145 7446 18179
rect 7388 18111 7400 18145
rect 7434 18111 7446 18145
rect 7388 18077 7446 18111
rect 7388 18043 7400 18077
rect 7434 18043 7446 18077
rect 7388 18009 7446 18043
rect 7388 17975 7400 18009
rect 7434 17975 7446 18009
rect 7388 17941 7446 17975
rect 7388 17907 7400 17941
rect 7434 17907 7446 17941
rect 7388 17873 7446 17907
rect 7388 17839 7400 17873
rect 7434 17839 7446 17873
rect 7388 17805 7446 17839
rect 7388 17771 7400 17805
rect 7434 17771 7446 17805
rect 7388 17737 7446 17771
rect 7388 17703 7400 17737
rect 7434 17703 7446 17737
rect 7388 17669 7446 17703
rect 7388 17635 7400 17669
rect 7434 17635 7446 17669
rect 7388 17592 7446 17635
rect 7846 18349 7904 18392
rect 7846 18315 7858 18349
rect 7892 18315 7904 18349
rect 7846 18281 7904 18315
rect 7846 18247 7858 18281
rect 7892 18247 7904 18281
rect 7846 18213 7904 18247
rect 7846 18179 7858 18213
rect 7892 18179 7904 18213
rect 7846 18145 7904 18179
rect 7846 18111 7858 18145
rect 7892 18111 7904 18145
rect 7846 18077 7904 18111
rect 7846 18043 7858 18077
rect 7892 18043 7904 18077
rect 7846 18009 7904 18043
rect 7846 17975 7858 18009
rect 7892 17975 7904 18009
rect 7846 17941 7904 17975
rect 7846 17907 7858 17941
rect 7892 17907 7904 17941
rect 7846 17873 7904 17907
rect 7846 17839 7858 17873
rect 7892 17839 7904 17873
rect 7846 17805 7904 17839
rect 7846 17771 7858 17805
rect 7892 17771 7904 17805
rect 7846 17737 7904 17771
rect 7846 17703 7858 17737
rect 7892 17703 7904 17737
rect 7846 17669 7904 17703
rect 7846 17635 7858 17669
rect 7892 17635 7904 17669
rect 7846 17592 7904 17635
rect 8304 18349 8362 18392
rect 8304 18315 8316 18349
rect 8350 18315 8362 18349
rect 8304 18281 8362 18315
rect 8304 18247 8316 18281
rect 8350 18247 8362 18281
rect 8304 18213 8362 18247
rect 8304 18179 8316 18213
rect 8350 18179 8362 18213
rect 8304 18145 8362 18179
rect 8304 18111 8316 18145
rect 8350 18111 8362 18145
rect 8304 18077 8362 18111
rect 8304 18043 8316 18077
rect 8350 18043 8362 18077
rect 8304 18009 8362 18043
rect 8304 17975 8316 18009
rect 8350 17975 8362 18009
rect 8304 17941 8362 17975
rect 8304 17907 8316 17941
rect 8350 17907 8362 17941
rect 8304 17873 8362 17907
rect 8304 17839 8316 17873
rect 8350 17839 8362 17873
rect 8304 17805 8362 17839
rect 8304 17771 8316 17805
rect 8350 17771 8362 17805
rect 8304 17737 8362 17771
rect 8304 17703 8316 17737
rect 8350 17703 8362 17737
rect 8304 17669 8362 17703
rect 8304 17635 8316 17669
rect 8350 17635 8362 17669
rect 8304 17592 8362 17635
rect 8762 18349 8820 18392
rect 8762 18315 8774 18349
rect 8808 18315 8820 18349
rect 8762 18281 8820 18315
rect 8762 18247 8774 18281
rect 8808 18247 8820 18281
rect 8762 18213 8820 18247
rect 8762 18179 8774 18213
rect 8808 18179 8820 18213
rect 8762 18145 8820 18179
rect 8762 18111 8774 18145
rect 8808 18111 8820 18145
rect 8762 18077 8820 18111
rect 8762 18043 8774 18077
rect 8808 18043 8820 18077
rect 8762 18009 8820 18043
rect 8762 17975 8774 18009
rect 8808 17975 8820 18009
rect 8762 17941 8820 17975
rect 8762 17907 8774 17941
rect 8808 17907 8820 17941
rect 8762 17873 8820 17907
rect 8762 17839 8774 17873
rect 8808 17839 8820 17873
rect 8762 17805 8820 17839
rect 8762 17771 8774 17805
rect 8808 17771 8820 17805
rect 8762 17737 8820 17771
rect 8762 17703 8774 17737
rect 8808 17703 8820 17737
rect 8762 17669 8820 17703
rect 8762 17635 8774 17669
rect 8808 17635 8820 17669
rect 8762 17592 8820 17635
rect 9220 18349 9278 18392
rect 9220 18315 9232 18349
rect 9266 18315 9278 18349
rect 9220 18281 9278 18315
rect 9220 18247 9232 18281
rect 9266 18247 9278 18281
rect 9220 18213 9278 18247
rect 9220 18179 9232 18213
rect 9266 18179 9278 18213
rect 9220 18145 9278 18179
rect 9220 18111 9232 18145
rect 9266 18111 9278 18145
rect 9220 18077 9278 18111
rect 9220 18043 9232 18077
rect 9266 18043 9278 18077
rect 9220 18009 9278 18043
rect 9220 17975 9232 18009
rect 9266 17975 9278 18009
rect 9220 17941 9278 17975
rect 9220 17907 9232 17941
rect 9266 17907 9278 17941
rect 9220 17873 9278 17907
rect 9220 17839 9232 17873
rect 9266 17839 9278 17873
rect 9220 17805 9278 17839
rect 9220 17771 9232 17805
rect 9266 17771 9278 17805
rect 9220 17737 9278 17771
rect 9220 17703 9232 17737
rect 9266 17703 9278 17737
rect 9220 17669 9278 17703
rect 9220 17635 9232 17669
rect 9266 17635 9278 17669
rect 9220 17592 9278 17635
rect 9678 18349 9736 18392
rect 9678 18315 9690 18349
rect 9724 18315 9736 18349
rect 9678 18281 9736 18315
rect 9678 18247 9690 18281
rect 9724 18247 9736 18281
rect 9678 18213 9736 18247
rect 9678 18179 9690 18213
rect 9724 18179 9736 18213
rect 9678 18145 9736 18179
rect 9678 18111 9690 18145
rect 9724 18111 9736 18145
rect 9678 18077 9736 18111
rect 9678 18043 9690 18077
rect 9724 18043 9736 18077
rect 9678 18009 9736 18043
rect 9678 17975 9690 18009
rect 9724 17975 9736 18009
rect 9678 17941 9736 17975
rect 9678 17907 9690 17941
rect 9724 17907 9736 17941
rect 9678 17873 9736 17907
rect 9678 17839 9690 17873
rect 9724 17839 9736 17873
rect 9678 17805 9736 17839
rect 9678 17771 9690 17805
rect 9724 17771 9736 17805
rect 9678 17737 9736 17771
rect 9678 17703 9690 17737
rect 9724 17703 9736 17737
rect 9678 17669 9736 17703
rect 9678 17635 9690 17669
rect 9724 17635 9736 17669
rect 9678 17592 9736 17635
rect 10136 18349 10194 18392
rect 10136 18315 10148 18349
rect 10182 18315 10194 18349
rect 10136 18281 10194 18315
rect 10136 18247 10148 18281
rect 10182 18247 10194 18281
rect 10136 18213 10194 18247
rect 10136 18179 10148 18213
rect 10182 18179 10194 18213
rect 10136 18145 10194 18179
rect 10136 18111 10148 18145
rect 10182 18111 10194 18145
rect 10136 18077 10194 18111
rect 10136 18043 10148 18077
rect 10182 18043 10194 18077
rect 10136 18009 10194 18043
rect 10136 17975 10148 18009
rect 10182 17975 10194 18009
rect 10136 17941 10194 17975
rect 10136 17907 10148 17941
rect 10182 17907 10194 17941
rect 10136 17873 10194 17907
rect 10136 17839 10148 17873
rect 10182 17839 10194 17873
rect 10136 17805 10194 17839
rect 10136 17771 10148 17805
rect 10182 17771 10194 17805
rect 10136 17737 10194 17771
rect 10136 17703 10148 17737
rect 10182 17703 10194 17737
rect 10136 17669 10194 17703
rect 10136 17635 10148 17669
rect 10182 17635 10194 17669
rect 10136 17592 10194 17635
<< pdiff >>
rect 15065 41181 15123 41197
rect 15065 41147 15077 41181
rect 15111 41147 15123 41181
rect 15065 41113 15123 41147
rect 15065 41079 15077 41113
rect 15111 41079 15123 41113
rect 15065 41045 15123 41079
rect 15065 41011 15077 41045
rect 15111 41011 15123 41045
rect 15065 40977 15123 41011
rect 15065 40943 15077 40977
rect 15111 40943 15123 40977
rect 15065 40909 15123 40943
rect 15065 40875 15077 40909
rect 15111 40875 15123 40909
rect 15065 40841 15123 40875
rect 15065 40807 15077 40841
rect 15111 40807 15123 40841
rect 15065 40773 15123 40807
rect 15065 40739 15077 40773
rect 15111 40739 15123 40773
rect 15065 40705 15123 40739
rect 15065 40671 15077 40705
rect 15111 40671 15123 40705
rect 15065 40637 15123 40671
rect 15065 40603 15077 40637
rect 15111 40603 15123 40637
rect 15065 40569 15123 40603
rect 15065 40535 15077 40569
rect 15111 40535 15123 40569
rect 15065 40501 15123 40535
rect 15065 40467 15077 40501
rect 15111 40467 15123 40501
rect 15065 40433 15123 40467
rect 15065 40399 15077 40433
rect 15111 40399 15123 40433
rect 15065 40365 15123 40399
rect 15065 40331 15077 40365
rect 15111 40331 15123 40365
rect 15065 40297 15123 40331
rect 15065 40263 15077 40297
rect 15111 40263 15123 40297
rect 15065 40229 15123 40263
rect 15065 40195 15077 40229
rect 15111 40195 15123 40229
rect 15065 40161 15123 40195
rect 15065 40127 15077 40161
rect 15111 40127 15123 40161
rect 15065 40093 15123 40127
rect 15065 40059 15077 40093
rect 15111 40059 15123 40093
rect 15065 40025 15123 40059
rect 15065 39991 15077 40025
rect 15111 39991 15123 40025
rect 15065 39957 15123 39991
rect 15065 39923 15077 39957
rect 15111 39923 15123 39957
rect 15065 39907 15123 39923
rect 15523 41181 15581 41197
rect 15523 41147 15535 41181
rect 15569 41147 15581 41181
rect 15523 41113 15581 41147
rect 15523 41079 15535 41113
rect 15569 41079 15581 41113
rect 15523 41045 15581 41079
rect 15523 41011 15535 41045
rect 15569 41011 15581 41045
rect 15523 40977 15581 41011
rect 15523 40943 15535 40977
rect 15569 40943 15581 40977
rect 15523 40909 15581 40943
rect 15523 40875 15535 40909
rect 15569 40875 15581 40909
rect 15523 40841 15581 40875
rect 15523 40807 15535 40841
rect 15569 40807 15581 40841
rect 15523 40773 15581 40807
rect 15523 40739 15535 40773
rect 15569 40739 15581 40773
rect 15523 40705 15581 40739
rect 15523 40671 15535 40705
rect 15569 40671 15581 40705
rect 15523 40637 15581 40671
rect 15523 40603 15535 40637
rect 15569 40603 15581 40637
rect 15523 40569 15581 40603
rect 15523 40535 15535 40569
rect 15569 40535 15581 40569
rect 15523 40501 15581 40535
rect 15523 40467 15535 40501
rect 15569 40467 15581 40501
rect 15523 40433 15581 40467
rect 15523 40399 15535 40433
rect 15569 40399 15581 40433
rect 15523 40365 15581 40399
rect 15523 40331 15535 40365
rect 15569 40331 15581 40365
rect 15523 40297 15581 40331
rect 15523 40263 15535 40297
rect 15569 40263 15581 40297
rect 15523 40229 15581 40263
rect 15523 40195 15535 40229
rect 15569 40195 15581 40229
rect 15523 40161 15581 40195
rect 15523 40127 15535 40161
rect 15569 40127 15581 40161
rect 15523 40093 15581 40127
rect 15523 40059 15535 40093
rect 15569 40059 15581 40093
rect 15523 40025 15581 40059
rect 15523 39991 15535 40025
rect 15569 39991 15581 40025
rect 15523 39957 15581 39991
rect 15523 39923 15535 39957
rect 15569 39923 15581 39957
rect 15523 39907 15581 39923
rect 15981 41181 16039 41197
rect 15981 41147 15993 41181
rect 16027 41147 16039 41181
rect 15981 41113 16039 41147
rect 15981 41079 15993 41113
rect 16027 41079 16039 41113
rect 15981 41045 16039 41079
rect 15981 41011 15993 41045
rect 16027 41011 16039 41045
rect 15981 40977 16039 41011
rect 15981 40943 15993 40977
rect 16027 40943 16039 40977
rect 15981 40909 16039 40943
rect 15981 40875 15993 40909
rect 16027 40875 16039 40909
rect 15981 40841 16039 40875
rect 15981 40807 15993 40841
rect 16027 40807 16039 40841
rect 15981 40773 16039 40807
rect 15981 40739 15993 40773
rect 16027 40739 16039 40773
rect 15981 40705 16039 40739
rect 15981 40671 15993 40705
rect 16027 40671 16039 40705
rect 15981 40637 16039 40671
rect 15981 40603 15993 40637
rect 16027 40603 16039 40637
rect 15981 40569 16039 40603
rect 15981 40535 15993 40569
rect 16027 40535 16039 40569
rect 15981 40501 16039 40535
rect 15981 40467 15993 40501
rect 16027 40467 16039 40501
rect 15981 40433 16039 40467
rect 15981 40399 15993 40433
rect 16027 40399 16039 40433
rect 15981 40365 16039 40399
rect 15981 40331 15993 40365
rect 16027 40331 16039 40365
rect 15981 40297 16039 40331
rect 15981 40263 15993 40297
rect 16027 40263 16039 40297
rect 15981 40229 16039 40263
rect 15981 40195 15993 40229
rect 16027 40195 16039 40229
rect 15981 40161 16039 40195
rect 15981 40127 15993 40161
rect 16027 40127 16039 40161
rect 15981 40093 16039 40127
rect 15981 40059 15993 40093
rect 16027 40059 16039 40093
rect 15981 40025 16039 40059
rect 15981 39991 15993 40025
rect 16027 39991 16039 40025
rect 15981 39957 16039 39991
rect 15981 39923 15993 39957
rect 16027 39923 16039 39957
rect 15981 39907 16039 39923
rect 16439 41181 16497 41197
rect 16439 41147 16451 41181
rect 16485 41147 16497 41181
rect 16439 41113 16497 41147
rect 16439 41079 16451 41113
rect 16485 41079 16497 41113
rect 16439 41045 16497 41079
rect 16439 41011 16451 41045
rect 16485 41011 16497 41045
rect 16439 40977 16497 41011
rect 16439 40943 16451 40977
rect 16485 40943 16497 40977
rect 16439 40909 16497 40943
rect 16439 40875 16451 40909
rect 16485 40875 16497 40909
rect 16439 40841 16497 40875
rect 16439 40807 16451 40841
rect 16485 40807 16497 40841
rect 16439 40773 16497 40807
rect 16439 40739 16451 40773
rect 16485 40739 16497 40773
rect 16439 40705 16497 40739
rect 16439 40671 16451 40705
rect 16485 40671 16497 40705
rect 16439 40637 16497 40671
rect 16439 40603 16451 40637
rect 16485 40603 16497 40637
rect 16439 40569 16497 40603
rect 16439 40535 16451 40569
rect 16485 40535 16497 40569
rect 16439 40501 16497 40535
rect 16439 40467 16451 40501
rect 16485 40467 16497 40501
rect 16439 40433 16497 40467
rect 16439 40399 16451 40433
rect 16485 40399 16497 40433
rect 16439 40365 16497 40399
rect 16439 40331 16451 40365
rect 16485 40331 16497 40365
rect 16439 40297 16497 40331
rect 16439 40263 16451 40297
rect 16485 40263 16497 40297
rect 16439 40229 16497 40263
rect 16439 40195 16451 40229
rect 16485 40195 16497 40229
rect 16439 40161 16497 40195
rect 16439 40127 16451 40161
rect 16485 40127 16497 40161
rect 16439 40093 16497 40127
rect 16439 40059 16451 40093
rect 16485 40059 16497 40093
rect 16439 40025 16497 40059
rect 16439 39991 16451 40025
rect 16485 39991 16497 40025
rect 16439 39957 16497 39991
rect 16439 39923 16451 39957
rect 16485 39923 16497 39957
rect 16439 39907 16497 39923
rect 16897 41181 16955 41197
rect 16897 41147 16909 41181
rect 16943 41147 16955 41181
rect 16897 41113 16955 41147
rect 16897 41079 16909 41113
rect 16943 41079 16955 41113
rect 16897 41045 16955 41079
rect 16897 41011 16909 41045
rect 16943 41011 16955 41045
rect 16897 40977 16955 41011
rect 16897 40943 16909 40977
rect 16943 40943 16955 40977
rect 16897 40909 16955 40943
rect 16897 40875 16909 40909
rect 16943 40875 16955 40909
rect 16897 40841 16955 40875
rect 16897 40807 16909 40841
rect 16943 40807 16955 40841
rect 16897 40773 16955 40807
rect 16897 40739 16909 40773
rect 16943 40739 16955 40773
rect 16897 40705 16955 40739
rect 16897 40671 16909 40705
rect 16943 40671 16955 40705
rect 16897 40637 16955 40671
rect 16897 40603 16909 40637
rect 16943 40603 16955 40637
rect 16897 40569 16955 40603
rect 16897 40535 16909 40569
rect 16943 40535 16955 40569
rect 16897 40501 16955 40535
rect 16897 40467 16909 40501
rect 16943 40467 16955 40501
rect 16897 40433 16955 40467
rect 16897 40399 16909 40433
rect 16943 40399 16955 40433
rect 16897 40365 16955 40399
rect 16897 40331 16909 40365
rect 16943 40331 16955 40365
rect 16897 40297 16955 40331
rect 16897 40263 16909 40297
rect 16943 40263 16955 40297
rect 16897 40229 16955 40263
rect 16897 40195 16909 40229
rect 16943 40195 16955 40229
rect 16897 40161 16955 40195
rect 16897 40127 16909 40161
rect 16943 40127 16955 40161
rect 16897 40093 16955 40127
rect 16897 40059 16909 40093
rect 16943 40059 16955 40093
rect 16897 40025 16955 40059
rect 16897 39991 16909 40025
rect 16943 39991 16955 40025
rect 16897 39957 16955 39991
rect 16897 39923 16909 39957
rect 16943 39923 16955 39957
rect 16897 39907 16955 39923
rect 17355 41181 17413 41197
rect 17355 41147 17367 41181
rect 17401 41147 17413 41181
rect 17355 41113 17413 41147
rect 17355 41079 17367 41113
rect 17401 41079 17413 41113
rect 17355 41045 17413 41079
rect 17355 41011 17367 41045
rect 17401 41011 17413 41045
rect 17355 40977 17413 41011
rect 17355 40943 17367 40977
rect 17401 40943 17413 40977
rect 17355 40909 17413 40943
rect 17355 40875 17367 40909
rect 17401 40875 17413 40909
rect 17355 40841 17413 40875
rect 17355 40807 17367 40841
rect 17401 40807 17413 40841
rect 17355 40773 17413 40807
rect 17355 40739 17367 40773
rect 17401 40739 17413 40773
rect 17355 40705 17413 40739
rect 17355 40671 17367 40705
rect 17401 40671 17413 40705
rect 17355 40637 17413 40671
rect 17355 40603 17367 40637
rect 17401 40603 17413 40637
rect 17355 40569 17413 40603
rect 17355 40535 17367 40569
rect 17401 40535 17413 40569
rect 17355 40501 17413 40535
rect 17355 40467 17367 40501
rect 17401 40467 17413 40501
rect 17355 40433 17413 40467
rect 17355 40399 17367 40433
rect 17401 40399 17413 40433
rect 17355 40365 17413 40399
rect 17355 40331 17367 40365
rect 17401 40331 17413 40365
rect 17355 40297 17413 40331
rect 17355 40263 17367 40297
rect 17401 40263 17413 40297
rect 17355 40229 17413 40263
rect 17355 40195 17367 40229
rect 17401 40195 17413 40229
rect 17355 40161 17413 40195
rect 17355 40127 17367 40161
rect 17401 40127 17413 40161
rect 17355 40093 17413 40127
rect 17355 40059 17367 40093
rect 17401 40059 17413 40093
rect 17355 40025 17413 40059
rect 17355 39991 17367 40025
rect 17401 39991 17413 40025
rect 17355 39957 17413 39991
rect 17355 39923 17367 39957
rect 17401 39923 17413 39957
rect 17355 39907 17413 39923
rect 17813 41181 17871 41197
rect 17813 41147 17825 41181
rect 17859 41147 17871 41181
rect 17813 41113 17871 41147
rect 17813 41079 17825 41113
rect 17859 41079 17871 41113
rect 17813 41045 17871 41079
rect 17813 41011 17825 41045
rect 17859 41011 17871 41045
rect 17813 40977 17871 41011
rect 17813 40943 17825 40977
rect 17859 40943 17871 40977
rect 17813 40909 17871 40943
rect 17813 40875 17825 40909
rect 17859 40875 17871 40909
rect 17813 40841 17871 40875
rect 17813 40807 17825 40841
rect 17859 40807 17871 40841
rect 17813 40773 17871 40807
rect 17813 40739 17825 40773
rect 17859 40739 17871 40773
rect 17813 40705 17871 40739
rect 17813 40671 17825 40705
rect 17859 40671 17871 40705
rect 17813 40637 17871 40671
rect 17813 40603 17825 40637
rect 17859 40603 17871 40637
rect 17813 40569 17871 40603
rect 17813 40535 17825 40569
rect 17859 40535 17871 40569
rect 17813 40501 17871 40535
rect 17813 40467 17825 40501
rect 17859 40467 17871 40501
rect 17813 40433 17871 40467
rect 17813 40399 17825 40433
rect 17859 40399 17871 40433
rect 17813 40365 17871 40399
rect 17813 40331 17825 40365
rect 17859 40331 17871 40365
rect 17813 40297 17871 40331
rect 17813 40263 17825 40297
rect 17859 40263 17871 40297
rect 17813 40229 17871 40263
rect 17813 40195 17825 40229
rect 17859 40195 17871 40229
rect 17813 40161 17871 40195
rect 17813 40127 17825 40161
rect 17859 40127 17871 40161
rect 17813 40093 17871 40127
rect 17813 40059 17825 40093
rect 17859 40059 17871 40093
rect 17813 40025 17871 40059
rect 17813 39991 17825 40025
rect 17859 39991 17871 40025
rect 17813 39957 17871 39991
rect 17813 39923 17825 39957
rect 17859 39923 17871 39957
rect 17813 39907 17871 39923
rect 18271 41181 18329 41197
rect 18271 41147 18283 41181
rect 18317 41147 18329 41181
rect 18271 41113 18329 41147
rect 18271 41079 18283 41113
rect 18317 41079 18329 41113
rect 18271 41045 18329 41079
rect 18271 41011 18283 41045
rect 18317 41011 18329 41045
rect 18271 40977 18329 41011
rect 18271 40943 18283 40977
rect 18317 40943 18329 40977
rect 18271 40909 18329 40943
rect 18271 40875 18283 40909
rect 18317 40875 18329 40909
rect 18271 40841 18329 40875
rect 18271 40807 18283 40841
rect 18317 40807 18329 40841
rect 18271 40773 18329 40807
rect 18271 40739 18283 40773
rect 18317 40739 18329 40773
rect 18271 40705 18329 40739
rect 18271 40671 18283 40705
rect 18317 40671 18329 40705
rect 18271 40637 18329 40671
rect 18271 40603 18283 40637
rect 18317 40603 18329 40637
rect 18271 40569 18329 40603
rect 18271 40535 18283 40569
rect 18317 40535 18329 40569
rect 18271 40501 18329 40535
rect 18271 40467 18283 40501
rect 18317 40467 18329 40501
rect 18271 40433 18329 40467
rect 18271 40399 18283 40433
rect 18317 40399 18329 40433
rect 18271 40365 18329 40399
rect 18271 40331 18283 40365
rect 18317 40331 18329 40365
rect 18271 40297 18329 40331
rect 18271 40263 18283 40297
rect 18317 40263 18329 40297
rect 18271 40229 18329 40263
rect 18271 40195 18283 40229
rect 18317 40195 18329 40229
rect 18271 40161 18329 40195
rect 18271 40127 18283 40161
rect 18317 40127 18329 40161
rect 18271 40093 18329 40127
rect 18271 40059 18283 40093
rect 18317 40059 18329 40093
rect 18271 40025 18329 40059
rect 18271 39991 18283 40025
rect 18317 39991 18329 40025
rect 18271 39957 18329 39991
rect 18271 39923 18283 39957
rect 18317 39923 18329 39957
rect 18271 39907 18329 39923
rect 18729 41181 18787 41197
rect 18729 41147 18741 41181
rect 18775 41147 18787 41181
rect 18729 41113 18787 41147
rect 18729 41079 18741 41113
rect 18775 41079 18787 41113
rect 18729 41045 18787 41079
rect 18729 41011 18741 41045
rect 18775 41011 18787 41045
rect 18729 40977 18787 41011
rect 18729 40943 18741 40977
rect 18775 40943 18787 40977
rect 18729 40909 18787 40943
rect 18729 40875 18741 40909
rect 18775 40875 18787 40909
rect 18729 40841 18787 40875
rect 18729 40807 18741 40841
rect 18775 40807 18787 40841
rect 18729 40773 18787 40807
rect 18729 40739 18741 40773
rect 18775 40739 18787 40773
rect 18729 40705 18787 40739
rect 18729 40671 18741 40705
rect 18775 40671 18787 40705
rect 18729 40637 18787 40671
rect 18729 40603 18741 40637
rect 18775 40603 18787 40637
rect 18729 40569 18787 40603
rect 18729 40535 18741 40569
rect 18775 40535 18787 40569
rect 18729 40501 18787 40535
rect 18729 40467 18741 40501
rect 18775 40467 18787 40501
rect 18729 40433 18787 40467
rect 18729 40399 18741 40433
rect 18775 40399 18787 40433
rect 18729 40365 18787 40399
rect 18729 40331 18741 40365
rect 18775 40331 18787 40365
rect 18729 40297 18787 40331
rect 18729 40263 18741 40297
rect 18775 40263 18787 40297
rect 18729 40229 18787 40263
rect 18729 40195 18741 40229
rect 18775 40195 18787 40229
rect 18729 40161 18787 40195
rect 18729 40127 18741 40161
rect 18775 40127 18787 40161
rect 18729 40093 18787 40127
rect 18729 40059 18741 40093
rect 18775 40059 18787 40093
rect 18729 40025 18787 40059
rect 18729 39991 18741 40025
rect 18775 39991 18787 40025
rect 18729 39957 18787 39991
rect 18729 39923 18741 39957
rect 18775 39923 18787 39957
rect 18729 39907 18787 39923
rect 19187 41181 19245 41197
rect 19187 41147 19199 41181
rect 19233 41147 19245 41181
rect 19187 41113 19245 41147
rect 19187 41079 19199 41113
rect 19233 41079 19245 41113
rect 19187 41045 19245 41079
rect 19187 41011 19199 41045
rect 19233 41011 19245 41045
rect 19187 40977 19245 41011
rect 19187 40943 19199 40977
rect 19233 40943 19245 40977
rect 19187 40909 19245 40943
rect 19187 40875 19199 40909
rect 19233 40875 19245 40909
rect 19187 40841 19245 40875
rect 19187 40807 19199 40841
rect 19233 40807 19245 40841
rect 19187 40773 19245 40807
rect 19187 40739 19199 40773
rect 19233 40739 19245 40773
rect 19187 40705 19245 40739
rect 19187 40671 19199 40705
rect 19233 40671 19245 40705
rect 19187 40637 19245 40671
rect 19187 40603 19199 40637
rect 19233 40603 19245 40637
rect 19187 40569 19245 40603
rect 19187 40535 19199 40569
rect 19233 40535 19245 40569
rect 19187 40501 19245 40535
rect 19187 40467 19199 40501
rect 19233 40467 19245 40501
rect 19187 40433 19245 40467
rect 19187 40399 19199 40433
rect 19233 40399 19245 40433
rect 19187 40365 19245 40399
rect 19187 40331 19199 40365
rect 19233 40331 19245 40365
rect 19187 40297 19245 40331
rect 19187 40263 19199 40297
rect 19233 40263 19245 40297
rect 19187 40229 19245 40263
rect 19187 40195 19199 40229
rect 19233 40195 19245 40229
rect 19187 40161 19245 40195
rect 19187 40127 19199 40161
rect 19233 40127 19245 40161
rect 19187 40093 19245 40127
rect 19187 40059 19199 40093
rect 19233 40059 19245 40093
rect 19187 40025 19245 40059
rect 19187 39991 19199 40025
rect 19233 39991 19245 40025
rect 19187 39957 19245 39991
rect 19187 39923 19199 39957
rect 19233 39923 19245 39957
rect 19187 39907 19245 39923
rect 19645 41181 19703 41197
rect 19645 41147 19657 41181
rect 19691 41147 19703 41181
rect 19645 41113 19703 41147
rect 19645 41079 19657 41113
rect 19691 41079 19703 41113
rect 19645 41045 19703 41079
rect 19645 41011 19657 41045
rect 19691 41011 19703 41045
rect 19645 40977 19703 41011
rect 19645 40943 19657 40977
rect 19691 40943 19703 40977
rect 19645 40909 19703 40943
rect 19645 40875 19657 40909
rect 19691 40875 19703 40909
rect 19645 40841 19703 40875
rect 19645 40807 19657 40841
rect 19691 40807 19703 40841
rect 19645 40773 19703 40807
rect 19645 40739 19657 40773
rect 19691 40739 19703 40773
rect 19645 40705 19703 40739
rect 19645 40671 19657 40705
rect 19691 40671 19703 40705
rect 19645 40637 19703 40671
rect 19645 40603 19657 40637
rect 19691 40603 19703 40637
rect 19645 40569 19703 40603
rect 19645 40535 19657 40569
rect 19691 40535 19703 40569
rect 19645 40501 19703 40535
rect 19645 40467 19657 40501
rect 19691 40467 19703 40501
rect 19645 40433 19703 40467
rect 19645 40399 19657 40433
rect 19691 40399 19703 40433
rect 19645 40365 19703 40399
rect 19645 40331 19657 40365
rect 19691 40331 19703 40365
rect 19645 40297 19703 40331
rect 19645 40263 19657 40297
rect 19691 40263 19703 40297
rect 19645 40229 19703 40263
rect 19645 40195 19657 40229
rect 19691 40195 19703 40229
rect 19645 40161 19703 40195
rect 19645 40127 19657 40161
rect 19691 40127 19703 40161
rect 19645 40093 19703 40127
rect 19645 40059 19657 40093
rect 19691 40059 19703 40093
rect 19645 40025 19703 40059
rect 19645 39991 19657 40025
rect 19691 39991 19703 40025
rect 19645 39957 19703 39991
rect 19645 39923 19657 39957
rect 19691 39923 19703 39957
rect 19645 39907 19703 39923
rect 20103 41181 20161 41197
rect 20103 41147 20115 41181
rect 20149 41147 20161 41181
rect 20103 41113 20161 41147
rect 20103 41079 20115 41113
rect 20149 41079 20161 41113
rect 20103 41045 20161 41079
rect 20103 41011 20115 41045
rect 20149 41011 20161 41045
rect 20103 40977 20161 41011
rect 20103 40943 20115 40977
rect 20149 40943 20161 40977
rect 20103 40909 20161 40943
rect 20103 40875 20115 40909
rect 20149 40875 20161 40909
rect 20103 40841 20161 40875
rect 20103 40807 20115 40841
rect 20149 40807 20161 40841
rect 20103 40773 20161 40807
rect 20103 40739 20115 40773
rect 20149 40739 20161 40773
rect 20103 40705 20161 40739
rect 20103 40671 20115 40705
rect 20149 40671 20161 40705
rect 20103 40637 20161 40671
rect 20103 40603 20115 40637
rect 20149 40603 20161 40637
rect 20103 40569 20161 40603
rect 20103 40535 20115 40569
rect 20149 40535 20161 40569
rect 20103 40501 20161 40535
rect 20103 40467 20115 40501
rect 20149 40467 20161 40501
rect 20103 40433 20161 40467
rect 20103 40399 20115 40433
rect 20149 40399 20161 40433
rect 20103 40365 20161 40399
rect 20103 40331 20115 40365
rect 20149 40331 20161 40365
rect 20103 40297 20161 40331
rect 20103 40263 20115 40297
rect 20149 40263 20161 40297
rect 20103 40229 20161 40263
rect 20103 40195 20115 40229
rect 20149 40195 20161 40229
rect 20103 40161 20161 40195
rect 20103 40127 20115 40161
rect 20149 40127 20161 40161
rect 20103 40093 20161 40127
rect 20103 40059 20115 40093
rect 20149 40059 20161 40093
rect 20103 40025 20161 40059
rect 20103 39991 20115 40025
rect 20149 39991 20161 40025
rect 20103 39957 20161 39991
rect 20103 39923 20115 39957
rect 20149 39923 20161 39957
rect 20103 39907 20161 39923
rect 20561 41181 20619 41197
rect 20561 41147 20573 41181
rect 20607 41147 20619 41181
rect 20561 41113 20619 41147
rect 20561 41079 20573 41113
rect 20607 41079 20619 41113
rect 20561 41045 20619 41079
rect 20561 41011 20573 41045
rect 20607 41011 20619 41045
rect 20561 40977 20619 41011
rect 20561 40943 20573 40977
rect 20607 40943 20619 40977
rect 20561 40909 20619 40943
rect 20561 40875 20573 40909
rect 20607 40875 20619 40909
rect 20561 40841 20619 40875
rect 20561 40807 20573 40841
rect 20607 40807 20619 40841
rect 20561 40773 20619 40807
rect 20561 40739 20573 40773
rect 20607 40739 20619 40773
rect 20561 40705 20619 40739
rect 20561 40671 20573 40705
rect 20607 40671 20619 40705
rect 20561 40637 20619 40671
rect 20561 40603 20573 40637
rect 20607 40603 20619 40637
rect 20561 40569 20619 40603
rect 20561 40535 20573 40569
rect 20607 40535 20619 40569
rect 20561 40501 20619 40535
rect 20561 40467 20573 40501
rect 20607 40467 20619 40501
rect 20561 40433 20619 40467
rect 20561 40399 20573 40433
rect 20607 40399 20619 40433
rect 20561 40365 20619 40399
rect 20561 40331 20573 40365
rect 20607 40331 20619 40365
rect 20561 40297 20619 40331
rect 20561 40263 20573 40297
rect 20607 40263 20619 40297
rect 20561 40229 20619 40263
rect 20561 40195 20573 40229
rect 20607 40195 20619 40229
rect 20561 40161 20619 40195
rect 20561 40127 20573 40161
rect 20607 40127 20619 40161
rect 20561 40093 20619 40127
rect 20561 40059 20573 40093
rect 20607 40059 20619 40093
rect 20561 40025 20619 40059
rect 20561 39991 20573 40025
rect 20607 39991 20619 40025
rect 20561 39957 20619 39991
rect 20561 39923 20573 39957
rect 20607 39923 20619 39957
rect 20561 39907 20619 39923
rect 21019 41181 21077 41197
rect 21019 41147 21031 41181
rect 21065 41147 21077 41181
rect 21019 41113 21077 41147
rect 21019 41079 21031 41113
rect 21065 41079 21077 41113
rect 21019 41045 21077 41079
rect 21019 41011 21031 41045
rect 21065 41011 21077 41045
rect 21019 40977 21077 41011
rect 21019 40943 21031 40977
rect 21065 40943 21077 40977
rect 21019 40909 21077 40943
rect 21019 40875 21031 40909
rect 21065 40875 21077 40909
rect 21019 40841 21077 40875
rect 21019 40807 21031 40841
rect 21065 40807 21077 40841
rect 21019 40773 21077 40807
rect 21019 40739 21031 40773
rect 21065 40739 21077 40773
rect 21019 40705 21077 40739
rect 21019 40671 21031 40705
rect 21065 40671 21077 40705
rect 21019 40637 21077 40671
rect 21019 40603 21031 40637
rect 21065 40603 21077 40637
rect 21019 40569 21077 40603
rect 21019 40535 21031 40569
rect 21065 40535 21077 40569
rect 21019 40501 21077 40535
rect 21019 40467 21031 40501
rect 21065 40467 21077 40501
rect 21019 40433 21077 40467
rect 21019 40399 21031 40433
rect 21065 40399 21077 40433
rect 21019 40365 21077 40399
rect 21019 40331 21031 40365
rect 21065 40331 21077 40365
rect 21019 40297 21077 40331
rect 21019 40263 21031 40297
rect 21065 40263 21077 40297
rect 21019 40229 21077 40263
rect 21019 40195 21031 40229
rect 21065 40195 21077 40229
rect 21019 40161 21077 40195
rect 21019 40127 21031 40161
rect 21065 40127 21077 40161
rect 21019 40093 21077 40127
rect 21019 40059 21031 40093
rect 21065 40059 21077 40093
rect 21019 40025 21077 40059
rect 21019 39991 21031 40025
rect 21065 39991 21077 40025
rect 21019 39957 21077 39991
rect 21019 39923 21031 39957
rect 21065 39923 21077 39957
rect 21019 39907 21077 39923
rect 21477 41181 21535 41197
rect 21477 41147 21489 41181
rect 21523 41147 21535 41181
rect 21477 41113 21535 41147
rect 21477 41079 21489 41113
rect 21523 41079 21535 41113
rect 21477 41045 21535 41079
rect 21477 41011 21489 41045
rect 21523 41011 21535 41045
rect 21477 40977 21535 41011
rect 21477 40943 21489 40977
rect 21523 40943 21535 40977
rect 21477 40909 21535 40943
rect 21477 40875 21489 40909
rect 21523 40875 21535 40909
rect 21477 40841 21535 40875
rect 21477 40807 21489 40841
rect 21523 40807 21535 40841
rect 21477 40773 21535 40807
rect 21477 40739 21489 40773
rect 21523 40739 21535 40773
rect 21477 40705 21535 40739
rect 21477 40671 21489 40705
rect 21523 40671 21535 40705
rect 21477 40637 21535 40671
rect 21477 40603 21489 40637
rect 21523 40603 21535 40637
rect 21477 40569 21535 40603
rect 21477 40535 21489 40569
rect 21523 40535 21535 40569
rect 21477 40501 21535 40535
rect 21477 40467 21489 40501
rect 21523 40467 21535 40501
rect 21477 40433 21535 40467
rect 21477 40399 21489 40433
rect 21523 40399 21535 40433
rect 21477 40365 21535 40399
rect 21477 40331 21489 40365
rect 21523 40331 21535 40365
rect 21477 40297 21535 40331
rect 21477 40263 21489 40297
rect 21523 40263 21535 40297
rect 21477 40229 21535 40263
rect 21477 40195 21489 40229
rect 21523 40195 21535 40229
rect 21477 40161 21535 40195
rect 21477 40127 21489 40161
rect 21523 40127 21535 40161
rect 21477 40093 21535 40127
rect 21477 40059 21489 40093
rect 21523 40059 21535 40093
rect 21477 40025 21535 40059
rect 21477 39991 21489 40025
rect 21523 39991 21535 40025
rect 21477 39957 21535 39991
rect 21477 39923 21489 39957
rect 21523 39923 21535 39957
rect 21477 39907 21535 39923
rect 21935 41181 21993 41197
rect 21935 41147 21947 41181
rect 21981 41147 21993 41181
rect 21935 41113 21993 41147
rect 21935 41079 21947 41113
rect 21981 41079 21993 41113
rect 21935 41045 21993 41079
rect 21935 41011 21947 41045
rect 21981 41011 21993 41045
rect 21935 40977 21993 41011
rect 21935 40943 21947 40977
rect 21981 40943 21993 40977
rect 21935 40909 21993 40943
rect 21935 40875 21947 40909
rect 21981 40875 21993 40909
rect 21935 40841 21993 40875
rect 21935 40807 21947 40841
rect 21981 40807 21993 40841
rect 21935 40773 21993 40807
rect 21935 40739 21947 40773
rect 21981 40739 21993 40773
rect 21935 40705 21993 40739
rect 21935 40671 21947 40705
rect 21981 40671 21993 40705
rect 21935 40637 21993 40671
rect 21935 40603 21947 40637
rect 21981 40603 21993 40637
rect 21935 40569 21993 40603
rect 21935 40535 21947 40569
rect 21981 40535 21993 40569
rect 21935 40501 21993 40535
rect 21935 40467 21947 40501
rect 21981 40467 21993 40501
rect 21935 40433 21993 40467
rect 21935 40399 21947 40433
rect 21981 40399 21993 40433
rect 21935 40365 21993 40399
rect 21935 40331 21947 40365
rect 21981 40331 21993 40365
rect 21935 40297 21993 40331
rect 21935 40263 21947 40297
rect 21981 40263 21993 40297
rect 21935 40229 21993 40263
rect 21935 40195 21947 40229
rect 21981 40195 21993 40229
rect 21935 40161 21993 40195
rect 21935 40127 21947 40161
rect 21981 40127 21993 40161
rect 21935 40093 21993 40127
rect 21935 40059 21947 40093
rect 21981 40059 21993 40093
rect 21935 40025 21993 40059
rect 21935 39991 21947 40025
rect 21981 39991 21993 40025
rect 21935 39957 21993 39991
rect 21935 39923 21947 39957
rect 21981 39923 21993 39957
rect 21935 39907 21993 39923
rect 22393 41181 22451 41197
rect 22393 41147 22405 41181
rect 22439 41147 22451 41181
rect 22393 41113 22451 41147
rect 22393 41079 22405 41113
rect 22439 41079 22451 41113
rect 22393 41045 22451 41079
rect 22393 41011 22405 41045
rect 22439 41011 22451 41045
rect 22393 40977 22451 41011
rect 22393 40943 22405 40977
rect 22439 40943 22451 40977
rect 22393 40909 22451 40943
rect 22393 40875 22405 40909
rect 22439 40875 22451 40909
rect 22393 40841 22451 40875
rect 22393 40807 22405 40841
rect 22439 40807 22451 40841
rect 22393 40773 22451 40807
rect 22393 40739 22405 40773
rect 22439 40739 22451 40773
rect 22393 40705 22451 40739
rect 22393 40671 22405 40705
rect 22439 40671 22451 40705
rect 22393 40637 22451 40671
rect 22393 40603 22405 40637
rect 22439 40603 22451 40637
rect 22393 40569 22451 40603
rect 22393 40535 22405 40569
rect 22439 40535 22451 40569
rect 22393 40501 22451 40535
rect 22393 40467 22405 40501
rect 22439 40467 22451 40501
rect 22393 40433 22451 40467
rect 22393 40399 22405 40433
rect 22439 40399 22451 40433
rect 22393 40365 22451 40399
rect 22393 40331 22405 40365
rect 22439 40331 22451 40365
rect 22393 40297 22451 40331
rect 22393 40263 22405 40297
rect 22439 40263 22451 40297
rect 22393 40229 22451 40263
rect 22393 40195 22405 40229
rect 22439 40195 22451 40229
rect 22393 40161 22451 40195
rect 22393 40127 22405 40161
rect 22439 40127 22451 40161
rect 22393 40093 22451 40127
rect 22393 40059 22405 40093
rect 22439 40059 22451 40093
rect 22393 40025 22451 40059
rect 22393 39991 22405 40025
rect 22439 39991 22451 40025
rect 22393 39957 22451 39991
rect 22393 39923 22405 39957
rect 22439 39923 22451 39957
rect 22393 39907 22451 39923
rect 22851 41181 22909 41197
rect 22851 41147 22863 41181
rect 22897 41147 22909 41181
rect 22851 41113 22909 41147
rect 22851 41079 22863 41113
rect 22897 41079 22909 41113
rect 22851 41045 22909 41079
rect 22851 41011 22863 41045
rect 22897 41011 22909 41045
rect 22851 40977 22909 41011
rect 22851 40943 22863 40977
rect 22897 40943 22909 40977
rect 22851 40909 22909 40943
rect 22851 40875 22863 40909
rect 22897 40875 22909 40909
rect 22851 40841 22909 40875
rect 22851 40807 22863 40841
rect 22897 40807 22909 40841
rect 22851 40773 22909 40807
rect 22851 40739 22863 40773
rect 22897 40739 22909 40773
rect 22851 40705 22909 40739
rect 22851 40671 22863 40705
rect 22897 40671 22909 40705
rect 22851 40637 22909 40671
rect 22851 40603 22863 40637
rect 22897 40603 22909 40637
rect 22851 40569 22909 40603
rect 22851 40535 22863 40569
rect 22897 40535 22909 40569
rect 22851 40501 22909 40535
rect 22851 40467 22863 40501
rect 22897 40467 22909 40501
rect 22851 40433 22909 40467
rect 22851 40399 22863 40433
rect 22897 40399 22909 40433
rect 22851 40365 22909 40399
rect 22851 40331 22863 40365
rect 22897 40331 22909 40365
rect 22851 40297 22909 40331
rect 22851 40263 22863 40297
rect 22897 40263 22909 40297
rect 22851 40229 22909 40263
rect 22851 40195 22863 40229
rect 22897 40195 22909 40229
rect 22851 40161 22909 40195
rect 22851 40127 22863 40161
rect 22897 40127 22909 40161
rect 22851 40093 22909 40127
rect 22851 40059 22863 40093
rect 22897 40059 22909 40093
rect 22851 40025 22909 40059
rect 22851 39991 22863 40025
rect 22897 39991 22909 40025
rect 22851 39957 22909 39991
rect 22851 39923 22863 39957
rect 22897 39923 22909 39957
rect 22851 39907 22909 39923
rect 23309 41181 23367 41197
rect 23309 41147 23321 41181
rect 23355 41147 23367 41181
rect 23309 41113 23367 41147
rect 23309 41079 23321 41113
rect 23355 41079 23367 41113
rect 23309 41045 23367 41079
rect 23309 41011 23321 41045
rect 23355 41011 23367 41045
rect 23309 40977 23367 41011
rect 23309 40943 23321 40977
rect 23355 40943 23367 40977
rect 23309 40909 23367 40943
rect 23309 40875 23321 40909
rect 23355 40875 23367 40909
rect 23309 40841 23367 40875
rect 23309 40807 23321 40841
rect 23355 40807 23367 40841
rect 23309 40773 23367 40807
rect 23309 40739 23321 40773
rect 23355 40739 23367 40773
rect 23309 40705 23367 40739
rect 23309 40671 23321 40705
rect 23355 40671 23367 40705
rect 23309 40637 23367 40671
rect 23309 40603 23321 40637
rect 23355 40603 23367 40637
rect 23309 40569 23367 40603
rect 23309 40535 23321 40569
rect 23355 40535 23367 40569
rect 23309 40501 23367 40535
rect 23309 40467 23321 40501
rect 23355 40467 23367 40501
rect 23309 40433 23367 40467
rect 23309 40399 23321 40433
rect 23355 40399 23367 40433
rect 23309 40365 23367 40399
rect 23309 40331 23321 40365
rect 23355 40331 23367 40365
rect 23309 40297 23367 40331
rect 23309 40263 23321 40297
rect 23355 40263 23367 40297
rect 23309 40229 23367 40263
rect 23309 40195 23321 40229
rect 23355 40195 23367 40229
rect 23309 40161 23367 40195
rect 23309 40127 23321 40161
rect 23355 40127 23367 40161
rect 23309 40093 23367 40127
rect 23309 40059 23321 40093
rect 23355 40059 23367 40093
rect 23309 40025 23367 40059
rect 23309 39991 23321 40025
rect 23355 39991 23367 40025
rect 23309 39957 23367 39991
rect 23309 39923 23321 39957
rect 23355 39923 23367 39957
rect 23309 39907 23367 39923
rect 23767 41181 23825 41197
rect 23767 41147 23779 41181
rect 23813 41147 23825 41181
rect 23767 41113 23825 41147
rect 23767 41079 23779 41113
rect 23813 41079 23825 41113
rect 23767 41045 23825 41079
rect 23767 41011 23779 41045
rect 23813 41011 23825 41045
rect 23767 40977 23825 41011
rect 23767 40943 23779 40977
rect 23813 40943 23825 40977
rect 23767 40909 23825 40943
rect 23767 40875 23779 40909
rect 23813 40875 23825 40909
rect 23767 40841 23825 40875
rect 23767 40807 23779 40841
rect 23813 40807 23825 40841
rect 23767 40773 23825 40807
rect 23767 40739 23779 40773
rect 23813 40739 23825 40773
rect 23767 40705 23825 40739
rect 23767 40671 23779 40705
rect 23813 40671 23825 40705
rect 23767 40637 23825 40671
rect 23767 40603 23779 40637
rect 23813 40603 23825 40637
rect 23767 40569 23825 40603
rect 23767 40535 23779 40569
rect 23813 40535 23825 40569
rect 23767 40501 23825 40535
rect 23767 40467 23779 40501
rect 23813 40467 23825 40501
rect 23767 40433 23825 40467
rect 23767 40399 23779 40433
rect 23813 40399 23825 40433
rect 23767 40365 23825 40399
rect 23767 40331 23779 40365
rect 23813 40331 23825 40365
rect 23767 40297 23825 40331
rect 23767 40263 23779 40297
rect 23813 40263 23825 40297
rect 23767 40229 23825 40263
rect 23767 40195 23779 40229
rect 23813 40195 23825 40229
rect 23767 40161 23825 40195
rect 23767 40127 23779 40161
rect 23813 40127 23825 40161
rect 23767 40093 23825 40127
rect 23767 40059 23779 40093
rect 23813 40059 23825 40093
rect 23767 40025 23825 40059
rect 23767 39991 23779 40025
rect 23813 39991 23825 40025
rect 23767 39957 23825 39991
rect 23767 39923 23779 39957
rect 23813 39923 23825 39957
rect 23767 39907 23825 39923
rect 24225 41181 24283 41197
rect 24225 41147 24237 41181
rect 24271 41147 24283 41181
rect 24225 41113 24283 41147
rect 24225 41079 24237 41113
rect 24271 41079 24283 41113
rect 24225 41045 24283 41079
rect 24225 41011 24237 41045
rect 24271 41011 24283 41045
rect 24225 40977 24283 41011
rect 24225 40943 24237 40977
rect 24271 40943 24283 40977
rect 24225 40909 24283 40943
rect 24225 40875 24237 40909
rect 24271 40875 24283 40909
rect 24225 40841 24283 40875
rect 24225 40807 24237 40841
rect 24271 40807 24283 40841
rect 24225 40773 24283 40807
rect 24225 40739 24237 40773
rect 24271 40739 24283 40773
rect 24225 40705 24283 40739
rect 24225 40671 24237 40705
rect 24271 40671 24283 40705
rect 24225 40637 24283 40671
rect 24225 40603 24237 40637
rect 24271 40603 24283 40637
rect 24225 40569 24283 40603
rect 24225 40535 24237 40569
rect 24271 40535 24283 40569
rect 24225 40501 24283 40535
rect 24225 40467 24237 40501
rect 24271 40467 24283 40501
rect 24225 40433 24283 40467
rect 24225 40399 24237 40433
rect 24271 40399 24283 40433
rect 24225 40365 24283 40399
rect 24225 40331 24237 40365
rect 24271 40331 24283 40365
rect 24225 40297 24283 40331
rect 24225 40263 24237 40297
rect 24271 40263 24283 40297
rect 24225 40229 24283 40263
rect 24225 40195 24237 40229
rect 24271 40195 24283 40229
rect 24225 40161 24283 40195
rect 24225 40127 24237 40161
rect 24271 40127 24283 40161
rect 24225 40093 24283 40127
rect 24225 40059 24237 40093
rect 24271 40059 24283 40093
rect 24225 40025 24283 40059
rect 24225 39991 24237 40025
rect 24271 39991 24283 40025
rect 24225 39957 24283 39991
rect 24225 39923 24237 39957
rect 24271 39923 24283 39957
rect 24225 39907 24283 39923
rect 24683 41181 24741 41197
rect 24683 41147 24695 41181
rect 24729 41147 24741 41181
rect 24683 41113 24741 41147
rect 24683 41079 24695 41113
rect 24729 41079 24741 41113
rect 24683 41045 24741 41079
rect 24683 41011 24695 41045
rect 24729 41011 24741 41045
rect 24683 40977 24741 41011
rect 24683 40943 24695 40977
rect 24729 40943 24741 40977
rect 24683 40909 24741 40943
rect 24683 40875 24695 40909
rect 24729 40875 24741 40909
rect 24683 40841 24741 40875
rect 24683 40807 24695 40841
rect 24729 40807 24741 40841
rect 24683 40773 24741 40807
rect 24683 40739 24695 40773
rect 24729 40739 24741 40773
rect 24683 40705 24741 40739
rect 24683 40671 24695 40705
rect 24729 40671 24741 40705
rect 24683 40637 24741 40671
rect 24683 40603 24695 40637
rect 24729 40603 24741 40637
rect 24683 40569 24741 40603
rect 24683 40535 24695 40569
rect 24729 40535 24741 40569
rect 24683 40501 24741 40535
rect 24683 40467 24695 40501
rect 24729 40467 24741 40501
rect 24683 40433 24741 40467
rect 24683 40399 24695 40433
rect 24729 40399 24741 40433
rect 24683 40365 24741 40399
rect 24683 40331 24695 40365
rect 24729 40331 24741 40365
rect 24683 40297 24741 40331
rect 24683 40263 24695 40297
rect 24729 40263 24741 40297
rect 24683 40229 24741 40263
rect 24683 40195 24695 40229
rect 24729 40195 24741 40229
rect 24683 40161 24741 40195
rect 24683 40127 24695 40161
rect 24729 40127 24741 40161
rect 24683 40093 24741 40127
rect 24683 40059 24695 40093
rect 24729 40059 24741 40093
rect 24683 40025 24741 40059
rect 24683 39991 24695 40025
rect 24729 39991 24741 40025
rect 24683 39957 24741 39991
rect 24683 39923 24695 39957
rect 24729 39923 24741 39957
rect 24683 39907 24741 39923
rect 25141 41181 25199 41197
rect 25141 41147 25153 41181
rect 25187 41147 25199 41181
rect 25141 41113 25199 41147
rect 25141 41079 25153 41113
rect 25187 41079 25199 41113
rect 25141 41045 25199 41079
rect 25141 41011 25153 41045
rect 25187 41011 25199 41045
rect 25141 40977 25199 41011
rect 25141 40943 25153 40977
rect 25187 40943 25199 40977
rect 25141 40909 25199 40943
rect 25141 40875 25153 40909
rect 25187 40875 25199 40909
rect 25141 40841 25199 40875
rect 25141 40807 25153 40841
rect 25187 40807 25199 40841
rect 25141 40773 25199 40807
rect 25141 40739 25153 40773
rect 25187 40739 25199 40773
rect 25141 40705 25199 40739
rect 25141 40671 25153 40705
rect 25187 40671 25199 40705
rect 25141 40637 25199 40671
rect 25141 40603 25153 40637
rect 25187 40603 25199 40637
rect 25141 40569 25199 40603
rect 25141 40535 25153 40569
rect 25187 40535 25199 40569
rect 25141 40501 25199 40535
rect 25141 40467 25153 40501
rect 25187 40467 25199 40501
rect 25141 40433 25199 40467
rect 25141 40399 25153 40433
rect 25187 40399 25199 40433
rect 25141 40365 25199 40399
rect 25141 40331 25153 40365
rect 25187 40331 25199 40365
rect 25141 40297 25199 40331
rect 25141 40263 25153 40297
rect 25187 40263 25199 40297
rect 25141 40229 25199 40263
rect 25141 40195 25153 40229
rect 25187 40195 25199 40229
rect 25141 40161 25199 40195
rect 25141 40127 25153 40161
rect 25187 40127 25199 40161
rect 25141 40093 25199 40127
rect 25141 40059 25153 40093
rect 25187 40059 25199 40093
rect 25141 40025 25199 40059
rect 25141 39991 25153 40025
rect 25187 39991 25199 40025
rect 25141 39957 25199 39991
rect 25141 39923 25153 39957
rect 25187 39923 25199 39957
rect 25141 39907 25199 39923
rect 25599 41181 25657 41197
rect 25599 41147 25611 41181
rect 25645 41147 25657 41181
rect 25599 41113 25657 41147
rect 25599 41079 25611 41113
rect 25645 41079 25657 41113
rect 25599 41045 25657 41079
rect 25599 41011 25611 41045
rect 25645 41011 25657 41045
rect 25599 40977 25657 41011
rect 25599 40943 25611 40977
rect 25645 40943 25657 40977
rect 25599 40909 25657 40943
rect 25599 40875 25611 40909
rect 25645 40875 25657 40909
rect 25599 40841 25657 40875
rect 25599 40807 25611 40841
rect 25645 40807 25657 40841
rect 25599 40773 25657 40807
rect 25599 40739 25611 40773
rect 25645 40739 25657 40773
rect 25599 40705 25657 40739
rect 25599 40671 25611 40705
rect 25645 40671 25657 40705
rect 25599 40637 25657 40671
rect 25599 40603 25611 40637
rect 25645 40603 25657 40637
rect 25599 40569 25657 40603
rect 25599 40535 25611 40569
rect 25645 40535 25657 40569
rect 25599 40501 25657 40535
rect 25599 40467 25611 40501
rect 25645 40467 25657 40501
rect 25599 40433 25657 40467
rect 25599 40399 25611 40433
rect 25645 40399 25657 40433
rect 25599 40365 25657 40399
rect 25599 40331 25611 40365
rect 25645 40331 25657 40365
rect 25599 40297 25657 40331
rect 25599 40263 25611 40297
rect 25645 40263 25657 40297
rect 25599 40229 25657 40263
rect 25599 40195 25611 40229
rect 25645 40195 25657 40229
rect 25599 40161 25657 40195
rect 25599 40127 25611 40161
rect 25645 40127 25657 40161
rect 25599 40093 25657 40127
rect 25599 40059 25611 40093
rect 25645 40059 25657 40093
rect 25599 40025 25657 40059
rect 25599 39991 25611 40025
rect 25645 39991 25657 40025
rect 25599 39957 25657 39991
rect 25599 39923 25611 39957
rect 25645 39923 25657 39957
rect 25599 39907 25657 39923
rect 26057 41181 26115 41197
rect 26057 41147 26069 41181
rect 26103 41147 26115 41181
rect 26057 41113 26115 41147
rect 26057 41079 26069 41113
rect 26103 41079 26115 41113
rect 26057 41045 26115 41079
rect 26057 41011 26069 41045
rect 26103 41011 26115 41045
rect 26057 40977 26115 41011
rect 26057 40943 26069 40977
rect 26103 40943 26115 40977
rect 26057 40909 26115 40943
rect 26057 40875 26069 40909
rect 26103 40875 26115 40909
rect 26057 40841 26115 40875
rect 26057 40807 26069 40841
rect 26103 40807 26115 40841
rect 26057 40773 26115 40807
rect 26057 40739 26069 40773
rect 26103 40739 26115 40773
rect 26057 40705 26115 40739
rect 26057 40671 26069 40705
rect 26103 40671 26115 40705
rect 26057 40637 26115 40671
rect 26057 40603 26069 40637
rect 26103 40603 26115 40637
rect 26057 40569 26115 40603
rect 26057 40535 26069 40569
rect 26103 40535 26115 40569
rect 26057 40501 26115 40535
rect 26057 40467 26069 40501
rect 26103 40467 26115 40501
rect 26057 40433 26115 40467
rect 26057 40399 26069 40433
rect 26103 40399 26115 40433
rect 26057 40365 26115 40399
rect 26057 40331 26069 40365
rect 26103 40331 26115 40365
rect 26057 40297 26115 40331
rect 26057 40263 26069 40297
rect 26103 40263 26115 40297
rect 26057 40229 26115 40263
rect 26057 40195 26069 40229
rect 26103 40195 26115 40229
rect 26057 40161 26115 40195
rect 26057 40127 26069 40161
rect 26103 40127 26115 40161
rect 26057 40093 26115 40127
rect 26057 40059 26069 40093
rect 26103 40059 26115 40093
rect 26057 40025 26115 40059
rect 26057 39991 26069 40025
rect 26103 39991 26115 40025
rect 26057 39957 26115 39991
rect 26057 39923 26069 39957
rect 26103 39923 26115 39957
rect 26057 39907 26115 39923
rect 26515 41181 26573 41197
rect 26515 41147 26527 41181
rect 26561 41147 26573 41181
rect 26515 41113 26573 41147
rect 26515 41079 26527 41113
rect 26561 41079 26573 41113
rect 26515 41045 26573 41079
rect 26515 41011 26527 41045
rect 26561 41011 26573 41045
rect 26515 40977 26573 41011
rect 26515 40943 26527 40977
rect 26561 40943 26573 40977
rect 26515 40909 26573 40943
rect 26515 40875 26527 40909
rect 26561 40875 26573 40909
rect 26515 40841 26573 40875
rect 26515 40807 26527 40841
rect 26561 40807 26573 40841
rect 26515 40773 26573 40807
rect 26515 40739 26527 40773
rect 26561 40739 26573 40773
rect 26515 40705 26573 40739
rect 26515 40671 26527 40705
rect 26561 40671 26573 40705
rect 26515 40637 26573 40671
rect 26515 40603 26527 40637
rect 26561 40603 26573 40637
rect 26515 40569 26573 40603
rect 26515 40535 26527 40569
rect 26561 40535 26573 40569
rect 26515 40501 26573 40535
rect 26515 40467 26527 40501
rect 26561 40467 26573 40501
rect 26515 40433 26573 40467
rect 26515 40399 26527 40433
rect 26561 40399 26573 40433
rect 26515 40365 26573 40399
rect 26515 40331 26527 40365
rect 26561 40331 26573 40365
rect 26515 40297 26573 40331
rect 26515 40263 26527 40297
rect 26561 40263 26573 40297
rect 26515 40229 26573 40263
rect 26515 40195 26527 40229
rect 26561 40195 26573 40229
rect 26515 40161 26573 40195
rect 26515 40127 26527 40161
rect 26561 40127 26573 40161
rect 26515 40093 26573 40127
rect 26515 40059 26527 40093
rect 26561 40059 26573 40093
rect 26515 40025 26573 40059
rect 26515 39991 26527 40025
rect 26561 39991 26573 40025
rect 26515 39957 26573 39991
rect 26515 39923 26527 39957
rect 26561 39923 26573 39957
rect 26515 39907 26573 39923
rect 26973 41181 27031 41197
rect 26973 41147 26985 41181
rect 27019 41147 27031 41181
rect 26973 41113 27031 41147
rect 26973 41079 26985 41113
rect 27019 41079 27031 41113
rect 26973 41045 27031 41079
rect 26973 41011 26985 41045
rect 27019 41011 27031 41045
rect 26973 40977 27031 41011
rect 26973 40943 26985 40977
rect 27019 40943 27031 40977
rect 26973 40909 27031 40943
rect 26973 40875 26985 40909
rect 27019 40875 27031 40909
rect 26973 40841 27031 40875
rect 26973 40807 26985 40841
rect 27019 40807 27031 40841
rect 26973 40773 27031 40807
rect 26973 40739 26985 40773
rect 27019 40739 27031 40773
rect 26973 40705 27031 40739
rect 26973 40671 26985 40705
rect 27019 40671 27031 40705
rect 26973 40637 27031 40671
rect 26973 40603 26985 40637
rect 27019 40603 27031 40637
rect 26973 40569 27031 40603
rect 26973 40535 26985 40569
rect 27019 40535 27031 40569
rect 26973 40501 27031 40535
rect 26973 40467 26985 40501
rect 27019 40467 27031 40501
rect 26973 40433 27031 40467
rect 26973 40399 26985 40433
rect 27019 40399 27031 40433
rect 26973 40365 27031 40399
rect 26973 40331 26985 40365
rect 27019 40331 27031 40365
rect 26973 40297 27031 40331
rect 26973 40263 26985 40297
rect 27019 40263 27031 40297
rect 26973 40229 27031 40263
rect 26973 40195 26985 40229
rect 27019 40195 27031 40229
rect 26973 40161 27031 40195
rect 26973 40127 26985 40161
rect 27019 40127 27031 40161
rect 26973 40093 27031 40127
rect 26973 40059 26985 40093
rect 27019 40059 27031 40093
rect 26973 40025 27031 40059
rect 26973 39991 26985 40025
rect 27019 39991 27031 40025
rect 26973 39957 27031 39991
rect 26973 39923 26985 39957
rect 27019 39923 27031 39957
rect 26973 39907 27031 39923
rect 27431 41181 27489 41197
rect 27431 41147 27443 41181
rect 27477 41147 27489 41181
rect 27431 41113 27489 41147
rect 27431 41079 27443 41113
rect 27477 41079 27489 41113
rect 27431 41045 27489 41079
rect 27431 41011 27443 41045
rect 27477 41011 27489 41045
rect 27431 40977 27489 41011
rect 27431 40943 27443 40977
rect 27477 40943 27489 40977
rect 27431 40909 27489 40943
rect 27431 40875 27443 40909
rect 27477 40875 27489 40909
rect 27431 40841 27489 40875
rect 27431 40807 27443 40841
rect 27477 40807 27489 40841
rect 27431 40773 27489 40807
rect 27431 40739 27443 40773
rect 27477 40739 27489 40773
rect 27431 40705 27489 40739
rect 27431 40671 27443 40705
rect 27477 40671 27489 40705
rect 27431 40637 27489 40671
rect 27431 40603 27443 40637
rect 27477 40603 27489 40637
rect 27431 40569 27489 40603
rect 27431 40535 27443 40569
rect 27477 40535 27489 40569
rect 27431 40501 27489 40535
rect 27431 40467 27443 40501
rect 27477 40467 27489 40501
rect 27431 40433 27489 40467
rect 27431 40399 27443 40433
rect 27477 40399 27489 40433
rect 27431 40365 27489 40399
rect 27431 40331 27443 40365
rect 27477 40331 27489 40365
rect 27431 40297 27489 40331
rect 27431 40263 27443 40297
rect 27477 40263 27489 40297
rect 27431 40229 27489 40263
rect 27431 40195 27443 40229
rect 27477 40195 27489 40229
rect 27431 40161 27489 40195
rect 27431 40127 27443 40161
rect 27477 40127 27489 40161
rect 27431 40093 27489 40127
rect 27431 40059 27443 40093
rect 27477 40059 27489 40093
rect 27431 40025 27489 40059
rect 27431 39991 27443 40025
rect 27477 39991 27489 40025
rect 27431 39957 27489 39991
rect 27431 39923 27443 39957
rect 27477 39923 27489 39957
rect 27431 39907 27489 39923
rect 27889 41181 27947 41197
rect 27889 41147 27901 41181
rect 27935 41147 27947 41181
rect 27889 41113 27947 41147
rect 27889 41079 27901 41113
rect 27935 41079 27947 41113
rect 27889 41045 27947 41079
rect 27889 41011 27901 41045
rect 27935 41011 27947 41045
rect 27889 40977 27947 41011
rect 27889 40943 27901 40977
rect 27935 40943 27947 40977
rect 27889 40909 27947 40943
rect 27889 40875 27901 40909
rect 27935 40875 27947 40909
rect 27889 40841 27947 40875
rect 27889 40807 27901 40841
rect 27935 40807 27947 40841
rect 27889 40773 27947 40807
rect 27889 40739 27901 40773
rect 27935 40739 27947 40773
rect 27889 40705 27947 40739
rect 27889 40671 27901 40705
rect 27935 40671 27947 40705
rect 27889 40637 27947 40671
rect 27889 40603 27901 40637
rect 27935 40603 27947 40637
rect 27889 40569 27947 40603
rect 27889 40535 27901 40569
rect 27935 40535 27947 40569
rect 27889 40501 27947 40535
rect 27889 40467 27901 40501
rect 27935 40467 27947 40501
rect 27889 40433 27947 40467
rect 27889 40399 27901 40433
rect 27935 40399 27947 40433
rect 27889 40365 27947 40399
rect 27889 40331 27901 40365
rect 27935 40331 27947 40365
rect 27889 40297 27947 40331
rect 27889 40263 27901 40297
rect 27935 40263 27947 40297
rect 27889 40229 27947 40263
rect 27889 40195 27901 40229
rect 27935 40195 27947 40229
rect 27889 40161 27947 40195
rect 27889 40127 27901 40161
rect 27935 40127 27947 40161
rect 27889 40093 27947 40127
rect 27889 40059 27901 40093
rect 27935 40059 27947 40093
rect 27889 40025 27947 40059
rect 27889 39991 27901 40025
rect 27935 39991 27947 40025
rect 27889 39957 27947 39991
rect 27889 39923 27901 39957
rect 27935 39923 27947 39957
rect 27889 39907 27947 39923
rect 28347 41181 28405 41197
rect 28347 41147 28359 41181
rect 28393 41147 28405 41181
rect 28347 41113 28405 41147
rect 28347 41079 28359 41113
rect 28393 41079 28405 41113
rect 28347 41045 28405 41079
rect 28347 41011 28359 41045
rect 28393 41011 28405 41045
rect 28347 40977 28405 41011
rect 28347 40943 28359 40977
rect 28393 40943 28405 40977
rect 28347 40909 28405 40943
rect 28347 40875 28359 40909
rect 28393 40875 28405 40909
rect 28347 40841 28405 40875
rect 28347 40807 28359 40841
rect 28393 40807 28405 40841
rect 28347 40773 28405 40807
rect 28347 40739 28359 40773
rect 28393 40739 28405 40773
rect 28347 40705 28405 40739
rect 28347 40671 28359 40705
rect 28393 40671 28405 40705
rect 28347 40637 28405 40671
rect 28347 40603 28359 40637
rect 28393 40603 28405 40637
rect 28347 40569 28405 40603
rect 28347 40535 28359 40569
rect 28393 40535 28405 40569
rect 28347 40501 28405 40535
rect 28347 40467 28359 40501
rect 28393 40467 28405 40501
rect 28347 40433 28405 40467
rect 28347 40399 28359 40433
rect 28393 40399 28405 40433
rect 28347 40365 28405 40399
rect 28347 40331 28359 40365
rect 28393 40331 28405 40365
rect 28347 40297 28405 40331
rect 28347 40263 28359 40297
rect 28393 40263 28405 40297
rect 28347 40229 28405 40263
rect 28347 40195 28359 40229
rect 28393 40195 28405 40229
rect 28347 40161 28405 40195
rect 28347 40127 28359 40161
rect 28393 40127 28405 40161
rect 28347 40093 28405 40127
rect 28347 40059 28359 40093
rect 28393 40059 28405 40093
rect 28347 40025 28405 40059
rect 28347 39991 28359 40025
rect 28393 39991 28405 40025
rect 28347 39957 28405 39991
rect 28347 39923 28359 39957
rect 28393 39923 28405 39957
rect 28347 39907 28405 39923
rect 28805 41181 28863 41197
rect 28805 41147 28817 41181
rect 28851 41147 28863 41181
rect 28805 41113 28863 41147
rect 28805 41079 28817 41113
rect 28851 41079 28863 41113
rect 28805 41045 28863 41079
rect 28805 41011 28817 41045
rect 28851 41011 28863 41045
rect 28805 40977 28863 41011
rect 28805 40943 28817 40977
rect 28851 40943 28863 40977
rect 28805 40909 28863 40943
rect 28805 40875 28817 40909
rect 28851 40875 28863 40909
rect 28805 40841 28863 40875
rect 28805 40807 28817 40841
rect 28851 40807 28863 40841
rect 28805 40773 28863 40807
rect 28805 40739 28817 40773
rect 28851 40739 28863 40773
rect 28805 40705 28863 40739
rect 28805 40671 28817 40705
rect 28851 40671 28863 40705
rect 28805 40637 28863 40671
rect 28805 40603 28817 40637
rect 28851 40603 28863 40637
rect 28805 40569 28863 40603
rect 28805 40535 28817 40569
rect 28851 40535 28863 40569
rect 28805 40501 28863 40535
rect 28805 40467 28817 40501
rect 28851 40467 28863 40501
rect 28805 40433 28863 40467
rect 28805 40399 28817 40433
rect 28851 40399 28863 40433
rect 28805 40365 28863 40399
rect 28805 40331 28817 40365
rect 28851 40331 28863 40365
rect 28805 40297 28863 40331
rect 28805 40263 28817 40297
rect 28851 40263 28863 40297
rect 28805 40229 28863 40263
rect 28805 40195 28817 40229
rect 28851 40195 28863 40229
rect 28805 40161 28863 40195
rect 28805 40127 28817 40161
rect 28851 40127 28863 40161
rect 28805 40093 28863 40127
rect 28805 40059 28817 40093
rect 28851 40059 28863 40093
rect 28805 40025 28863 40059
rect 28805 39991 28817 40025
rect 28851 39991 28863 40025
rect 28805 39957 28863 39991
rect 28805 39923 28817 39957
rect 28851 39923 28863 39957
rect 28805 39907 28863 39923
rect 29263 41181 29321 41197
rect 29263 41147 29275 41181
rect 29309 41147 29321 41181
rect 29263 41113 29321 41147
rect 29263 41079 29275 41113
rect 29309 41079 29321 41113
rect 29263 41045 29321 41079
rect 29263 41011 29275 41045
rect 29309 41011 29321 41045
rect 29263 40977 29321 41011
rect 29263 40943 29275 40977
rect 29309 40943 29321 40977
rect 29263 40909 29321 40943
rect 29263 40875 29275 40909
rect 29309 40875 29321 40909
rect 29263 40841 29321 40875
rect 29263 40807 29275 40841
rect 29309 40807 29321 40841
rect 29263 40773 29321 40807
rect 29263 40739 29275 40773
rect 29309 40739 29321 40773
rect 29263 40705 29321 40739
rect 29263 40671 29275 40705
rect 29309 40671 29321 40705
rect 29263 40637 29321 40671
rect 29263 40603 29275 40637
rect 29309 40603 29321 40637
rect 29263 40569 29321 40603
rect 29263 40535 29275 40569
rect 29309 40535 29321 40569
rect 29263 40501 29321 40535
rect 29263 40467 29275 40501
rect 29309 40467 29321 40501
rect 29263 40433 29321 40467
rect 29263 40399 29275 40433
rect 29309 40399 29321 40433
rect 29263 40365 29321 40399
rect 29263 40331 29275 40365
rect 29309 40331 29321 40365
rect 29263 40297 29321 40331
rect 29263 40263 29275 40297
rect 29309 40263 29321 40297
rect 29263 40229 29321 40263
rect 29263 40195 29275 40229
rect 29309 40195 29321 40229
rect 29263 40161 29321 40195
rect 29263 40127 29275 40161
rect 29309 40127 29321 40161
rect 29263 40093 29321 40127
rect 29263 40059 29275 40093
rect 29309 40059 29321 40093
rect 29263 40025 29321 40059
rect 29263 39991 29275 40025
rect 29309 39991 29321 40025
rect 29263 39957 29321 39991
rect 29263 39923 29275 39957
rect 29309 39923 29321 39957
rect 29263 39907 29321 39923
rect 29721 41181 29779 41197
rect 29721 41147 29733 41181
rect 29767 41147 29779 41181
rect 29721 41113 29779 41147
rect 29721 41079 29733 41113
rect 29767 41079 29779 41113
rect 29721 41045 29779 41079
rect 29721 41011 29733 41045
rect 29767 41011 29779 41045
rect 29721 40977 29779 41011
rect 29721 40943 29733 40977
rect 29767 40943 29779 40977
rect 29721 40909 29779 40943
rect 29721 40875 29733 40909
rect 29767 40875 29779 40909
rect 29721 40841 29779 40875
rect 29721 40807 29733 40841
rect 29767 40807 29779 40841
rect 29721 40773 29779 40807
rect 29721 40739 29733 40773
rect 29767 40739 29779 40773
rect 29721 40705 29779 40739
rect 29721 40671 29733 40705
rect 29767 40671 29779 40705
rect 29721 40637 29779 40671
rect 29721 40603 29733 40637
rect 29767 40603 29779 40637
rect 29721 40569 29779 40603
rect 29721 40535 29733 40569
rect 29767 40535 29779 40569
rect 29721 40501 29779 40535
rect 29721 40467 29733 40501
rect 29767 40467 29779 40501
rect 29721 40433 29779 40467
rect 29721 40399 29733 40433
rect 29767 40399 29779 40433
rect 29721 40365 29779 40399
rect 29721 40331 29733 40365
rect 29767 40331 29779 40365
rect 29721 40297 29779 40331
rect 29721 40263 29733 40297
rect 29767 40263 29779 40297
rect 29721 40229 29779 40263
rect 29721 40195 29733 40229
rect 29767 40195 29779 40229
rect 29721 40161 29779 40195
rect 29721 40127 29733 40161
rect 29767 40127 29779 40161
rect 29721 40093 29779 40127
rect 29721 40059 29733 40093
rect 29767 40059 29779 40093
rect 29721 40025 29779 40059
rect 29721 39991 29733 40025
rect 29767 39991 29779 40025
rect 29721 39957 29779 39991
rect 29721 39923 29733 39957
rect 29767 39923 29779 39957
rect 29721 39907 29779 39923
rect 30179 41181 30237 41197
rect 30179 41147 30191 41181
rect 30225 41147 30237 41181
rect 30179 41113 30237 41147
rect 30179 41079 30191 41113
rect 30225 41079 30237 41113
rect 30179 41045 30237 41079
rect 30179 41011 30191 41045
rect 30225 41011 30237 41045
rect 30179 40977 30237 41011
rect 30179 40943 30191 40977
rect 30225 40943 30237 40977
rect 30179 40909 30237 40943
rect 30179 40875 30191 40909
rect 30225 40875 30237 40909
rect 30179 40841 30237 40875
rect 30179 40807 30191 40841
rect 30225 40807 30237 40841
rect 30179 40773 30237 40807
rect 30179 40739 30191 40773
rect 30225 40739 30237 40773
rect 30179 40705 30237 40739
rect 30179 40671 30191 40705
rect 30225 40671 30237 40705
rect 30179 40637 30237 40671
rect 30179 40603 30191 40637
rect 30225 40603 30237 40637
rect 30179 40569 30237 40603
rect 30179 40535 30191 40569
rect 30225 40535 30237 40569
rect 30179 40501 30237 40535
rect 30179 40467 30191 40501
rect 30225 40467 30237 40501
rect 30179 40433 30237 40467
rect 30179 40399 30191 40433
rect 30225 40399 30237 40433
rect 30179 40365 30237 40399
rect 30179 40331 30191 40365
rect 30225 40331 30237 40365
rect 30179 40297 30237 40331
rect 30179 40263 30191 40297
rect 30225 40263 30237 40297
rect 30179 40229 30237 40263
rect 30179 40195 30191 40229
rect 30225 40195 30237 40229
rect 30179 40161 30237 40195
rect 30179 40127 30191 40161
rect 30225 40127 30237 40161
rect 30179 40093 30237 40127
rect 30179 40059 30191 40093
rect 30225 40059 30237 40093
rect 30179 40025 30237 40059
rect 30179 39991 30191 40025
rect 30225 39991 30237 40025
rect 30179 39957 30237 39991
rect 30179 39923 30191 39957
rect 30225 39923 30237 39957
rect 30179 39907 30237 39923
rect 30637 41181 30695 41197
rect 30637 41147 30649 41181
rect 30683 41147 30695 41181
rect 30637 41113 30695 41147
rect 30637 41079 30649 41113
rect 30683 41079 30695 41113
rect 30637 41045 30695 41079
rect 30637 41011 30649 41045
rect 30683 41011 30695 41045
rect 30637 40977 30695 41011
rect 30637 40943 30649 40977
rect 30683 40943 30695 40977
rect 30637 40909 30695 40943
rect 30637 40875 30649 40909
rect 30683 40875 30695 40909
rect 30637 40841 30695 40875
rect 30637 40807 30649 40841
rect 30683 40807 30695 40841
rect 30637 40773 30695 40807
rect 30637 40739 30649 40773
rect 30683 40739 30695 40773
rect 30637 40705 30695 40739
rect 30637 40671 30649 40705
rect 30683 40671 30695 40705
rect 30637 40637 30695 40671
rect 30637 40603 30649 40637
rect 30683 40603 30695 40637
rect 30637 40569 30695 40603
rect 30637 40535 30649 40569
rect 30683 40535 30695 40569
rect 30637 40501 30695 40535
rect 30637 40467 30649 40501
rect 30683 40467 30695 40501
rect 30637 40433 30695 40467
rect 30637 40399 30649 40433
rect 30683 40399 30695 40433
rect 30637 40365 30695 40399
rect 30637 40331 30649 40365
rect 30683 40331 30695 40365
rect 30637 40297 30695 40331
rect 30637 40263 30649 40297
rect 30683 40263 30695 40297
rect 30637 40229 30695 40263
rect 30637 40195 30649 40229
rect 30683 40195 30695 40229
rect 30637 40161 30695 40195
rect 30637 40127 30649 40161
rect 30683 40127 30695 40161
rect 30637 40093 30695 40127
rect 30637 40059 30649 40093
rect 30683 40059 30695 40093
rect 30637 40025 30695 40059
rect 30637 39991 30649 40025
rect 30683 39991 30695 40025
rect 30637 39957 30695 39991
rect 30637 39923 30649 39957
rect 30683 39923 30695 39957
rect 30637 39907 30695 39923
rect 31095 41181 31153 41197
rect 31095 41147 31107 41181
rect 31141 41147 31153 41181
rect 31095 41113 31153 41147
rect 31095 41079 31107 41113
rect 31141 41079 31153 41113
rect 31095 41045 31153 41079
rect 31095 41011 31107 41045
rect 31141 41011 31153 41045
rect 31095 40977 31153 41011
rect 31095 40943 31107 40977
rect 31141 40943 31153 40977
rect 31095 40909 31153 40943
rect 31095 40875 31107 40909
rect 31141 40875 31153 40909
rect 31095 40841 31153 40875
rect 31095 40807 31107 40841
rect 31141 40807 31153 40841
rect 31095 40773 31153 40807
rect 31095 40739 31107 40773
rect 31141 40739 31153 40773
rect 31095 40705 31153 40739
rect 31095 40671 31107 40705
rect 31141 40671 31153 40705
rect 31095 40637 31153 40671
rect 31095 40603 31107 40637
rect 31141 40603 31153 40637
rect 31095 40569 31153 40603
rect 31095 40535 31107 40569
rect 31141 40535 31153 40569
rect 31095 40501 31153 40535
rect 31095 40467 31107 40501
rect 31141 40467 31153 40501
rect 31095 40433 31153 40467
rect 31095 40399 31107 40433
rect 31141 40399 31153 40433
rect 31095 40365 31153 40399
rect 31095 40331 31107 40365
rect 31141 40331 31153 40365
rect 31095 40297 31153 40331
rect 31095 40263 31107 40297
rect 31141 40263 31153 40297
rect 31095 40229 31153 40263
rect 31095 40195 31107 40229
rect 31141 40195 31153 40229
rect 31095 40161 31153 40195
rect 31095 40127 31107 40161
rect 31141 40127 31153 40161
rect 31095 40093 31153 40127
rect 31095 40059 31107 40093
rect 31141 40059 31153 40093
rect 31095 40025 31153 40059
rect 31095 39991 31107 40025
rect 31141 39991 31153 40025
rect 31095 39957 31153 39991
rect 31095 39923 31107 39957
rect 31141 39923 31153 39957
rect 31095 39907 31153 39923
rect 31553 41181 31611 41197
rect 31553 41147 31565 41181
rect 31599 41147 31611 41181
rect 31553 41113 31611 41147
rect 31553 41079 31565 41113
rect 31599 41079 31611 41113
rect 31553 41045 31611 41079
rect 31553 41011 31565 41045
rect 31599 41011 31611 41045
rect 31553 40977 31611 41011
rect 31553 40943 31565 40977
rect 31599 40943 31611 40977
rect 31553 40909 31611 40943
rect 31553 40875 31565 40909
rect 31599 40875 31611 40909
rect 31553 40841 31611 40875
rect 31553 40807 31565 40841
rect 31599 40807 31611 40841
rect 31553 40773 31611 40807
rect 31553 40739 31565 40773
rect 31599 40739 31611 40773
rect 31553 40705 31611 40739
rect 31553 40671 31565 40705
rect 31599 40671 31611 40705
rect 31553 40637 31611 40671
rect 31553 40603 31565 40637
rect 31599 40603 31611 40637
rect 31553 40569 31611 40603
rect 31553 40535 31565 40569
rect 31599 40535 31611 40569
rect 31553 40501 31611 40535
rect 31553 40467 31565 40501
rect 31599 40467 31611 40501
rect 31553 40433 31611 40467
rect 31553 40399 31565 40433
rect 31599 40399 31611 40433
rect 31553 40365 31611 40399
rect 31553 40331 31565 40365
rect 31599 40331 31611 40365
rect 31553 40297 31611 40331
rect 31553 40263 31565 40297
rect 31599 40263 31611 40297
rect 31553 40229 31611 40263
rect 31553 40195 31565 40229
rect 31599 40195 31611 40229
rect 31553 40161 31611 40195
rect 31553 40127 31565 40161
rect 31599 40127 31611 40161
rect 31553 40093 31611 40127
rect 31553 40059 31565 40093
rect 31599 40059 31611 40093
rect 31553 40025 31611 40059
rect 31553 39991 31565 40025
rect 31599 39991 31611 40025
rect 31553 39957 31611 39991
rect 31553 39923 31565 39957
rect 31599 39923 31611 39957
rect 31553 39907 31611 39923
rect 32011 41181 32069 41197
rect 32011 41147 32023 41181
rect 32057 41147 32069 41181
rect 32011 41113 32069 41147
rect 32011 41079 32023 41113
rect 32057 41079 32069 41113
rect 32011 41045 32069 41079
rect 32011 41011 32023 41045
rect 32057 41011 32069 41045
rect 32011 40977 32069 41011
rect 32011 40943 32023 40977
rect 32057 40943 32069 40977
rect 32011 40909 32069 40943
rect 32011 40875 32023 40909
rect 32057 40875 32069 40909
rect 32011 40841 32069 40875
rect 32011 40807 32023 40841
rect 32057 40807 32069 40841
rect 32011 40773 32069 40807
rect 32011 40739 32023 40773
rect 32057 40739 32069 40773
rect 32011 40705 32069 40739
rect 32011 40671 32023 40705
rect 32057 40671 32069 40705
rect 32011 40637 32069 40671
rect 32011 40603 32023 40637
rect 32057 40603 32069 40637
rect 32011 40569 32069 40603
rect 32011 40535 32023 40569
rect 32057 40535 32069 40569
rect 32011 40501 32069 40535
rect 32011 40467 32023 40501
rect 32057 40467 32069 40501
rect 32011 40433 32069 40467
rect 32011 40399 32023 40433
rect 32057 40399 32069 40433
rect 32011 40365 32069 40399
rect 32011 40331 32023 40365
rect 32057 40331 32069 40365
rect 32011 40297 32069 40331
rect 32011 40263 32023 40297
rect 32057 40263 32069 40297
rect 32011 40229 32069 40263
rect 32011 40195 32023 40229
rect 32057 40195 32069 40229
rect 32011 40161 32069 40195
rect 32011 40127 32023 40161
rect 32057 40127 32069 40161
rect 32011 40093 32069 40127
rect 32011 40059 32023 40093
rect 32057 40059 32069 40093
rect 32011 40025 32069 40059
rect 32011 39991 32023 40025
rect 32057 39991 32069 40025
rect 32011 39957 32069 39991
rect 32011 39923 32023 39957
rect 32057 39923 32069 39957
rect 32011 39907 32069 39923
rect 32469 41181 32527 41197
rect 32469 41147 32481 41181
rect 32515 41147 32527 41181
rect 32469 41113 32527 41147
rect 32469 41079 32481 41113
rect 32515 41079 32527 41113
rect 32469 41045 32527 41079
rect 32469 41011 32481 41045
rect 32515 41011 32527 41045
rect 32469 40977 32527 41011
rect 32469 40943 32481 40977
rect 32515 40943 32527 40977
rect 32469 40909 32527 40943
rect 32469 40875 32481 40909
rect 32515 40875 32527 40909
rect 32469 40841 32527 40875
rect 32469 40807 32481 40841
rect 32515 40807 32527 40841
rect 32469 40773 32527 40807
rect 32469 40739 32481 40773
rect 32515 40739 32527 40773
rect 32469 40705 32527 40739
rect 32469 40671 32481 40705
rect 32515 40671 32527 40705
rect 32469 40637 32527 40671
rect 32469 40603 32481 40637
rect 32515 40603 32527 40637
rect 32469 40569 32527 40603
rect 32469 40535 32481 40569
rect 32515 40535 32527 40569
rect 32469 40501 32527 40535
rect 32469 40467 32481 40501
rect 32515 40467 32527 40501
rect 32469 40433 32527 40467
rect 32469 40399 32481 40433
rect 32515 40399 32527 40433
rect 32469 40365 32527 40399
rect 32469 40331 32481 40365
rect 32515 40331 32527 40365
rect 32469 40297 32527 40331
rect 32469 40263 32481 40297
rect 32515 40263 32527 40297
rect 32469 40229 32527 40263
rect 32469 40195 32481 40229
rect 32515 40195 32527 40229
rect 32469 40161 32527 40195
rect 32469 40127 32481 40161
rect 32515 40127 32527 40161
rect 32469 40093 32527 40127
rect 32469 40059 32481 40093
rect 32515 40059 32527 40093
rect 32469 40025 32527 40059
rect 32469 39991 32481 40025
rect 32515 39991 32527 40025
rect 32469 39957 32527 39991
rect 32469 39923 32481 39957
rect 32515 39923 32527 39957
rect 32469 39907 32527 39923
rect 32927 41181 32985 41197
rect 32927 41147 32939 41181
rect 32973 41147 32985 41181
rect 32927 41113 32985 41147
rect 32927 41079 32939 41113
rect 32973 41079 32985 41113
rect 32927 41045 32985 41079
rect 32927 41011 32939 41045
rect 32973 41011 32985 41045
rect 32927 40977 32985 41011
rect 32927 40943 32939 40977
rect 32973 40943 32985 40977
rect 32927 40909 32985 40943
rect 32927 40875 32939 40909
rect 32973 40875 32985 40909
rect 32927 40841 32985 40875
rect 32927 40807 32939 40841
rect 32973 40807 32985 40841
rect 32927 40773 32985 40807
rect 32927 40739 32939 40773
rect 32973 40739 32985 40773
rect 32927 40705 32985 40739
rect 32927 40671 32939 40705
rect 32973 40671 32985 40705
rect 32927 40637 32985 40671
rect 32927 40603 32939 40637
rect 32973 40603 32985 40637
rect 32927 40569 32985 40603
rect 32927 40535 32939 40569
rect 32973 40535 32985 40569
rect 32927 40501 32985 40535
rect 32927 40467 32939 40501
rect 32973 40467 32985 40501
rect 32927 40433 32985 40467
rect 32927 40399 32939 40433
rect 32973 40399 32985 40433
rect 32927 40365 32985 40399
rect 32927 40331 32939 40365
rect 32973 40331 32985 40365
rect 32927 40297 32985 40331
rect 32927 40263 32939 40297
rect 32973 40263 32985 40297
rect 32927 40229 32985 40263
rect 32927 40195 32939 40229
rect 32973 40195 32985 40229
rect 32927 40161 32985 40195
rect 32927 40127 32939 40161
rect 32973 40127 32985 40161
rect 32927 40093 32985 40127
rect 32927 40059 32939 40093
rect 32973 40059 32985 40093
rect 32927 40025 32985 40059
rect 32927 39991 32939 40025
rect 32973 39991 32985 40025
rect 32927 39957 32985 39991
rect 32927 39923 32939 39957
rect 32973 39923 32985 39957
rect 32927 39907 32985 39923
rect 33385 41181 33443 41197
rect 33385 41147 33397 41181
rect 33431 41147 33443 41181
rect 33385 41113 33443 41147
rect 33385 41079 33397 41113
rect 33431 41079 33443 41113
rect 33385 41045 33443 41079
rect 33385 41011 33397 41045
rect 33431 41011 33443 41045
rect 33385 40977 33443 41011
rect 33385 40943 33397 40977
rect 33431 40943 33443 40977
rect 33385 40909 33443 40943
rect 33385 40875 33397 40909
rect 33431 40875 33443 40909
rect 33385 40841 33443 40875
rect 33385 40807 33397 40841
rect 33431 40807 33443 40841
rect 33385 40773 33443 40807
rect 33385 40739 33397 40773
rect 33431 40739 33443 40773
rect 33385 40705 33443 40739
rect 33385 40671 33397 40705
rect 33431 40671 33443 40705
rect 33385 40637 33443 40671
rect 33385 40603 33397 40637
rect 33431 40603 33443 40637
rect 33385 40569 33443 40603
rect 33385 40535 33397 40569
rect 33431 40535 33443 40569
rect 33385 40501 33443 40535
rect 33385 40467 33397 40501
rect 33431 40467 33443 40501
rect 33385 40433 33443 40467
rect 33385 40399 33397 40433
rect 33431 40399 33443 40433
rect 33385 40365 33443 40399
rect 33385 40331 33397 40365
rect 33431 40331 33443 40365
rect 33385 40297 33443 40331
rect 33385 40263 33397 40297
rect 33431 40263 33443 40297
rect 33385 40229 33443 40263
rect 33385 40195 33397 40229
rect 33431 40195 33443 40229
rect 33385 40161 33443 40195
rect 33385 40127 33397 40161
rect 33431 40127 33443 40161
rect 33385 40093 33443 40127
rect 33385 40059 33397 40093
rect 33431 40059 33443 40093
rect 33385 40025 33443 40059
rect 33385 39991 33397 40025
rect 33431 39991 33443 40025
rect 33385 39957 33443 39991
rect 33385 39923 33397 39957
rect 33431 39923 33443 39957
rect 33385 39907 33443 39923
rect 33843 41181 33901 41197
rect 33843 41147 33855 41181
rect 33889 41147 33901 41181
rect 33843 41113 33901 41147
rect 33843 41079 33855 41113
rect 33889 41079 33901 41113
rect 33843 41045 33901 41079
rect 33843 41011 33855 41045
rect 33889 41011 33901 41045
rect 33843 40977 33901 41011
rect 33843 40943 33855 40977
rect 33889 40943 33901 40977
rect 33843 40909 33901 40943
rect 33843 40875 33855 40909
rect 33889 40875 33901 40909
rect 33843 40841 33901 40875
rect 33843 40807 33855 40841
rect 33889 40807 33901 40841
rect 33843 40773 33901 40807
rect 33843 40739 33855 40773
rect 33889 40739 33901 40773
rect 33843 40705 33901 40739
rect 33843 40671 33855 40705
rect 33889 40671 33901 40705
rect 33843 40637 33901 40671
rect 33843 40603 33855 40637
rect 33889 40603 33901 40637
rect 33843 40569 33901 40603
rect 33843 40535 33855 40569
rect 33889 40535 33901 40569
rect 33843 40501 33901 40535
rect 33843 40467 33855 40501
rect 33889 40467 33901 40501
rect 33843 40433 33901 40467
rect 33843 40399 33855 40433
rect 33889 40399 33901 40433
rect 33843 40365 33901 40399
rect 33843 40331 33855 40365
rect 33889 40331 33901 40365
rect 33843 40297 33901 40331
rect 33843 40263 33855 40297
rect 33889 40263 33901 40297
rect 33843 40229 33901 40263
rect 33843 40195 33855 40229
rect 33889 40195 33901 40229
rect 33843 40161 33901 40195
rect 33843 40127 33855 40161
rect 33889 40127 33901 40161
rect 33843 40093 33901 40127
rect 33843 40059 33855 40093
rect 33889 40059 33901 40093
rect 33843 40025 33901 40059
rect 33843 39991 33855 40025
rect 33889 39991 33901 40025
rect 33843 39957 33901 39991
rect 33843 39923 33855 39957
rect 33889 39923 33901 39957
rect 33843 39907 33901 39923
rect 34301 41181 34359 41197
rect 34301 41147 34313 41181
rect 34347 41147 34359 41181
rect 34301 41113 34359 41147
rect 34301 41079 34313 41113
rect 34347 41079 34359 41113
rect 34301 41045 34359 41079
rect 34301 41011 34313 41045
rect 34347 41011 34359 41045
rect 34301 40977 34359 41011
rect 34301 40943 34313 40977
rect 34347 40943 34359 40977
rect 34301 40909 34359 40943
rect 34301 40875 34313 40909
rect 34347 40875 34359 40909
rect 34301 40841 34359 40875
rect 34301 40807 34313 40841
rect 34347 40807 34359 40841
rect 34301 40773 34359 40807
rect 34301 40739 34313 40773
rect 34347 40739 34359 40773
rect 34301 40705 34359 40739
rect 34301 40671 34313 40705
rect 34347 40671 34359 40705
rect 34301 40637 34359 40671
rect 34301 40603 34313 40637
rect 34347 40603 34359 40637
rect 34301 40569 34359 40603
rect 34301 40535 34313 40569
rect 34347 40535 34359 40569
rect 34301 40501 34359 40535
rect 34301 40467 34313 40501
rect 34347 40467 34359 40501
rect 34301 40433 34359 40467
rect 34301 40399 34313 40433
rect 34347 40399 34359 40433
rect 34301 40365 34359 40399
rect 34301 40331 34313 40365
rect 34347 40331 34359 40365
rect 34301 40297 34359 40331
rect 34301 40263 34313 40297
rect 34347 40263 34359 40297
rect 34301 40229 34359 40263
rect 34301 40195 34313 40229
rect 34347 40195 34359 40229
rect 34301 40161 34359 40195
rect 34301 40127 34313 40161
rect 34347 40127 34359 40161
rect 34301 40093 34359 40127
rect 34301 40059 34313 40093
rect 34347 40059 34359 40093
rect 34301 40025 34359 40059
rect 34301 39991 34313 40025
rect 34347 39991 34359 40025
rect 34301 39957 34359 39991
rect 34301 39923 34313 39957
rect 34347 39923 34359 39957
rect 34301 39907 34359 39923
rect 34759 41181 34817 41197
rect 34759 41147 34771 41181
rect 34805 41147 34817 41181
rect 34759 41113 34817 41147
rect 34759 41079 34771 41113
rect 34805 41079 34817 41113
rect 34759 41045 34817 41079
rect 34759 41011 34771 41045
rect 34805 41011 34817 41045
rect 34759 40977 34817 41011
rect 34759 40943 34771 40977
rect 34805 40943 34817 40977
rect 34759 40909 34817 40943
rect 34759 40875 34771 40909
rect 34805 40875 34817 40909
rect 34759 40841 34817 40875
rect 34759 40807 34771 40841
rect 34805 40807 34817 40841
rect 34759 40773 34817 40807
rect 34759 40739 34771 40773
rect 34805 40739 34817 40773
rect 34759 40705 34817 40739
rect 34759 40671 34771 40705
rect 34805 40671 34817 40705
rect 34759 40637 34817 40671
rect 34759 40603 34771 40637
rect 34805 40603 34817 40637
rect 34759 40569 34817 40603
rect 34759 40535 34771 40569
rect 34805 40535 34817 40569
rect 34759 40501 34817 40535
rect 34759 40467 34771 40501
rect 34805 40467 34817 40501
rect 34759 40433 34817 40467
rect 34759 40399 34771 40433
rect 34805 40399 34817 40433
rect 34759 40365 34817 40399
rect 34759 40331 34771 40365
rect 34805 40331 34817 40365
rect 34759 40297 34817 40331
rect 34759 40263 34771 40297
rect 34805 40263 34817 40297
rect 34759 40229 34817 40263
rect 34759 40195 34771 40229
rect 34805 40195 34817 40229
rect 34759 40161 34817 40195
rect 34759 40127 34771 40161
rect 34805 40127 34817 40161
rect 34759 40093 34817 40127
rect 34759 40059 34771 40093
rect 34805 40059 34817 40093
rect 34759 40025 34817 40059
rect 34759 39991 34771 40025
rect 34805 39991 34817 40025
rect 34759 39957 34817 39991
rect 34759 39923 34771 39957
rect 34805 39923 34817 39957
rect 34759 39907 34817 39923
rect 35217 41181 35275 41197
rect 35217 41147 35229 41181
rect 35263 41147 35275 41181
rect 35217 41113 35275 41147
rect 35217 41079 35229 41113
rect 35263 41079 35275 41113
rect 35217 41045 35275 41079
rect 35217 41011 35229 41045
rect 35263 41011 35275 41045
rect 35217 40977 35275 41011
rect 35217 40943 35229 40977
rect 35263 40943 35275 40977
rect 35217 40909 35275 40943
rect 35217 40875 35229 40909
rect 35263 40875 35275 40909
rect 35217 40841 35275 40875
rect 35217 40807 35229 40841
rect 35263 40807 35275 40841
rect 35217 40773 35275 40807
rect 35217 40739 35229 40773
rect 35263 40739 35275 40773
rect 35217 40705 35275 40739
rect 35217 40671 35229 40705
rect 35263 40671 35275 40705
rect 35217 40637 35275 40671
rect 35217 40603 35229 40637
rect 35263 40603 35275 40637
rect 35217 40569 35275 40603
rect 35217 40535 35229 40569
rect 35263 40535 35275 40569
rect 35217 40501 35275 40535
rect 35217 40467 35229 40501
rect 35263 40467 35275 40501
rect 35217 40433 35275 40467
rect 35217 40399 35229 40433
rect 35263 40399 35275 40433
rect 35217 40365 35275 40399
rect 35217 40331 35229 40365
rect 35263 40331 35275 40365
rect 35217 40297 35275 40331
rect 35217 40263 35229 40297
rect 35263 40263 35275 40297
rect 35217 40229 35275 40263
rect 35217 40195 35229 40229
rect 35263 40195 35275 40229
rect 35217 40161 35275 40195
rect 35217 40127 35229 40161
rect 35263 40127 35275 40161
rect 35217 40093 35275 40127
rect 35217 40059 35229 40093
rect 35263 40059 35275 40093
rect 35217 40025 35275 40059
rect 35217 39991 35229 40025
rect 35263 39991 35275 40025
rect 35217 39957 35275 39991
rect 35217 39923 35229 39957
rect 35263 39923 35275 39957
rect 35217 39907 35275 39923
rect 35675 41181 35733 41197
rect 35675 41147 35687 41181
rect 35721 41147 35733 41181
rect 35675 41113 35733 41147
rect 35675 41079 35687 41113
rect 35721 41079 35733 41113
rect 35675 41045 35733 41079
rect 35675 41011 35687 41045
rect 35721 41011 35733 41045
rect 35675 40977 35733 41011
rect 35675 40943 35687 40977
rect 35721 40943 35733 40977
rect 35675 40909 35733 40943
rect 35675 40875 35687 40909
rect 35721 40875 35733 40909
rect 35675 40841 35733 40875
rect 35675 40807 35687 40841
rect 35721 40807 35733 40841
rect 35675 40773 35733 40807
rect 35675 40739 35687 40773
rect 35721 40739 35733 40773
rect 35675 40705 35733 40739
rect 35675 40671 35687 40705
rect 35721 40671 35733 40705
rect 35675 40637 35733 40671
rect 35675 40603 35687 40637
rect 35721 40603 35733 40637
rect 35675 40569 35733 40603
rect 35675 40535 35687 40569
rect 35721 40535 35733 40569
rect 35675 40501 35733 40535
rect 35675 40467 35687 40501
rect 35721 40467 35733 40501
rect 35675 40433 35733 40467
rect 35675 40399 35687 40433
rect 35721 40399 35733 40433
rect 35675 40365 35733 40399
rect 35675 40331 35687 40365
rect 35721 40331 35733 40365
rect 35675 40297 35733 40331
rect 35675 40263 35687 40297
rect 35721 40263 35733 40297
rect 35675 40229 35733 40263
rect 35675 40195 35687 40229
rect 35721 40195 35733 40229
rect 35675 40161 35733 40195
rect 35675 40127 35687 40161
rect 35721 40127 35733 40161
rect 35675 40093 35733 40127
rect 35675 40059 35687 40093
rect 35721 40059 35733 40093
rect 35675 40025 35733 40059
rect 35675 39991 35687 40025
rect 35721 39991 35733 40025
rect 35675 39957 35733 39991
rect 35675 39923 35687 39957
rect 35721 39923 35733 39957
rect 35675 39907 35733 39923
rect 36133 41181 36191 41197
rect 36133 41147 36145 41181
rect 36179 41147 36191 41181
rect 36133 41113 36191 41147
rect 36133 41079 36145 41113
rect 36179 41079 36191 41113
rect 36133 41045 36191 41079
rect 36133 41011 36145 41045
rect 36179 41011 36191 41045
rect 36133 40977 36191 41011
rect 36133 40943 36145 40977
rect 36179 40943 36191 40977
rect 36133 40909 36191 40943
rect 36133 40875 36145 40909
rect 36179 40875 36191 40909
rect 36133 40841 36191 40875
rect 36133 40807 36145 40841
rect 36179 40807 36191 40841
rect 36133 40773 36191 40807
rect 36133 40739 36145 40773
rect 36179 40739 36191 40773
rect 36133 40705 36191 40739
rect 36133 40671 36145 40705
rect 36179 40671 36191 40705
rect 36133 40637 36191 40671
rect 36133 40603 36145 40637
rect 36179 40603 36191 40637
rect 36133 40569 36191 40603
rect 36133 40535 36145 40569
rect 36179 40535 36191 40569
rect 36133 40501 36191 40535
rect 36133 40467 36145 40501
rect 36179 40467 36191 40501
rect 36133 40433 36191 40467
rect 36133 40399 36145 40433
rect 36179 40399 36191 40433
rect 36133 40365 36191 40399
rect 36133 40331 36145 40365
rect 36179 40331 36191 40365
rect 36133 40297 36191 40331
rect 36133 40263 36145 40297
rect 36179 40263 36191 40297
rect 36133 40229 36191 40263
rect 36133 40195 36145 40229
rect 36179 40195 36191 40229
rect 36133 40161 36191 40195
rect 36133 40127 36145 40161
rect 36179 40127 36191 40161
rect 36133 40093 36191 40127
rect 36133 40059 36145 40093
rect 36179 40059 36191 40093
rect 36133 40025 36191 40059
rect 36133 39991 36145 40025
rect 36179 39991 36191 40025
rect 36133 39957 36191 39991
rect 36133 39923 36145 39957
rect 36179 39923 36191 39957
rect 36133 39907 36191 39923
rect 36591 41181 36649 41197
rect 36591 41147 36603 41181
rect 36637 41147 36649 41181
rect 36591 41113 36649 41147
rect 36591 41079 36603 41113
rect 36637 41079 36649 41113
rect 36591 41045 36649 41079
rect 36591 41011 36603 41045
rect 36637 41011 36649 41045
rect 36591 40977 36649 41011
rect 36591 40943 36603 40977
rect 36637 40943 36649 40977
rect 36591 40909 36649 40943
rect 36591 40875 36603 40909
rect 36637 40875 36649 40909
rect 36591 40841 36649 40875
rect 36591 40807 36603 40841
rect 36637 40807 36649 40841
rect 36591 40773 36649 40807
rect 36591 40739 36603 40773
rect 36637 40739 36649 40773
rect 36591 40705 36649 40739
rect 36591 40671 36603 40705
rect 36637 40671 36649 40705
rect 36591 40637 36649 40671
rect 36591 40603 36603 40637
rect 36637 40603 36649 40637
rect 36591 40569 36649 40603
rect 36591 40535 36603 40569
rect 36637 40535 36649 40569
rect 36591 40501 36649 40535
rect 36591 40467 36603 40501
rect 36637 40467 36649 40501
rect 36591 40433 36649 40467
rect 36591 40399 36603 40433
rect 36637 40399 36649 40433
rect 36591 40365 36649 40399
rect 36591 40331 36603 40365
rect 36637 40331 36649 40365
rect 36591 40297 36649 40331
rect 36591 40263 36603 40297
rect 36637 40263 36649 40297
rect 36591 40229 36649 40263
rect 36591 40195 36603 40229
rect 36637 40195 36649 40229
rect 36591 40161 36649 40195
rect 36591 40127 36603 40161
rect 36637 40127 36649 40161
rect 36591 40093 36649 40127
rect 36591 40059 36603 40093
rect 36637 40059 36649 40093
rect 36591 40025 36649 40059
rect 36591 39991 36603 40025
rect 36637 39991 36649 40025
rect 36591 39957 36649 39991
rect 36591 39923 36603 39957
rect 36637 39923 36649 39957
rect 36591 39907 36649 39923
rect 37049 41181 37107 41197
rect 37049 41147 37061 41181
rect 37095 41147 37107 41181
rect 37049 41113 37107 41147
rect 37049 41079 37061 41113
rect 37095 41079 37107 41113
rect 37049 41045 37107 41079
rect 37049 41011 37061 41045
rect 37095 41011 37107 41045
rect 37049 40977 37107 41011
rect 37049 40943 37061 40977
rect 37095 40943 37107 40977
rect 37049 40909 37107 40943
rect 37049 40875 37061 40909
rect 37095 40875 37107 40909
rect 37049 40841 37107 40875
rect 37049 40807 37061 40841
rect 37095 40807 37107 40841
rect 37049 40773 37107 40807
rect 37049 40739 37061 40773
rect 37095 40739 37107 40773
rect 37049 40705 37107 40739
rect 37049 40671 37061 40705
rect 37095 40671 37107 40705
rect 37049 40637 37107 40671
rect 37049 40603 37061 40637
rect 37095 40603 37107 40637
rect 37049 40569 37107 40603
rect 37049 40535 37061 40569
rect 37095 40535 37107 40569
rect 37049 40501 37107 40535
rect 37049 40467 37061 40501
rect 37095 40467 37107 40501
rect 37049 40433 37107 40467
rect 37049 40399 37061 40433
rect 37095 40399 37107 40433
rect 37049 40365 37107 40399
rect 37049 40331 37061 40365
rect 37095 40331 37107 40365
rect 37049 40297 37107 40331
rect 37049 40263 37061 40297
rect 37095 40263 37107 40297
rect 37049 40229 37107 40263
rect 37049 40195 37061 40229
rect 37095 40195 37107 40229
rect 37049 40161 37107 40195
rect 37049 40127 37061 40161
rect 37095 40127 37107 40161
rect 37049 40093 37107 40127
rect 37049 40059 37061 40093
rect 37095 40059 37107 40093
rect 37049 40025 37107 40059
rect 37049 39991 37061 40025
rect 37095 39991 37107 40025
rect 37049 39957 37107 39991
rect 37049 39923 37061 39957
rect 37095 39923 37107 39957
rect 37049 39907 37107 39923
rect 37507 41181 37565 41197
rect 37507 41147 37519 41181
rect 37553 41147 37565 41181
rect 37507 41113 37565 41147
rect 37507 41079 37519 41113
rect 37553 41079 37565 41113
rect 37507 41045 37565 41079
rect 37507 41011 37519 41045
rect 37553 41011 37565 41045
rect 37507 40977 37565 41011
rect 37507 40943 37519 40977
rect 37553 40943 37565 40977
rect 37507 40909 37565 40943
rect 37507 40875 37519 40909
rect 37553 40875 37565 40909
rect 37507 40841 37565 40875
rect 37507 40807 37519 40841
rect 37553 40807 37565 40841
rect 37507 40773 37565 40807
rect 37507 40739 37519 40773
rect 37553 40739 37565 40773
rect 37507 40705 37565 40739
rect 37507 40671 37519 40705
rect 37553 40671 37565 40705
rect 37507 40637 37565 40671
rect 37507 40603 37519 40637
rect 37553 40603 37565 40637
rect 37507 40569 37565 40603
rect 37507 40535 37519 40569
rect 37553 40535 37565 40569
rect 37507 40501 37565 40535
rect 37507 40467 37519 40501
rect 37553 40467 37565 40501
rect 37507 40433 37565 40467
rect 37507 40399 37519 40433
rect 37553 40399 37565 40433
rect 37507 40365 37565 40399
rect 37507 40331 37519 40365
rect 37553 40331 37565 40365
rect 37507 40297 37565 40331
rect 37507 40263 37519 40297
rect 37553 40263 37565 40297
rect 37507 40229 37565 40263
rect 37507 40195 37519 40229
rect 37553 40195 37565 40229
rect 37507 40161 37565 40195
rect 37507 40127 37519 40161
rect 37553 40127 37565 40161
rect 37507 40093 37565 40127
rect 37507 40059 37519 40093
rect 37553 40059 37565 40093
rect 37507 40025 37565 40059
rect 37507 39991 37519 40025
rect 37553 39991 37565 40025
rect 37507 39957 37565 39991
rect 37507 39923 37519 39957
rect 37553 39923 37565 39957
rect 37507 39907 37565 39923
rect 37965 41181 38023 41197
rect 37965 41147 37977 41181
rect 38011 41147 38023 41181
rect 37965 41113 38023 41147
rect 37965 41079 37977 41113
rect 38011 41079 38023 41113
rect 37965 41045 38023 41079
rect 37965 41011 37977 41045
rect 38011 41011 38023 41045
rect 37965 40977 38023 41011
rect 37965 40943 37977 40977
rect 38011 40943 38023 40977
rect 37965 40909 38023 40943
rect 37965 40875 37977 40909
rect 38011 40875 38023 40909
rect 37965 40841 38023 40875
rect 37965 40807 37977 40841
rect 38011 40807 38023 40841
rect 37965 40773 38023 40807
rect 37965 40739 37977 40773
rect 38011 40739 38023 40773
rect 37965 40705 38023 40739
rect 37965 40671 37977 40705
rect 38011 40671 38023 40705
rect 37965 40637 38023 40671
rect 37965 40603 37977 40637
rect 38011 40603 38023 40637
rect 37965 40569 38023 40603
rect 37965 40535 37977 40569
rect 38011 40535 38023 40569
rect 37965 40501 38023 40535
rect 37965 40467 37977 40501
rect 38011 40467 38023 40501
rect 37965 40433 38023 40467
rect 37965 40399 37977 40433
rect 38011 40399 38023 40433
rect 37965 40365 38023 40399
rect 37965 40331 37977 40365
rect 38011 40331 38023 40365
rect 37965 40297 38023 40331
rect 37965 40263 37977 40297
rect 38011 40263 38023 40297
rect 37965 40229 38023 40263
rect 37965 40195 37977 40229
rect 38011 40195 38023 40229
rect 37965 40161 38023 40195
rect 37965 40127 37977 40161
rect 38011 40127 38023 40161
rect 37965 40093 38023 40127
rect 37965 40059 37977 40093
rect 38011 40059 38023 40093
rect 37965 40025 38023 40059
rect 37965 39991 37977 40025
rect 38011 39991 38023 40025
rect 37965 39957 38023 39991
rect 37965 39923 37977 39957
rect 38011 39923 38023 39957
rect 37965 39907 38023 39923
rect 38423 41181 38481 41197
rect 38423 41147 38435 41181
rect 38469 41147 38481 41181
rect 38423 41113 38481 41147
rect 38423 41079 38435 41113
rect 38469 41079 38481 41113
rect 38423 41045 38481 41079
rect 38423 41011 38435 41045
rect 38469 41011 38481 41045
rect 38423 40977 38481 41011
rect 38423 40943 38435 40977
rect 38469 40943 38481 40977
rect 38423 40909 38481 40943
rect 38423 40875 38435 40909
rect 38469 40875 38481 40909
rect 38423 40841 38481 40875
rect 38423 40807 38435 40841
rect 38469 40807 38481 40841
rect 38423 40773 38481 40807
rect 38423 40739 38435 40773
rect 38469 40739 38481 40773
rect 38423 40705 38481 40739
rect 38423 40671 38435 40705
rect 38469 40671 38481 40705
rect 38423 40637 38481 40671
rect 38423 40603 38435 40637
rect 38469 40603 38481 40637
rect 38423 40569 38481 40603
rect 38423 40535 38435 40569
rect 38469 40535 38481 40569
rect 38423 40501 38481 40535
rect 38423 40467 38435 40501
rect 38469 40467 38481 40501
rect 38423 40433 38481 40467
rect 38423 40399 38435 40433
rect 38469 40399 38481 40433
rect 38423 40365 38481 40399
rect 38423 40331 38435 40365
rect 38469 40331 38481 40365
rect 38423 40297 38481 40331
rect 38423 40263 38435 40297
rect 38469 40263 38481 40297
rect 38423 40229 38481 40263
rect 38423 40195 38435 40229
rect 38469 40195 38481 40229
rect 38423 40161 38481 40195
rect 38423 40127 38435 40161
rect 38469 40127 38481 40161
rect 38423 40093 38481 40127
rect 38423 40059 38435 40093
rect 38469 40059 38481 40093
rect 38423 40025 38481 40059
rect 38423 39991 38435 40025
rect 38469 39991 38481 40025
rect 38423 39957 38481 39991
rect 38423 39923 38435 39957
rect 38469 39923 38481 39957
rect 38423 39907 38481 39923
rect 38881 41181 38939 41197
rect 38881 41147 38893 41181
rect 38927 41147 38939 41181
rect 38881 41113 38939 41147
rect 38881 41079 38893 41113
rect 38927 41079 38939 41113
rect 38881 41045 38939 41079
rect 38881 41011 38893 41045
rect 38927 41011 38939 41045
rect 38881 40977 38939 41011
rect 38881 40943 38893 40977
rect 38927 40943 38939 40977
rect 38881 40909 38939 40943
rect 38881 40875 38893 40909
rect 38927 40875 38939 40909
rect 38881 40841 38939 40875
rect 38881 40807 38893 40841
rect 38927 40807 38939 40841
rect 38881 40773 38939 40807
rect 38881 40739 38893 40773
rect 38927 40739 38939 40773
rect 38881 40705 38939 40739
rect 38881 40671 38893 40705
rect 38927 40671 38939 40705
rect 38881 40637 38939 40671
rect 38881 40603 38893 40637
rect 38927 40603 38939 40637
rect 38881 40569 38939 40603
rect 38881 40535 38893 40569
rect 38927 40535 38939 40569
rect 38881 40501 38939 40535
rect 38881 40467 38893 40501
rect 38927 40467 38939 40501
rect 38881 40433 38939 40467
rect 38881 40399 38893 40433
rect 38927 40399 38939 40433
rect 38881 40365 38939 40399
rect 38881 40331 38893 40365
rect 38927 40331 38939 40365
rect 38881 40297 38939 40331
rect 38881 40263 38893 40297
rect 38927 40263 38939 40297
rect 38881 40229 38939 40263
rect 38881 40195 38893 40229
rect 38927 40195 38939 40229
rect 38881 40161 38939 40195
rect 38881 40127 38893 40161
rect 38927 40127 38939 40161
rect 38881 40093 38939 40127
rect 38881 40059 38893 40093
rect 38927 40059 38939 40093
rect 38881 40025 38939 40059
rect 38881 39991 38893 40025
rect 38927 39991 38939 40025
rect 38881 39957 38939 39991
rect 38881 39923 38893 39957
rect 38927 39923 38939 39957
rect 38881 39907 38939 39923
rect 39339 41181 39397 41197
rect 39339 41147 39351 41181
rect 39385 41147 39397 41181
rect 39339 41113 39397 41147
rect 39339 41079 39351 41113
rect 39385 41079 39397 41113
rect 39339 41045 39397 41079
rect 39339 41011 39351 41045
rect 39385 41011 39397 41045
rect 39339 40977 39397 41011
rect 39339 40943 39351 40977
rect 39385 40943 39397 40977
rect 39339 40909 39397 40943
rect 39339 40875 39351 40909
rect 39385 40875 39397 40909
rect 39339 40841 39397 40875
rect 39339 40807 39351 40841
rect 39385 40807 39397 40841
rect 39339 40773 39397 40807
rect 39339 40739 39351 40773
rect 39385 40739 39397 40773
rect 39339 40705 39397 40739
rect 39339 40671 39351 40705
rect 39385 40671 39397 40705
rect 39339 40637 39397 40671
rect 39339 40603 39351 40637
rect 39385 40603 39397 40637
rect 39339 40569 39397 40603
rect 39339 40535 39351 40569
rect 39385 40535 39397 40569
rect 39339 40501 39397 40535
rect 39339 40467 39351 40501
rect 39385 40467 39397 40501
rect 39339 40433 39397 40467
rect 39339 40399 39351 40433
rect 39385 40399 39397 40433
rect 39339 40365 39397 40399
rect 39339 40331 39351 40365
rect 39385 40331 39397 40365
rect 39339 40297 39397 40331
rect 39339 40263 39351 40297
rect 39385 40263 39397 40297
rect 39339 40229 39397 40263
rect 39339 40195 39351 40229
rect 39385 40195 39397 40229
rect 39339 40161 39397 40195
rect 39339 40127 39351 40161
rect 39385 40127 39397 40161
rect 39339 40093 39397 40127
rect 39339 40059 39351 40093
rect 39385 40059 39397 40093
rect 39339 40025 39397 40059
rect 39339 39991 39351 40025
rect 39385 39991 39397 40025
rect 39339 39957 39397 39991
rect 39339 39923 39351 39957
rect 39385 39923 39397 39957
rect 39339 39907 39397 39923
rect 39797 41181 39855 41197
rect 39797 41147 39809 41181
rect 39843 41147 39855 41181
rect 39797 41113 39855 41147
rect 39797 41079 39809 41113
rect 39843 41079 39855 41113
rect 39797 41045 39855 41079
rect 39797 41011 39809 41045
rect 39843 41011 39855 41045
rect 39797 40977 39855 41011
rect 39797 40943 39809 40977
rect 39843 40943 39855 40977
rect 39797 40909 39855 40943
rect 39797 40875 39809 40909
rect 39843 40875 39855 40909
rect 39797 40841 39855 40875
rect 39797 40807 39809 40841
rect 39843 40807 39855 40841
rect 39797 40773 39855 40807
rect 39797 40739 39809 40773
rect 39843 40739 39855 40773
rect 39797 40705 39855 40739
rect 39797 40671 39809 40705
rect 39843 40671 39855 40705
rect 39797 40637 39855 40671
rect 39797 40603 39809 40637
rect 39843 40603 39855 40637
rect 39797 40569 39855 40603
rect 39797 40535 39809 40569
rect 39843 40535 39855 40569
rect 39797 40501 39855 40535
rect 39797 40467 39809 40501
rect 39843 40467 39855 40501
rect 39797 40433 39855 40467
rect 39797 40399 39809 40433
rect 39843 40399 39855 40433
rect 39797 40365 39855 40399
rect 39797 40331 39809 40365
rect 39843 40331 39855 40365
rect 39797 40297 39855 40331
rect 39797 40263 39809 40297
rect 39843 40263 39855 40297
rect 39797 40229 39855 40263
rect 39797 40195 39809 40229
rect 39843 40195 39855 40229
rect 39797 40161 39855 40195
rect 39797 40127 39809 40161
rect 39843 40127 39855 40161
rect 39797 40093 39855 40127
rect 39797 40059 39809 40093
rect 39843 40059 39855 40093
rect 39797 40025 39855 40059
rect 39797 39991 39809 40025
rect 39843 39991 39855 40025
rect 39797 39957 39855 39991
rect 39797 39923 39809 39957
rect 39843 39923 39855 39957
rect 39797 39907 39855 39923
rect 40255 41181 40313 41197
rect 40255 41147 40267 41181
rect 40301 41147 40313 41181
rect 40255 41113 40313 41147
rect 40255 41079 40267 41113
rect 40301 41079 40313 41113
rect 40255 41045 40313 41079
rect 40255 41011 40267 41045
rect 40301 41011 40313 41045
rect 40255 40977 40313 41011
rect 40255 40943 40267 40977
rect 40301 40943 40313 40977
rect 40255 40909 40313 40943
rect 40255 40875 40267 40909
rect 40301 40875 40313 40909
rect 40255 40841 40313 40875
rect 40255 40807 40267 40841
rect 40301 40807 40313 40841
rect 40255 40773 40313 40807
rect 40255 40739 40267 40773
rect 40301 40739 40313 40773
rect 40255 40705 40313 40739
rect 40255 40671 40267 40705
rect 40301 40671 40313 40705
rect 40255 40637 40313 40671
rect 40255 40603 40267 40637
rect 40301 40603 40313 40637
rect 40255 40569 40313 40603
rect 40255 40535 40267 40569
rect 40301 40535 40313 40569
rect 40255 40501 40313 40535
rect 40255 40467 40267 40501
rect 40301 40467 40313 40501
rect 40255 40433 40313 40467
rect 40255 40399 40267 40433
rect 40301 40399 40313 40433
rect 40255 40365 40313 40399
rect 40255 40331 40267 40365
rect 40301 40331 40313 40365
rect 40255 40297 40313 40331
rect 40255 40263 40267 40297
rect 40301 40263 40313 40297
rect 40255 40229 40313 40263
rect 40255 40195 40267 40229
rect 40301 40195 40313 40229
rect 40255 40161 40313 40195
rect 40255 40127 40267 40161
rect 40301 40127 40313 40161
rect 40255 40093 40313 40127
rect 40255 40059 40267 40093
rect 40301 40059 40313 40093
rect 40255 40025 40313 40059
rect 40255 39991 40267 40025
rect 40301 39991 40313 40025
rect 40255 39957 40313 39991
rect 40255 39923 40267 39957
rect 40301 39923 40313 39957
rect 40255 39907 40313 39923
rect 40713 41181 40771 41197
rect 40713 41147 40725 41181
rect 40759 41147 40771 41181
rect 40713 41113 40771 41147
rect 40713 41079 40725 41113
rect 40759 41079 40771 41113
rect 40713 41045 40771 41079
rect 40713 41011 40725 41045
rect 40759 41011 40771 41045
rect 40713 40977 40771 41011
rect 40713 40943 40725 40977
rect 40759 40943 40771 40977
rect 40713 40909 40771 40943
rect 40713 40875 40725 40909
rect 40759 40875 40771 40909
rect 40713 40841 40771 40875
rect 40713 40807 40725 40841
rect 40759 40807 40771 40841
rect 40713 40773 40771 40807
rect 40713 40739 40725 40773
rect 40759 40739 40771 40773
rect 40713 40705 40771 40739
rect 40713 40671 40725 40705
rect 40759 40671 40771 40705
rect 40713 40637 40771 40671
rect 40713 40603 40725 40637
rect 40759 40603 40771 40637
rect 40713 40569 40771 40603
rect 40713 40535 40725 40569
rect 40759 40535 40771 40569
rect 40713 40501 40771 40535
rect 40713 40467 40725 40501
rect 40759 40467 40771 40501
rect 40713 40433 40771 40467
rect 40713 40399 40725 40433
rect 40759 40399 40771 40433
rect 40713 40365 40771 40399
rect 40713 40331 40725 40365
rect 40759 40331 40771 40365
rect 40713 40297 40771 40331
rect 40713 40263 40725 40297
rect 40759 40263 40771 40297
rect 40713 40229 40771 40263
rect 40713 40195 40725 40229
rect 40759 40195 40771 40229
rect 40713 40161 40771 40195
rect 40713 40127 40725 40161
rect 40759 40127 40771 40161
rect 40713 40093 40771 40127
rect 40713 40059 40725 40093
rect 40759 40059 40771 40093
rect 40713 40025 40771 40059
rect 40713 39991 40725 40025
rect 40759 39991 40771 40025
rect 40713 39957 40771 39991
rect 40713 39923 40725 39957
rect 40759 39923 40771 39957
rect 40713 39907 40771 39923
rect 41171 41181 41229 41197
rect 41171 41147 41183 41181
rect 41217 41147 41229 41181
rect 41171 41113 41229 41147
rect 41171 41079 41183 41113
rect 41217 41079 41229 41113
rect 41171 41045 41229 41079
rect 41171 41011 41183 41045
rect 41217 41011 41229 41045
rect 41171 40977 41229 41011
rect 41171 40943 41183 40977
rect 41217 40943 41229 40977
rect 41171 40909 41229 40943
rect 41171 40875 41183 40909
rect 41217 40875 41229 40909
rect 41171 40841 41229 40875
rect 41171 40807 41183 40841
rect 41217 40807 41229 40841
rect 41171 40773 41229 40807
rect 41171 40739 41183 40773
rect 41217 40739 41229 40773
rect 41171 40705 41229 40739
rect 41171 40671 41183 40705
rect 41217 40671 41229 40705
rect 41171 40637 41229 40671
rect 41171 40603 41183 40637
rect 41217 40603 41229 40637
rect 41171 40569 41229 40603
rect 41171 40535 41183 40569
rect 41217 40535 41229 40569
rect 41171 40501 41229 40535
rect 41171 40467 41183 40501
rect 41217 40467 41229 40501
rect 41171 40433 41229 40467
rect 41171 40399 41183 40433
rect 41217 40399 41229 40433
rect 41171 40365 41229 40399
rect 41171 40331 41183 40365
rect 41217 40331 41229 40365
rect 41171 40297 41229 40331
rect 41171 40263 41183 40297
rect 41217 40263 41229 40297
rect 41171 40229 41229 40263
rect 41171 40195 41183 40229
rect 41217 40195 41229 40229
rect 41171 40161 41229 40195
rect 41171 40127 41183 40161
rect 41217 40127 41229 40161
rect 41171 40093 41229 40127
rect 41171 40059 41183 40093
rect 41217 40059 41229 40093
rect 41171 40025 41229 40059
rect 41171 39991 41183 40025
rect 41217 39991 41229 40025
rect 41171 39957 41229 39991
rect 41171 39923 41183 39957
rect 41217 39923 41229 39957
rect 41171 39907 41229 39923
rect 41629 41181 41687 41197
rect 41629 41147 41641 41181
rect 41675 41147 41687 41181
rect 41629 41113 41687 41147
rect 41629 41079 41641 41113
rect 41675 41079 41687 41113
rect 41629 41045 41687 41079
rect 41629 41011 41641 41045
rect 41675 41011 41687 41045
rect 41629 40977 41687 41011
rect 41629 40943 41641 40977
rect 41675 40943 41687 40977
rect 41629 40909 41687 40943
rect 41629 40875 41641 40909
rect 41675 40875 41687 40909
rect 41629 40841 41687 40875
rect 41629 40807 41641 40841
rect 41675 40807 41687 40841
rect 41629 40773 41687 40807
rect 41629 40739 41641 40773
rect 41675 40739 41687 40773
rect 41629 40705 41687 40739
rect 41629 40671 41641 40705
rect 41675 40671 41687 40705
rect 41629 40637 41687 40671
rect 41629 40603 41641 40637
rect 41675 40603 41687 40637
rect 41629 40569 41687 40603
rect 41629 40535 41641 40569
rect 41675 40535 41687 40569
rect 41629 40501 41687 40535
rect 41629 40467 41641 40501
rect 41675 40467 41687 40501
rect 41629 40433 41687 40467
rect 41629 40399 41641 40433
rect 41675 40399 41687 40433
rect 41629 40365 41687 40399
rect 41629 40331 41641 40365
rect 41675 40331 41687 40365
rect 41629 40297 41687 40331
rect 41629 40263 41641 40297
rect 41675 40263 41687 40297
rect 41629 40229 41687 40263
rect 41629 40195 41641 40229
rect 41675 40195 41687 40229
rect 41629 40161 41687 40195
rect 41629 40127 41641 40161
rect 41675 40127 41687 40161
rect 41629 40093 41687 40127
rect 41629 40059 41641 40093
rect 41675 40059 41687 40093
rect 41629 40025 41687 40059
rect 41629 39991 41641 40025
rect 41675 39991 41687 40025
rect 41629 39957 41687 39991
rect 41629 39923 41641 39957
rect 41675 39923 41687 39957
rect 41629 39907 41687 39923
rect 42087 41181 42145 41197
rect 42087 41147 42099 41181
rect 42133 41147 42145 41181
rect 42087 41113 42145 41147
rect 42087 41079 42099 41113
rect 42133 41079 42145 41113
rect 42087 41045 42145 41079
rect 42087 41011 42099 41045
rect 42133 41011 42145 41045
rect 42087 40977 42145 41011
rect 42087 40943 42099 40977
rect 42133 40943 42145 40977
rect 42087 40909 42145 40943
rect 42087 40875 42099 40909
rect 42133 40875 42145 40909
rect 42087 40841 42145 40875
rect 42087 40807 42099 40841
rect 42133 40807 42145 40841
rect 42087 40773 42145 40807
rect 42087 40739 42099 40773
rect 42133 40739 42145 40773
rect 42087 40705 42145 40739
rect 42087 40671 42099 40705
rect 42133 40671 42145 40705
rect 42087 40637 42145 40671
rect 42087 40603 42099 40637
rect 42133 40603 42145 40637
rect 42087 40569 42145 40603
rect 42087 40535 42099 40569
rect 42133 40535 42145 40569
rect 42087 40501 42145 40535
rect 42087 40467 42099 40501
rect 42133 40467 42145 40501
rect 42087 40433 42145 40467
rect 42087 40399 42099 40433
rect 42133 40399 42145 40433
rect 42087 40365 42145 40399
rect 42087 40331 42099 40365
rect 42133 40331 42145 40365
rect 42087 40297 42145 40331
rect 42087 40263 42099 40297
rect 42133 40263 42145 40297
rect 42087 40229 42145 40263
rect 42087 40195 42099 40229
rect 42133 40195 42145 40229
rect 42087 40161 42145 40195
rect 42087 40127 42099 40161
rect 42133 40127 42145 40161
rect 42087 40093 42145 40127
rect 42087 40059 42099 40093
rect 42133 40059 42145 40093
rect 42087 40025 42145 40059
rect 42087 39991 42099 40025
rect 42133 39991 42145 40025
rect 42087 39957 42145 39991
rect 42087 39923 42099 39957
rect 42133 39923 42145 39957
rect 42087 39907 42145 39923
rect 42545 41181 42603 41197
rect 42545 41147 42557 41181
rect 42591 41147 42603 41181
rect 42545 41113 42603 41147
rect 42545 41079 42557 41113
rect 42591 41079 42603 41113
rect 42545 41045 42603 41079
rect 42545 41011 42557 41045
rect 42591 41011 42603 41045
rect 42545 40977 42603 41011
rect 42545 40943 42557 40977
rect 42591 40943 42603 40977
rect 42545 40909 42603 40943
rect 42545 40875 42557 40909
rect 42591 40875 42603 40909
rect 42545 40841 42603 40875
rect 42545 40807 42557 40841
rect 42591 40807 42603 40841
rect 42545 40773 42603 40807
rect 42545 40739 42557 40773
rect 42591 40739 42603 40773
rect 42545 40705 42603 40739
rect 42545 40671 42557 40705
rect 42591 40671 42603 40705
rect 42545 40637 42603 40671
rect 42545 40603 42557 40637
rect 42591 40603 42603 40637
rect 42545 40569 42603 40603
rect 42545 40535 42557 40569
rect 42591 40535 42603 40569
rect 42545 40501 42603 40535
rect 42545 40467 42557 40501
rect 42591 40467 42603 40501
rect 42545 40433 42603 40467
rect 42545 40399 42557 40433
rect 42591 40399 42603 40433
rect 42545 40365 42603 40399
rect 42545 40331 42557 40365
rect 42591 40331 42603 40365
rect 42545 40297 42603 40331
rect 42545 40263 42557 40297
rect 42591 40263 42603 40297
rect 42545 40229 42603 40263
rect 42545 40195 42557 40229
rect 42591 40195 42603 40229
rect 42545 40161 42603 40195
rect 42545 40127 42557 40161
rect 42591 40127 42603 40161
rect 42545 40093 42603 40127
rect 42545 40059 42557 40093
rect 42591 40059 42603 40093
rect 42545 40025 42603 40059
rect 42545 39991 42557 40025
rect 42591 39991 42603 40025
rect 42545 39957 42603 39991
rect 42545 39923 42557 39957
rect 42591 39923 42603 39957
rect 42545 39907 42603 39923
rect 30354 37020 31034 37072
rect 30354 36986 30408 37020
rect 30442 36986 30498 37020
rect 30532 36986 30588 37020
rect 30622 36986 30678 37020
rect 30712 36986 30768 37020
rect 30802 36986 30858 37020
rect 30892 36986 30948 37020
rect 30982 36986 31034 37020
rect 30354 36930 31034 36986
rect 30354 36896 30408 36930
rect 30442 36896 30498 36930
rect 30532 36896 30588 36930
rect 30622 36896 30678 36930
rect 30712 36896 30768 36930
rect 30802 36896 30858 36930
rect 30892 36896 30948 36930
rect 30982 36896 31034 36930
rect 30354 36840 31034 36896
rect 30354 36806 30408 36840
rect 30442 36806 30498 36840
rect 30532 36806 30588 36840
rect 30622 36806 30678 36840
rect 30712 36806 30768 36840
rect 30802 36806 30858 36840
rect 30892 36806 30948 36840
rect 30982 36806 31034 36840
rect 30354 36750 31034 36806
rect 30354 36716 30408 36750
rect 30442 36716 30498 36750
rect 30532 36716 30588 36750
rect 30622 36716 30678 36750
rect 30712 36716 30768 36750
rect 30802 36716 30858 36750
rect 30892 36716 30948 36750
rect 30982 36716 31034 36750
rect 30354 36660 31034 36716
rect 30354 36626 30408 36660
rect 30442 36626 30498 36660
rect 30532 36626 30588 36660
rect 30622 36626 30678 36660
rect 30712 36626 30768 36660
rect 30802 36626 30858 36660
rect 30892 36626 30948 36660
rect 30982 36626 31034 36660
rect 30354 36570 31034 36626
rect 30354 36536 30408 36570
rect 30442 36536 30498 36570
rect 30532 36536 30588 36570
rect 30622 36536 30678 36570
rect 30712 36536 30768 36570
rect 30802 36536 30858 36570
rect 30892 36536 30948 36570
rect 30982 36536 31034 36570
rect 30354 36480 31034 36536
rect 30354 36446 30408 36480
rect 30442 36446 30498 36480
rect 30532 36446 30588 36480
rect 30622 36446 30678 36480
rect 30712 36446 30768 36480
rect 30802 36446 30858 36480
rect 30892 36446 30948 36480
rect 30982 36446 31034 36480
rect 30354 36392 31034 36446
rect 31694 37020 32374 37072
rect 31694 36986 31748 37020
rect 31782 36986 31838 37020
rect 31872 36986 31928 37020
rect 31962 36986 32018 37020
rect 32052 36986 32108 37020
rect 32142 36986 32198 37020
rect 32232 36986 32288 37020
rect 32322 36986 32374 37020
rect 31694 36930 32374 36986
rect 31694 36896 31748 36930
rect 31782 36896 31838 36930
rect 31872 36896 31928 36930
rect 31962 36896 32018 36930
rect 32052 36896 32108 36930
rect 32142 36896 32198 36930
rect 32232 36896 32288 36930
rect 32322 36896 32374 36930
rect 31694 36840 32374 36896
rect 31694 36806 31748 36840
rect 31782 36806 31838 36840
rect 31872 36806 31928 36840
rect 31962 36806 32018 36840
rect 32052 36806 32108 36840
rect 32142 36806 32198 36840
rect 32232 36806 32288 36840
rect 32322 36806 32374 36840
rect 31694 36750 32374 36806
rect 31694 36716 31748 36750
rect 31782 36716 31838 36750
rect 31872 36716 31928 36750
rect 31962 36716 32018 36750
rect 32052 36716 32108 36750
rect 32142 36716 32198 36750
rect 32232 36716 32288 36750
rect 32322 36716 32374 36750
rect 31694 36660 32374 36716
rect 31694 36626 31748 36660
rect 31782 36626 31838 36660
rect 31872 36626 31928 36660
rect 31962 36626 32018 36660
rect 32052 36626 32108 36660
rect 32142 36626 32198 36660
rect 32232 36626 32288 36660
rect 32322 36626 32374 36660
rect 31694 36570 32374 36626
rect 31694 36536 31748 36570
rect 31782 36536 31838 36570
rect 31872 36536 31928 36570
rect 31962 36536 32018 36570
rect 32052 36536 32108 36570
rect 32142 36536 32198 36570
rect 32232 36536 32288 36570
rect 32322 36536 32374 36570
rect 31694 36480 32374 36536
rect 31694 36446 31748 36480
rect 31782 36446 31838 36480
rect 31872 36446 31928 36480
rect 31962 36446 32018 36480
rect 32052 36446 32108 36480
rect 32142 36446 32198 36480
rect 32232 36446 32288 36480
rect 32322 36446 32374 36480
rect 31694 36392 32374 36446
rect 33034 37020 33714 37072
rect 33034 36986 33088 37020
rect 33122 36986 33178 37020
rect 33212 36986 33268 37020
rect 33302 36986 33358 37020
rect 33392 36986 33448 37020
rect 33482 36986 33538 37020
rect 33572 36986 33628 37020
rect 33662 36986 33714 37020
rect 33034 36930 33714 36986
rect 33034 36896 33088 36930
rect 33122 36896 33178 36930
rect 33212 36896 33268 36930
rect 33302 36896 33358 36930
rect 33392 36896 33448 36930
rect 33482 36896 33538 36930
rect 33572 36896 33628 36930
rect 33662 36896 33714 36930
rect 33034 36840 33714 36896
rect 33034 36806 33088 36840
rect 33122 36806 33178 36840
rect 33212 36806 33268 36840
rect 33302 36806 33358 36840
rect 33392 36806 33448 36840
rect 33482 36806 33538 36840
rect 33572 36806 33628 36840
rect 33662 36806 33714 36840
rect 33034 36750 33714 36806
rect 33034 36716 33088 36750
rect 33122 36716 33178 36750
rect 33212 36716 33268 36750
rect 33302 36716 33358 36750
rect 33392 36716 33448 36750
rect 33482 36716 33538 36750
rect 33572 36716 33628 36750
rect 33662 36716 33714 36750
rect 33034 36660 33714 36716
rect 33034 36626 33088 36660
rect 33122 36626 33178 36660
rect 33212 36626 33268 36660
rect 33302 36626 33358 36660
rect 33392 36626 33448 36660
rect 33482 36626 33538 36660
rect 33572 36626 33628 36660
rect 33662 36626 33714 36660
rect 33034 36570 33714 36626
rect 33034 36536 33088 36570
rect 33122 36536 33178 36570
rect 33212 36536 33268 36570
rect 33302 36536 33358 36570
rect 33392 36536 33448 36570
rect 33482 36536 33538 36570
rect 33572 36536 33628 36570
rect 33662 36536 33714 36570
rect 33034 36480 33714 36536
rect 33034 36446 33088 36480
rect 33122 36446 33178 36480
rect 33212 36446 33268 36480
rect 33302 36446 33358 36480
rect 33392 36446 33448 36480
rect 33482 36446 33538 36480
rect 33572 36446 33628 36480
rect 33662 36446 33714 36480
rect 33034 36392 33714 36446
rect 34374 37020 35054 37072
rect 34374 36986 34428 37020
rect 34462 36986 34518 37020
rect 34552 36986 34608 37020
rect 34642 36986 34698 37020
rect 34732 36986 34788 37020
rect 34822 36986 34878 37020
rect 34912 36986 34968 37020
rect 35002 36986 35054 37020
rect 34374 36930 35054 36986
rect 34374 36896 34428 36930
rect 34462 36896 34518 36930
rect 34552 36896 34608 36930
rect 34642 36896 34698 36930
rect 34732 36896 34788 36930
rect 34822 36896 34878 36930
rect 34912 36896 34968 36930
rect 35002 36896 35054 36930
rect 34374 36840 35054 36896
rect 34374 36806 34428 36840
rect 34462 36806 34518 36840
rect 34552 36806 34608 36840
rect 34642 36806 34698 36840
rect 34732 36806 34788 36840
rect 34822 36806 34878 36840
rect 34912 36806 34968 36840
rect 35002 36806 35054 36840
rect 34374 36750 35054 36806
rect 34374 36716 34428 36750
rect 34462 36716 34518 36750
rect 34552 36716 34608 36750
rect 34642 36716 34698 36750
rect 34732 36716 34788 36750
rect 34822 36716 34878 36750
rect 34912 36716 34968 36750
rect 35002 36716 35054 36750
rect 34374 36660 35054 36716
rect 34374 36626 34428 36660
rect 34462 36626 34518 36660
rect 34552 36626 34608 36660
rect 34642 36626 34698 36660
rect 34732 36626 34788 36660
rect 34822 36626 34878 36660
rect 34912 36626 34968 36660
rect 35002 36626 35054 36660
rect 34374 36570 35054 36626
rect 34374 36536 34428 36570
rect 34462 36536 34518 36570
rect 34552 36536 34608 36570
rect 34642 36536 34698 36570
rect 34732 36536 34788 36570
rect 34822 36536 34878 36570
rect 34912 36536 34968 36570
rect 35002 36536 35054 36570
rect 34374 36480 35054 36536
rect 34374 36446 34428 36480
rect 34462 36446 34518 36480
rect 34552 36446 34608 36480
rect 34642 36446 34698 36480
rect 34732 36446 34788 36480
rect 34822 36446 34878 36480
rect 34912 36446 34968 36480
rect 35002 36446 35054 36480
rect 34374 36392 35054 36446
rect 35714 37020 36394 37072
rect 35714 36986 35768 37020
rect 35802 36986 35858 37020
rect 35892 36986 35948 37020
rect 35982 36986 36038 37020
rect 36072 36986 36128 37020
rect 36162 36986 36218 37020
rect 36252 36986 36308 37020
rect 36342 36986 36394 37020
rect 35714 36930 36394 36986
rect 35714 36896 35768 36930
rect 35802 36896 35858 36930
rect 35892 36896 35948 36930
rect 35982 36896 36038 36930
rect 36072 36896 36128 36930
rect 36162 36896 36218 36930
rect 36252 36896 36308 36930
rect 36342 36896 36394 36930
rect 35714 36840 36394 36896
rect 35714 36806 35768 36840
rect 35802 36806 35858 36840
rect 35892 36806 35948 36840
rect 35982 36806 36038 36840
rect 36072 36806 36128 36840
rect 36162 36806 36218 36840
rect 36252 36806 36308 36840
rect 36342 36806 36394 36840
rect 35714 36750 36394 36806
rect 35714 36716 35768 36750
rect 35802 36716 35858 36750
rect 35892 36716 35948 36750
rect 35982 36716 36038 36750
rect 36072 36716 36128 36750
rect 36162 36716 36218 36750
rect 36252 36716 36308 36750
rect 36342 36716 36394 36750
rect 35714 36660 36394 36716
rect 35714 36626 35768 36660
rect 35802 36626 35858 36660
rect 35892 36626 35948 36660
rect 35982 36626 36038 36660
rect 36072 36626 36128 36660
rect 36162 36626 36218 36660
rect 36252 36626 36308 36660
rect 36342 36626 36394 36660
rect 35714 36570 36394 36626
rect 35714 36536 35768 36570
rect 35802 36536 35858 36570
rect 35892 36536 35948 36570
rect 35982 36536 36038 36570
rect 36072 36536 36128 36570
rect 36162 36536 36218 36570
rect 36252 36536 36308 36570
rect 36342 36536 36394 36570
rect 35714 36480 36394 36536
rect 35714 36446 35768 36480
rect 35802 36446 35858 36480
rect 35892 36446 35948 36480
rect 35982 36446 36038 36480
rect 36072 36446 36128 36480
rect 36162 36446 36218 36480
rect 36252 36446 36308 36480
rect 36342 36446 36394 36480
rect 35714 36392 36394 36446
rect 37054 37020 37734 37072
rect 37054 36986 37108 37020
rect 37142 36986 37198 37020
rect 37232 36986 37288 37020
rect 37322 36986 37378 37020
rect 37412 36986 37468 37020
rect 37502 36986 37558 37020
rect 37592 36986 37648 37020
rect 37682 36986 37734 37020
rect 37054 36930 37734 36986
rect 37054 36896 37108 36930
rect 37142 36896 37198 36930
rect 37232 36896 37288 36930
rect 37322 36896 37378 36930
rect 37412 36896 37468 36930
rect 37502 36896 37558 36930
rect 37592 36896 37648 36930
rect 37682 36896 37734 36930
rect 37054 36840 37734 36896
rect 37054 36806 37108 36840
rect 37142 36806 37198 36840
rect 37232 36806 37288 36840
rect 37322 36806 37378 36840
rect 37412 36806 37468 36840
rect 37502 36806 37558 36840
rect 37592 36806 37648 36840
rect 37682 36806 37734 36840
rect 37054 36750 37734 36806
rect 37054 36716 37108 36750
rect 37142 36716 37198 36750
rect 37232 36716 37288 36750
rect 37322 36716 37378 36750
rect 37412 36716 37468 36750
rect 37502 36716 37558 36750
rect 37592 36716 37648 36750
rect 37682 36716 37734 36750
rect 37054 36660 37734 36716
rect 37054 36626 37108 36660
rect 37142 36626 37198 36660
rect 37232 36626 37288 36660
rect 37322 36626 37378 36660
rect 37412 36626 37468 36660
rect 37502 36626 37558 36660
rect 37592 36626 37648 36660
rect 37682 36626 37734 36660
rect 37054 36570 37734 36626
rect 37054 36536 37108 36570
rect 37142 36536 37198 36570
rect 37232 36536 37288 36570
rect 37322 36536 37378 36570
rect 37412 36536 37468 36570
rect 37502 36536 37558 36570
rect 37592 36536 37648 36570
rect 37682 36536 37734 36570
rect 37054 36480 37734 36536
rect 37054 36446 37108 36480
rect 37142 36446 37198 36480
rect 37232 36446 37288 36480
rect 37322 36446 37378 36480
rect 37412 36446 37468 36480
rect 37502 36446 37558 36480
rect 37592 36446 37648 36480
rect 37682 36446 37734 36480
rect 37054 36392 37734 36446
rect 38394 37020 39074 37072
rect 38394 36986 38448 37020
rect 38482 36986 38538 37020
rect 38572 36986 38628 37020
rect 38662 36986 38718 37020
rect 38752 36986 38808 37020
rect 38842 36986 38898 37020
rect 38932 36986 38988 37020
rect 39022 36986 39074 37020
rect 38394 36930 39074 36986
rect 38394 36896 38448 36930
rect 38482 36896 38538 36930
rect 38572 36896 38628 36930
rect 38662 36896 38718 36930
rect 38752 36896 38808 36930
rect 38842 36896 38898 36930
rect 38932 36896 38988 36930
rect 39022 36896 39074 36930
rect 38394 36840 39074 36896
rect 38394 36806 38448 36840
rect 38482 36806 38538 36840
rect 38572 36806 38628 36840
rect 38662 36806 38718 36840
rect 38752 36806 38808 36840
rect 38842 36806 38898 36840
rect 38932 36806 38988 36840
rect 39022 36806 39074 36840
rect 38394 36750 39074 36806
rect 38394 36716 38448 36750
rect 38482 36716 38538 36750
rect 38572 36716 38628 36750
rect 38662 36716 38718 36750
rect 38752 36716 38808 36750
rect 38842 36716 38898 36750
rect 38932 36716 38988 36750
rect 39022 36716 39074 36750
rect 38394 36660 39074 36716
rect 38394 36626 38448 36660
rect 38482 36626 38538 36660
rect 38572 36626 38628 36660
rect 38662 36626 38718 36660
rect 38752 36626 38808 36660
rect 38842 36626 38898 36660
rect 38932 36626 38988 36660
rect 39022 36626 39074 36660
rect 38394 36570 39074 36626
rect 38394 36536 38448 36570
rect 38482 36536 38538 36570
rect 38572 36536 38628 36570
rect 38662 36536 38718 36570
rect 38752 36536 38808 36570
rect 38842 36536 38898 36570
rect 38932 36536 38988 36570
rect 39022 36536 39074 36570
rect 38394 36480 39074 36536
rect 38394 36446 38448 36480
rect 38482 36446 38538 36480
rect 38572 36446 38628 36480
rect 38662 36446 38718 36480
rect 38752 36446 38808 36480
rect 38842 36446 38898 36480
rect 38932 36446 38988 36480
rect 39022 36446 39074 36480
rect 38394 36392 39074 36446
rect 14183 33661 14241 33677
rect 14183 33627 14195 33661
rect 14229 33627 14241 33661
rect 14183 33593 14241 33627
rect 14183 33559 14195 33593
rect 14229 33559 14241 33593
rect 14183 33525 14241 33559
rect 14183 33491 14195 33525
rect 14229 33491 14241 33525
rect 14183 33457 14241 33491
rect 14183 33423 14195 33457
rect 14229 33423 14241 33457
rect 14183 33389 14241 33423
rect 14183 33355 14195 33389
rect 14229 33355 14241 33389
rect 14183 33321 14241 33355
rect 14183 33287 14195 33321
rect 14229 33287 14241 33321
rect 14183 33253 14241 33287
rect 14183 33219 14195 33253
rect 14229 33219 14241 33253
rect 14183 33185 14241 33219
rect 14183 33151 14195 33185
rect 14229 33151 14241 33185
rect 14183 33117 14241 33151
rect 14183 33083 14195 33117
rect 14229 33083 14241 33117
rect 14183 33049 14241 33083
rect 14183 33015 14195 33049
rect 14229 33015 14241 33049
rect 14183 32981 14241 33015
rect 14183 32947 14195 32981
rect 14229 32947 14241 32981
rect 14183 32913 14241 32947
rect 14183 32879 14195 32913
rect 14229 32879 14241 32913
rect 14183 32845 14241 32879
rect 14183 32811 14195 32845
rect 14229 32811 14241 32845
rect 14183 32777 14241 32811
rect 14183 32743 14195 32777
rect 14229 32743 14241 32777
rect 14183 32709 14241 32743
rect 14183 32675 14195 32709
rect 14229 32675 14241 32709
rect 14183 32641 14241 32675
rect 14183 32607 14195 32641
rect 14229 32607 14241 32641
rect 14183 32573 14241 32607
rect 14183 32539 14195 32573
rect 14229 32539 14241 32573
rect 14183 32505 14241 32539
rect 14183 32471 14195 32505
rect 14229 32471 14241 32505
rect 14183 32437 14241 32471
rect 14183 32403 14195 32437
rect 14229 32403 14241 32437
rect 14183 32387 14241 32403
rect 14641 33661 14699 33677
rect 14641 33627 14653 33661
rect 14687 33627 14699 33661
rect 14641 33593 14699 33627
rect 14641 33559 14653 33593
rect 14687 33559 14699 33593
rect 14641 33525 14699 33559
rect 14641 33491 14653 33525
rect 14687 33491 14699 33525
rect 14641 33457 14699 33491
rect 14641 33423 14653 33457
rect 14687 33423 14699 33457
rect 14641 33389 14699 33423
rect 14641 33355 14653 33389
rect 14687 33355 14699 33389
rect 14641 33321 14699 33355
rect 14641 33287 14653 33321
rect 14687 33287 14699 33321
rect 14641 33253 14699 33287
rect 14641 33219 14653 33253
rect 14687 33219 14699 33253
rect 14641 33185 14699 33219
rect 14641 33151 14653 33185
rect 14687 33151 14699 33185
rect 14641 33117 14699 33151
rect 14641 33083 14653 33117
rect 14687 33083 14699 33117
rect 14641 33049 14699 33083
rect 14641 33015 14653 33049
rect 14687 33015 14699 33049
rect 14641 32981 14699 33015
rect 14641 32947 14653 32981
rect 14687 32947 14699 32981
rect 14641 32913 14699 32947
rect 14641 32879 14653 32913
rect 14687 32879 14699 32913
rect 14641 32845 14699 32879
rect 14641 32811 14653 32845
rect 14687 32811 14699 32845
rect 14641 32777 14699 32811
rect 14641 32743 14653 32777
rect 14687 32743 14699 32777
rect 14641 32709 14699 32743
rect 14641 32675 14653 32709
rect 14687 32675 14699 32709
rect 14641 32641 14699 32675
rect 14641 32607 14653 32641
rect 14687 32607 14699 32641
rect 14641 32573 14699 32607
rect 14641 32539 14653 32573
rect 14687 32539 14699 32573
rect 14641 32505 14699 32539
rect 14641 32471 14653 32505
rect 14687 32471 14699 32505
rect 14641 32437 14699 32471
rect 14641 32403 14653 32437
rect 14687 32403 14699 32437
rect 14641 32387 14699 32403
rect 15099 33661 15157 33677
rect 15099 33627 15111 33661
rect 15145 33627 15157 33661
rect 15099 33593 15157 33627
rect 15099 33559 15111 33593
rect 15145 33559 15157 33593
rect 15099 33525 15157 33559
rect 15099 33491 15111 33525
rect 15145 33491 15157 33525
rect 15099 33457 15157 33491
rect 15099 33423 15111 33457
rect 15145 33423 15157 33457
rect 15099 33389 15157 33423
rect 15099 33355 15111 33389
rect 15145 33355 15157 33389
rect 15099 33321 15157 33355
rect 15099 33287 15111 33321
rect 15145 33287 15157 33321
rect 15099 33253 15157 33287
rect 15099 33219 15111 33253
rect 15145 33219 15157 33253
rect 15099 33185 15157 33219
rect 15099 33151 15111 33185
rect 15145 33151 15157 33185
rect 15099 33117 15157 33151
rect 15099 33083 15111 33117
rect 15145 33083 15157 33117
rect 15099 33049 15157 33083
rect 15099 33015 15111 33049
rect 15145 33015 15157 33049
rect 15099 32981 15157 33015
rect 15099 32947 15111 32981
rect 15145 32947 15157 32981
rect 15099 32913 15157 32947
rect 15099 32879 15111 32913
rect 15145 32879 15157 32913
rect 15099 32845 15157 32879
rect 15099 32811 15111 32845
rect 15145 32811 15157 32845
rect 15099 32777 15157 32811
rect 15099 32743 15111 32777
rect 15145 32743 15157 32777
rect 15099 32709 15157 32743
rect 15099 32675 15111 32709
rect 15145 32675 15157 32709
rect 15099 32641 15157 32675
rect 15099 32607 15111 32641
rect 15145 32607 15157 32641
rect 15099 32573 15157 32607
rect 15099 32539 15111 32573
rect 15145 32539 15157 32573
rect 15099 32505 15157 32539
rect 15099 32471 15111 32505
rect 15145 32471 15157 32505
rect 15099 32437 15157 32471
rect 15099 32403 15111 32437
rect 15145 32403 15157 32437
rect 15099 32387 15157 32403
rect 15557 33661 15615 33677
rect 15557 33627 15569 33661
rect 15603 33627 15615 33661
rect 15557 33593 15615 33627
rect 15557 33559 15569 33593
rect 15603 33559 15615 33593
rect 15557 33525 15615 33559
rect 15557 33491 15569 33525
rect 15603 33491 15615 33525
rect 15557 33457 15615 33491
rect 15557 33423 15569 33457
rect 15603 33423 15615 33457
rect 15557 33389 15615 33423
rect 15557 33355 15569 33389
rect 15603 33355 15615 33389
rect 15557 33321 15615 33355
rect 15557 33287 15569 33321
rect 15603 33287 15615 33321
rect 15557 33253 15615 33287
rect 15557 33219 15569 33253
rect 15603 33219 15615 33253
rect 15557 33185 15615 33219
rect 15557 33151 15569 33185
rect 15603 33151 15615 33185
rect 15557 33117 15615 33151
rect 15557 33083 15569 33117
rect 15603 33083 15615 33117
rect 15557 33049 15615 33083
rect 15557 33015 15569 33049
rect 15603 33015 15615 33049
rect 15557 32981 15615 33015
rect 15557 32947 15569 32981
rect 15603 32947 15615 32981
rect 15557 32913 15615 32947
rect 15557 32879 15569 32913
rect 15603 32879 15615 32913
rect 15557 32845 15615 32879
rect 15557 32811 15569 32845
rect 15603 32811 15615 32845
rect 15557 32777 15615 32811
rect 15557 32743 15569 32777
rect 15603 32743 15615 32777
rect 15557 32709 15615 32743
rect 15557 32675 15569 32709
rect 15603 32675 15615 32709
rect 15557 32641 15615 32675
rect 15557 32607 15569 32641
rect 15603 32607 15615 32641
rect 15557 32573 15615 32607
rect 15557 32539 15569 32573
rect 15603 32539 15615 32573
rect 15557 32505 15615 32539
rect 15557 32471 15569 32505
rect 15603 32471 15615 32505
rect 15557 32437 15615 32471
rect 15557 32403 15569 32437
rect 15603 32403 15615 32437
rect 15557 32387 15615 32403
rect 16015 33661 16073 33677
rect 16015 33627 16027 33661
rect 16061 33627 16073 33661
rect 16015 33593 16073 33627
rect 16015 33559 16027 33593
rect 16061 33559 16073 33593
rect 16015 33525 16073 33559
rect 16015 33491 16027 33525
rect 16061 33491 16073 33525
rect 16015 33457 16073 33491
rect 16015 33423 16027 33457
rect 16061 33423 16073 33457
rect 16015 33389 16073 33423
rect 16015 33355 16027 33389
rect 16061 33355 16073 33389
rect 16015 33321 16073 33355
rect 16015 33287 16027 33321
rect 16061 33287 16073 33321
rect 16015 33253 16073 33287
rect 16015 33219 16027 33253
rect 16061 33219 16073 33253
rect 16015 33185 16073 33219
rect 16015 33151 16027 33185
rect 16061 33151 16073 33185
rect 16015 33117 16073 33151
rect 16015 33083 16027 33117
rect 16061 33083 16073 33117
rect 16015 33049 16073 33083
rect 16015 33015 16027 33049
rect 16061 33015 16073 33049
rect 16015 32981 16073 33015
rect 16015 32947 16027 32981
rect 16061 32947 16073 32981
rect 16015 32913 16073 32947
rect 16015 32879 16027 32913
rect 16061 32879 16073 32913
rect 16015 32845 16073 32879
rect 16015 32811 16027 32845
rect 16061 32811 16073 32845
rect 16015 32777 16073 32811
rect 16015 32743 16027 32777
rect 16061 32743 16073 32777
rect 16015 32709 16073 32743
rect 16015 32675 16027 32709
rect 16061 32675 16073 32709
rect 16015 32641 16073 32675
rect 16015 32607 16027 32641
rect 16061 32607 16073 32641
rect 16015 32573 16073 32607
rect 16015 32539 16027 32573
rect 16061 32539 16073 32573
rect 16015 32505 16073 32539
rect 16015 32471 16027 32505
rect 16061 32471 16073 32505
rect 16015 32437 16073 32471
rect 16015 32403 16027 32437
rect 16061 32403 16073 32437
rect 16015 32387 16073 32403
rect 16473 33661 16531 33677
rect 16473 33627 16485 33661
rect 16519 33627 16531 33661
rect 16473 33593 16531 33627
rect 16473 33559 16485 33593
rect 16519 33559 16531 33593
rect 16473 33525 16531 33559
rect 16473 33491 16485 33525
rect 16519 33491 16531 33525
rect 16473 33457 16531 33491
rect 16473 33423 16485 33457
rect 16519 33423 16531 33457
rect 16473 33389 16531 33423
rect 16473 33355 16485 33389
rect 16519 33355 16531 33389
rect 16473 33321 16531 33355
rect 16473 33287 16485 33321
rect 16519 33287 16531 33321
rect 16473 33253 16531 33287
rect 16473 33219 16485 33253
rect 16519 33219 16531 33253
rect 16473 33185 16531 33219
rect 16473 33151 16485 33185
rect 16519 33151 16531 33185
rect 16473 33117 16531 33151
rect 16473 33083 16485 33117
rect 16519 33083 16531 33117
rect 16473 33049 16531 33083
rect 16473 33015 16485 33049
rect 16519 33015 16531 33049
rect 16473 32981 16531 33015
rect 16473 32947 16485 32981
rect 16519 32947 16531 32981
rect 16473 32913 16531 32947
rect 16473 32879 16485 32913
rect 16519 32879 16531 32913
rect 16473 32845 16531 32879
rect 16473 32811 16485 32845
rect 16519 32811 16531 32845
rect 16473 32777 16531 32811
rect 16473 32743 16485 32777
rect 16519 32743 16531 32777
rect 16473 32709 16531 32743
rect 16473 32675 16485 32709
rect 16519 32675 16531 32709
rect 16473 32641 16531 32675
rect 16473 32607 16485 32641
rect 16519 32607 16531 32641
rect 16473 32573 16531 32607
rect 16473 32539 16485 32573
rect 16519 32539 16531 32573
rect 16473 32505 16531 32539
rect 16473 32471 16485 32505
rect 16519 32471 16531 32505
rect 16473 32437 16531 32471
rect 16473 32403 16485 32437
rect 16519 32403 16531 32437
rect 16473 32387 16531 32403
rect 16931 33661 16989 33677
rect 16931 33627 16943 33661
rect 16977 33627 16989 33661
rect 16931 33593 16989 33627
rect 16931 33559 16943 33593
rect 16977 33559 16989 33593
rect 16931 33525 16989 33559
rect 16931 33491 16943 33525
rect 16977 33491 16989 33525
rect 16931 33457 16989 33491
rect 16931 33423 16943 33457
rect 16977 33423 16989 33457
rect 16931 33389 16989 33423
rect 16931 33355 16943 33389
rect 16977 33355 16989 33389
rect 16931 33321 16989 33355
rect 16931 33287 16943 33321
rect 16977 33287 16989 33321
rect 16931 33253 16989 33287
rect 16931 33219 16943 33253
rect 16977 33219 16989 33253
rect 16931 33185 16989 33219
rect 16931 33151 16943 33185
rect 16977 33151 16989 33185
rect 16931 33117 16989 33151
rect 16931 33083 16943 33117
rect 16977 33083 16989 33117
rect 16931 33049 16989 33083
rect 16931 33015 16943 33049
rect 16977 33015 16989 33049
rect 16931 32981 16989 33015
rect 16931 32947 16943 32981
rect 16977 32947 16989 32981
rect 16931 32913 16989 32947
rect 16931 32879 16943 32913
rect 16977 32879 16989 32913
rect 16931 32845 16989 32879
rect 16931 32811 16943 32845
rect 16977 32811 16989 32845
rect 16931 32777 16989 32811
rect 16931 32743 16943 32777
rect 16977 32743 16989 32777
rect 16931 32709 16989 32743
rect 16931 32675 16943 32709
rect 16977 32675 16989 32709
rect 16931 32641 16989 32675
rect 16931 32607 16943 32641
rect 16977 32607 16989 32641
rect 16931 32573 16989 32607
rect 16931 32539 16943 32573
rect 16977 32539 16989 32573
rect 16931 32505 16989 32539
rect 16931 32471 16943 32505
rect 16977 32471 16989 32505
rect 16931 32437 16989 32471
rect 16931 32403 16943 32437
rect 16977 32403 16989 32437
rect 16931 32387 16989 32403
rect 17389 33661 17447 33677
rect 17389 33627 17401 33661
rect 17435 33627 17447 33661
rect 17389 33593 17447 33627
rect 17389 33559 17401 33593
rect 17435 33559 17447 33593
rect 17389 33525 17447 33559
rect 17389 33491 17401 33525
rect 17435 33491 17447 33525
rect 17389 33457 17447 33491
rect 17389 33423 17401 33457
rect 17435 33423 17447 33457
rect 17389 33389 17447 33423
rect 17389 33355 17401 33389
rect 17435 33355 17447 33389
rect 17389 33321 17447 33355
rect 17389 33287 17401 33321
rect 17435 33287 17447 33321
rect 17389 33253 17447 33287
rect 17389 33219 17401 33253
rect 17435 33219 17447 33253
rect 17389 33185 17447 33219
rect 17389 33151 17401 33185
rect 17435 33151 17447 33185
rect 17389 33117 17447 33151
rect 17389 33083 17401 33117
rect 17435 33083 17447 33117
rect 17389 33049 17447 33083
rect 17389 33015 17401 33049
rect 17435 33015 17447 33049
rect 17389 32981 17447 33015
rect 17389 32947 17401 32981
rect 17435 32947 17447 32981
rect 17389 32913 17447 32947
rect 17389 32879 17401 32913
rect 17435 32879 17447 32913
rect 17389 32845 17447 32879
rect 17389 32811 17401 32845
rect 17435 32811 17447 32845
rect 17389 32777 17447 32811
rect 17389 32743 17401 32777
rect 17435 32743 17447 32777
rect 17389 32709 17447 32743
rect 17389 32675 17401 32709
rect 17435 32675 17447 32709
rect 17389 32641 17447 32675
rect 17389 32607 17401 32641
rect 17435 32607 17447 32641
rect 17389 32573 17447 32607
rect 17389 32539 17401 32573
rect 17435 32539 17447 32573
rect 17389 32505 17447 32539
rect 17389 32471 17401 32505
rect 17435 32471 17447 32505
rect 17389 32437 17447 32471
rect 17389 32403 17401 32437
rect 17435 32403 17447 32437
rect 17389 32387 17447 32403
rect 17847 33661 17905 33677
rect 17847 33627 17859 33661
rect 17893 33627 17905 33661
rect 17847 33593 17905 33627
rect 17847 33559 17859 33593
rect 17893 33559 17905 33593
rect 17847 33525 17905 33559
rect 17847 33491 17859 33525
rect 17893 33491 17905 33525
rect 17847 33457 17905 33491
rect 17847 33423 17859 33457
rect 17893 33423 17905 33457
rect 17847 33389 17905 33423
rect 17847 33355 17859 33389
rect 17893 33355 17905 33389
rect 17847 33321 17905 33355
rect 17847 33287 17859 33321
rect 17893 33287 17905 33321
rect 17847 33253 17905 33287
rect 17847 33219 17859 33253
rect 17893 33219 17905 33253
rect 17847 33185 17905 33219
rect 17847 33151 17859 33185
rect 17893 33151 17905 33185
rect 17847 33117 17905 33151
rect 17847 33083 17859 33117
rect 17893 33083 17905 33117
rect 17847 33049 17905 33083
rect 17847 33015 17859 33049
rect 17893 33015 17905 33049
rect 17847 32981 17905 33015
rect 17847 32947 17859 32981
rect 17893 32947 17905 32981
rect 17847 32913 17905 32947
rect 17847 32879 17859 32913
rect 17893 32879 17905 32913
rect 17847 32845 17905 32879
rect 17847 32811 17859 32845
rect 17893 32811 17905 32845
rect 17847 32777 17905 32811
rect 17847 32743 17859 32777
rect 17893 32743 17905 32777
rect 17847 32709 17905 32743
rect 17847 32675 17859 32709
rect 17893 32675 17905 32709
rect 17847 32641 17905 32675
rect 17847 32607 17859 32641
rect 17893 32607 17905 32641
rect 17847 32573 17905 32607
rect 17847 32539 17859 32573
rect 17893 32539 17905 32573
rect 17847 32505 17905 32539
rect 17847 32471 17859 32505
rect 17893 32471 17905 32505
rect 17847 32437 17905 32471
rect 17847 32403 17859 32437
rect 17893 32403 17905 32437
rect 17847 32387 17905 32403
rect 18305 33661 18363 33677
rect 18305 33627 18317 33661
rect 18351 33627 18363 33661
rect 18305 33593 18363 33627
rect 18305 33559 18317 33593
rect 18351 33559 18363 33593
rect 18305 33525 18363 33559
rect 18305 33491 18317 33525
rect 18351 33491 18363 33525
rect 18305 33457 18363 33491
rect 18305 33423 18317 33457
rect 18351 33423 18363 33457
rect 18305 33389 18363 33423
rect 18305 33355 18317 33389
rect 18351 33355 18363 33389
rect 18305 33321 18363 33355
rect 18305 33287 18317 33321
rect 18351 33287 18363 33321
rect 18305 33253 18363 33287
rect 18305 33219 18317 33253
rect 18351 33219 18363 33253
rect 18305 33185 18363 33219
rect 18305 33151 18317 33185
rect 18351 33151 18363 33185
rect 18305 33117 18363 33151
rect 18305 33083 18317 33117
rect 18351 33083 18363 33117
rect 18305 33049 18363 33083
rect 18305 33015 18317 33049
rect 18351 33015 18363 33049
rect 18305 32981 18363 33015
rect 18305 32947 18317 32981
rect 18351 32947 18363 32981
rect 18305 32913 18363 32947
rect 18305 32879 18317 32913
rect 18351 32879 18363 32913
rect 18305 32845 18363 32879
rect 18305 32811 18317 32845
rect 18351 32811 18363 32845
rect 18305 32777 18363 32811
rect 18305 32743 18317 32777
rect 18351 32743 18363 32777
rect 18305 32709 18363 32743
rect 18305 32675 18317 32709
rect 18351 32675 18363 32709
rect 18305 32641 18363 32675
rect 18305 32607 18317 32641
rect 18351 32607 18363 32641
rect 18305 32573 18363 32607
rect 18305 32539 18317 32573
rect 18351 32539 18363 32573
rect 18305 32505 18363 32539
rect 18305 32471 18317 32505
rect 18351 32471 18363 32505
rect 18305 32437 18363 32471
rect 18305 32403 18317 32437
rect 18351 32403 18363 32437
rect 18305 32387 18363 32403
rect 18763 33661 18821 33677
rect 18763 33627 18775 33661
rect 18809 33627 18821 33661
rect 18763 33593 18821 33627
rect 18763 33559 18775 33593
rect 18809 33559 18821 33593
rect 18763 33525 18821 33559
rect 18763 33491 18775 33525
rect 18809 33491 18821 33525
rect 18763 33457 18821 33491
rect 18763 33423 18775 33457
rect 18809 33423 18821 33457
rect 18763 33389 18821 33423
rect 18763 33355 18775 33389
rect 18809 33355 18821 33389
rect 18763 33321 18821 33355
rect 18763 33287 18775 33321
rect 18809 33287 18821 33321
rect 18763 33253 18821 33287
rect 18763 33219 18775 33253
rect 18809 33219 18821 33253
rect 18763 33185 18821 33219
rect 18763 33151 18775 33185
rect 18809 33151 18821 33185
rect 18763 33117 18821 33151
rect 18763 33083 18775 33117
rect 18809 33083 18821 33117
rect 18763 33049 18821 33083
rect 18763 33015 18775 33049
rect 18809 33015 18821 33049
rect 18763 32981 18821 33015
rect 18763 32947 18775 32981
rect 18809 32947 18821 32981
rect 18763 32913 18821 32947
rect 18763 32879 18775 32913
rect 18809 32879 18821 32913
rect 18763 32845 18821 32879
rect 18763 32811 18775 32845
rect 18809 32811 18821 32845
rect 18763 32777 18821 32811
rect 18763 32743 18775 32777
rect 18809 32743 18821 32777
rect 18763 32709 18821 32743
rect 18763 32675 18775 32709
rect 18809 32675 18821 32709
rect 18763 32641 18821 32675
rect 18763 32607 18775 32641
rect 18809 32607 18821 32641
rect 18763 32573 18821 32607
rect 18763 32539 18775 32573
rect 18809 32539 18821 32573
rect 18763 32505 18821 32539
rect 18763 32471 18775 32505
rect 18809 32471 18821 32505
rect 18763 32437 18821 32471
rect 18763 32403 18775 32437
rect 18809 32403 18821 32437
rect 18763 32387 18821 32403
rect 19221 33661 19279 33677
rect 19221 33627 19233 33661
rect 19267 33627 19279 33661
rect 19221 33593 19279 33627
rect 19221 33559 19233 33593
rect 19267 33559 19279 33593
rect 19221 33525 19279 33559
rect 19221 33491 19233 33525
rect 19267 33491 19279 33525
rect 19221 33457 19279 33491
rect 19221 33423 19233 33457
rect 19267 33423 19279 33457
rect 19221 33389 19279 33423
rect 19221 33355 19233 33389
rect 19267 33355 19279 33389
rect 19221 33321 19279 33355
rect 19221 33287 19233 33321
rect 19267 33287 19279 33321
rect 19221 33253 19279 33287
rect 19221 33219 19233 33253
rect 19267 33219 19279 33253
rect 19221 33185 19279 33219
rect 19221 33151 19233 33185
rect 19267 33151 19279 33185
rect 19221 33117 19279 33151
rect 19221 33083 19233 33117
rect 19267 33083 19279 33117
rect 19221 33049 19279 33083
rect 19221 33015 19233 33049
rect 19267 33015 19279 33049
rect 19221 32981 19279 33015
rect 19221 32947 19233 32981
rect 19267 32947 19279 32981
rect 19221 32913 19279 32947
rect 19221 32879 19233 32913
rect 19267 32879 19279 32913
rect 19221 32845 19279 32879
rect 19221 32811 19233 32845
rect 19267 32811 19279 32845
rect 19221 32777 19279 32811
rect 19221 32743 19233 32777
rect 19267 32743 19279 32777
rect 19221 32709 19279 32743
rect 19221 32675 19233 32709
rect 19267 32675 19279 32709
rect 19221 32641 19279 32675
rect 19221 32607 19233 32641
rect 19267 32607 19279 32641
rect 19221 32573 19279 32607
rect 19221 32539 19233 32573
rect 19267 32539 19279 32573
rect 19221 32505 19279 32539
rect 19221 32471 19233 32505
rect 19267 32471 19279 32505
rect 19221 32437 19279 32471
rect 19221 32403 19233 32437
rect 19267 32403 19279 32437
rect 19221 32387 19279 32403
rect 19679 33661 19737 33677
rect 19679 33627 19691 33661
rect 19725 33627 19737 33661
rect 19679 33593 19737 33627
rect 19679 33559 19691 33593
rect 19725 33559 19737 33593
rect 19679 33525 19737 33559
rect 19679 33491 19691 33525
rect 19725 33491 19737 33525
rect 19679 33457 19737 33491
rect 19679 33423 19691 33457
rect 19725 33423 19737 33457
rect 19679 33389 19737 33423
rect 19679 33355 19691 33389
rect 19725 33355 19737 33389
rect 19679 33321 19737 33355
rect 19679 33287 19691 33321
rect 19725 33287 19737 33321
rect 19679 33253 19737 33287
rect 19679 33219 19691 33253
rect 19725 33219 19737 33253
rect 19679 33185 19737 33219
rect 19679 33151 19691 33185
rect 19725 33151 19737 33185
rect 19679 33117 19737 33151
rect 19679 33083 19691 33117
rect 19725 33083 19737 33117
rect 19679 33049 19737 33083
rect 19679 33015 19691 33049
rect 19725 33015 19737 33049
rect 19679 32981 19737 33015
rect 19679 32947 19691 32981
rect 19725 32947 19737 32981
rect 19679 32913 19737 32947
rect 19679 32879 19691 32913
rect 19725 32879 19737 32913
rect 19679 32845 19737 32879
rect 19679 32811 19691 32845
rect 19725 32811 19737 32845
rect 19679 32777 19737 32811
rect 19679 32743 19691 32777
rect 19725 32743 19737 32777
rect 19679 32709 19737 32743
rect 19679 32675 19691 32709
rect 19725 32675 19737 32709
rect 19679 32641 19737 32675
rect 19679 32607 19691 32641
rect 19725 32607 19737 32641
rect 19679 32573 19737 32607
rect 19679 32539 19691 32573
rect 19725 32539 19737 32573
rect 19679 32505 19737 32539
rect 19679 32471 19691 32505
rect 19725 32471 19737 32505
rect 19679 32437 19737 32471
rect 19679 32403 19691 32437
rect 19725 32403 19737 32437
rect 19679 32387 19737 32403
rect 20137 33661 20195 33677
rect 20137 33627 20149 33661
rect 20183 33627 20195 33661
rect 20137 33593 20195 33627
rect 20137 33559 20149 33593
rect 20183 33559 20195 33593
rect 20137 33525 20195 33559
rect 20137 33491 20149 33525
rect 20183 33491 20195 33525
rect 20137 33457 20195 33491
rect 20137 33423 20149 33457
rect 20183 33423 20195 33457
rect 20137 33389 20195 33423
rect 20137 33355 20149 33389
rect 20183 33355 20195 33389
rect 20137 33321 20195 33355
rect 20137 33287 20149 33321
rect 20183 33287 20195 33321
rect 20137 33253 20195 33287
rect 20137 33219 20149 33253
rect 20183 33219 20195 33253
rect 20137 33185 20195 33219
rect 20137 33151 20149 33185
rect 20183 33151 20195 33185
rect 20137 33117 20195 33151
rect 20137 33083 20149 33117
rect 20183 33083 20195 33117
rect 20137 33049 20195 33083
rect 20137 33015 20149 33049
rect 20183 33015 20195 33049
rect 20137 32981 20195 33015
rect 20137 32947 20149 32981
rect 20183 32947 20195 32981
rect 20137 32913 20195 32947
rect 20137 32879 20149 32913
rect 20183 32879 20195 32913
rect 20137 32845 20195 32879
rect 20137 32811 20149 32845
rect 20183 32811 20195 32845
rect 20137 32777 20195 32811
rect 20137 32743 20149 32777
rect 20183 32743 20195 32777
rect 20137 32709 20195 32743
rect 20137 32675 20149 32709
rect 20183 32675 20195 32709
rect 20137 32641 20195 32675
rect 20137 32607 20149 32641
rect 20183 32607 20195 32641
rect 20137 32573 20195 32607
rect 20137 32539 20149 32573
rect 20183 32539 20195 32573
rect 20137 32505 20195 32539
rect 20137 32471 20149 32505
rect 20183 32471 20195 32505
rect 20137 32437 20195 32471
rect 20137 32403 20149 32437
rect 20183 32403 20195 32437
rect 20137 32387 20195 32403
rect 20595 33661 20653 33677
rect 20595 33627 20607 33661
rect 20641 33627 20653 33661
rect 20595 33593 20653 33627
rect 20595 33559 20607 33593
rect 20641 33559 20653 33593
rect 20595 33525 20653 33559
rect 20595 33491 20607 33525
rect 20641 33491 20653 33525
rect 20595 33457 20653 33491
rect 20595 33423 20607 33457
rect 20641 33423 20653 33457
rect 20595 33389 20653 33423
rect 20595 33355 20607 33389
rect 20641 33355 20653 33389
rect 20595 33321 20653 33355
rect 20595 33287 20607 33321
rect 20641 33287 20653 33321
rect 20595 33253 20653 33287
rect 20595 33219 20607 33253
rect 20641 33219 20653 33253
rect 20595 33185 20653 33219
rect 20595 33151 20607 33185
rect 20641 33151 20653 33185
rect 20595 33117 20653 33151
rect 20595 33083 20607 33117
rect 20641 33083 20653 33117
rect 20595 33049 20653 33083
rect 20595 33015 20607 33049
rect 20641 33015 20653 33049
rect 20595 32981 20653 33015
rect 20595 32947 20607 32981
rect 20641 32947 20653 32981
rect 20595 32913 20653 32947
rect 20595 32879 20607 32913
rect 20641 32879 20653 32913
rect 20595 32845 20653 32879
rect 20595 32811 20607 32845
rect 20641 32811 20653 32845
rect 20595 32777 20653 32811
rect 20595 32743 20607 32777
rect 20641 32743 20653 32777
rect 20595 32709 20653 32743
rect 20595 32675 20607 32709
rect 20641 32675 20653 32709
rect 20595 32641 20653 32675
rect 20595 32607 20607 32641
rect 20641 32607 20653 32641
rect 20595 32573 20653 32607
rect 20595 32539 20607 32573
rect 20641 32539 20653 32573
rect 20595 32505 20653 32539
rect 20595 32471 20607 32505
rect 20641 32471 20653 32505
rect 20595 32437 20653 32471
rect 20595 32403 20607 32437
rect 20641 32403 20653 32437
rect 20595 32387 20653 32403
rect 21053 33661 21111 33677
rect 21053 33627 21065 33661
rect 21099 33627 21111 33661
rect 21053 33593 21111 33627
rect 21053 33559 21065 33593
rect 21099 33559 21111 33593
rect 21053 33525 21111 33559
rect 21053 33491 21065 33525
rect 21099 33491 21111 33525
rect 21053 33457 21111 33491
rect 21053 33423 21065 33457
rect 21099 33423 21111 33457
rect 21053 33389 21111 33423
rect 21053 33355 21065 33389
rect 21099 33355 21111 33389
rect 21053 33321 21111 33355
rect 21053 33287 21065 33321
rect 21099 33287 21111 33321
rect 21053 33253 21111 33287
rect 21053 33219 21065 33253
rect 21099 33219 21111 33253
rect 21053 33185 21111 33219
rect 21053 33151 21065 33185
rect 21099 33151 21111 33185
rect 21053 33117 21111 33151
rect 21053 33083 21065 33117
rect 21099 33083 21111 33117
rect 21053 33049 21111 33083
rect 21053 33015 21065 33049
rect 21099 33015 21111 33049
rect 21053 32981 21111 33015
rect 21053 32947 21065 32981
rect 21099 32947 21111 32981
rect 21053 32913 21111 32947
rect 21053 32879 21065 32913
rect 21099 32879 21111 32913
rect 21053 32845 21111 32879
rect 21053 32811 21065 32845
rect 21099 32811 21111 32845
rect 21053 32777 21111 32811
rect 21053 32743 21065 32777
rect 21099 32743 21111 32777
rect 21053 32709 21111 32743
rect 21053 32675 21065 32709
rect 21099 32675 21111 32709
rect 21053 32641 21111 32675
rect 21053 32607 21065 32641
rect 21099 32607 21111 32641
rect 21053 32573 21111 32607
rect 21053 32539 21065 32573
rect 21099 32539 21111 32573
rect 21053 32505 21111 32539
rect 21053 32471 21065 32505
rect 21099 32471 21111 32505
rect 21053 32437 21111 32471
rect 21053 32403 21065 32437
rect 21099 32403 21111 32437
rect 21053 32387 21111 32403
rect 21511 33661 21569 33677
rect 21511 33627 21523 33661
rect 21557 33627 21569 33661
rect 21511 33593 21569 33627
rect 21511 33559 21523 33593
rect 21557 33559 21569 33593
rect 21511 33525 21569 33559
rect 21511 33491 21523 33525
rect 21557 33491 21569 33525
rect 21511 33457 21569 33491
rect 21511 33423 21523 33457
rect 21557 33423 21569 33457
rect 21511 33389 21569 33423
rect 21511 33355 21523 33389
rect 21557 33355 21569 33389
rect 21511 33321 21569 33355
rect 21511 33287 21523 33321
rect 21557 33287 21569 33321
rect 21511 33253 21569 33287
rect 21511 33219 21523 33253
rect 21557 33219 21569 33253
rect 21511 33185 21569 33219
rect 21511 33151 21523 33185
rect 21557 33151 21569 33185
rect 21511 33117 21569 33151
rect 21511 33083 21523 33117
rect 21557 33083 21569 33117
rect 21511 33049 21569 33083
rect 21511 33015 21523 33049
rect 21557 33015 21569 33049
rect 21511 32981 21569 33015
rect 21511 32947 21523 32981
rect 21557 32947 21569 32981
rect 21511 32913 21569 32947
rect 21511 32879 21523 32913
rect 21557 32879 21569 32913
rect 21511 32845 21569 32879
rect 21511 32811 21523 32845
rect 21557 32811 21569 32845
rect 21511 32777 21569 32811
rect 21511 32743 21523 32777
rect 21557 32743 21569 32777
rect 21511 32709 21569 32743
rect 21511 32675 21523 32709
rect 21557 32675 21569 32709
rect 21511 32641 21569 32675
rect 21511 32607 21523 32641
rect 21557 32607 21569 32641
rect 21511 32573 21569 32607
rect 21511 32539 21523 32573
rect 21557 32539 21569 32573
rect 21511 32505 21569 32539
rect 21511 32471 21523 32505
rect 21557 32471 21569 32505
rect 21511 32437 21569 32471
rect 21511 32403 21523 32437
rect 21557 32403 21569 32437
rect 21511 32387 21569 32403
rect 21969 33661 22027 33677
rect 21969 33627 21981 33661
rect 22015 33627 22027 33661
rect 21969 33593 22027 33627
rect 21969 33559 21981 33593
rect 22015 33559 22027 33593
rect 21969 33525 22027 33559
rect 21969 33491 21981 33525
rect 22015 33491 22027 33525
rect 21969 33457 22027 33491
rect 21969 33423 21981 33457
rect 22015 33423 22027 33457
rect 21969 33389 22027 33423
rect 21969 33355 21981 33389
rect 22015 33355 22027 33389
rect 21969 33321 22027 33355
rect 21969 33287 21981 33321
rect 22015 33287 22027 33321
rect 21969 33253 22027 33287
rect 21969 33219 21981 33253
rect 22015 33219 22027 33253
rect 21969 33185 22027 33219
rect 21969 33151 21981 33185
rect 22015 33151 22027 33185
rect 21969 33117 22027 33151
rect 21969 33083 21981 33117
rect 22015 33083 22027 33117
rect 21969 33049 22027 33083
rect 21969 33015 21981 33049
rect 22015 33015 22027 33049
rect 21969 32981 22027 33015
rect 21969 32947 21981 32981
rect 22015 32947 22027 32981
rect 21969 32913 22027 32947
rect 21969 32879 21981 32913
rect 22015 32879 22027 32913
rect 21969 32845 22027 32879
rect 21969 32811 21981 32845
rect 22015 32811 22027 32845
rect 21969 32777 22027 32811
rect 21969 32743 21981 32777
rect 22015 32743 22027 32777
rect 21969 32709 22027 32743
rect 21969 32675 21981 32709
rect 22015 32675 22027 32709
rect 21969 32641 22027 32675
rect 21969 32607 21981 32641
rect 22015 32607 22027 32641
rect 21969 32573 22027 32607
rect 21969 32539 21981 32573
rect 22015 32539 22027 32573
rect 21969 32505 22027 32539
rect 21969 32471 21981 32505
rect 22015 32471 22027 32505
rect 21969 32437 22027 32471
rect 21969 32403 21981 32437
rect 22015 32403 22027 32437
rect 21969 32387 22027 32403
rect 22427 33661 22485 33677
rect 22427 33627 22439 33661
rect 22473 33627 22485 33661
rect 22427 33593 22485 33627
rect 22427 33559 22439 33593
rect 22473 33559 22485 33593
rect 22427 33525 22485 33559
rect 22427 33491 22439 33525
rect 22473 33491 22485 33525
rect 22427 33457 22485 33491
rect 22427 33423 22439 33457
rect 22473 33423 22485 33457
rect 22427 33389 22485 33423
rect 22427 33355 22439 33389
rect 22473 33355 22485 33389
rect 22427 33321 22485 33355
rect 22427 33287 22439 33321
rect 22473 33287 22485 33321
rect 22427 33253 22485 33287
rect 22427 33219 22439 33253
rect 22473 33219 22485 33253
rect 22427 33185 22485 33219
rect 22427 33151 22439 33185
rect 22473 33151 22485 33185
rect 22427 33117 22485 33151
rect 22427 33083 22439 33117
rect 22473 33083 22485 33117
rect 22427 33049 22485 33083
rect 22427 33015 22439 33049
rect 22473 33015 22485 33049
rect 22427 32981 22485 33015
rect 22427 32947 22439 32981
rect 22473 32947 22485 32981
rect 22427 32913 22485 32947
rect 22427 32879 22439 32913
rect 22473 32879 22485 32913
rect 22427 32845 22485 32879
rect 22427 32811 22439 32845
rect 22473 32811 22485 32845
rect 22427 32777 22485 32811
rect 22427 32743 22439 32777
rect 22473 32743 22485 32777
rect 22427 32709 22485 32743
rect 22427 32675 22439 32709
rect 22473 32675 22485 32709
rect 22427 32641 22485 32675
rect 22427 32607 22439 32641
rect 22473 32607 22485 32641
rect 22427 32573 22485 32607
rect 22427 32539 22439 32573
rect 22473 32539 22485 32573
rect 22427 32505 22485 32539
rect 22427 32471 22439 32505
rect 22473 32471 22485 32505
rect 22427 32437 22485 32471
rect 22427 32403 22439 32437
rect 22473 32403 22485 32437
rect 22427 32387 22485 32403
rect 22885 33661 22943 33677
rect 22885 33627 22897 33661
rect 22931 33627 22943 33661
rect 22885 33593 22943 33627
rect 22885 33559 22897 33593
rect 22931 33559 22943 33593
rect 22885 33525 22943 33559
rect 22885 33491 22897 33525
rect 22931 33491 22943 33525
rect 22885 33457 22943 33491
rect 22885 33423 22897 33457
rect 22931 33423 22943 33457
rect 22885 33389 22943 33423
rect 22885 33355 22897 33389
rect 22931 33355 22943 33389
rect 22885 33321 22943 33355
rect 22885 33287 22897 33321
rect 22931 33287 22943 33321
rect 22885 33253 22943 33287
rect 22885 33219 22897 33253
rect 22931 33219 22943 33253
rect 22885 33185 22943 33219
rect 22885 33151 22897 33185
rect 22931 33151 22943 33185
rect 22885 33117 22943 33151
rect 22885 33083 22897 33117
rect 22931 33083 22943 33117
rect 22885 33049 22943 33083
rect 22885 33015 22897 33049
rect 22931 33015 22943 33049
rect 22885 32981 22943 33015
rect 22885 32947 22897 32981
rect 22931 32947 22943 32981
rect 22885 32913 22943 32947
rect 22885 32879 22897 32913
rect 22931 32879 22943 32913
rect 22885 32845 22943 32879
rect 22885 32811 22897 32845
rect 22931 32811 22943 32845
rect 22885 32777 22943 32811
rect 22885 32743 22897 32777
rect 22931 32743 22943 32777
rect 22885 32709 22943 32743
rect 22885 32675 22897 32709
rect 22931 32675 22943 32709
rect 22885 32641 22943 32675
rect 22885 32607 22897 32641
rect 22931 32607 22943 32641
rect 22885 32573 22943 32607
rect 22885 32539 22897 32573
rect 22931 32539 22943 32573
rect 22885 32505 22943 32539
rect 22885 32471 22897 32505
rect 22931 32471 22943 32505
rect 22885 32437 22943 32471
rect 22885 32403 22897 32437
rect 22931 32403 22943 32437
rect 22885 32387 22943 32403
rect 23343 33661 23401 33677
rect 23343 33627 23355 33661
rect 23389 33627 23401 33661
rect 23343 33593 23401 33627
rect 23343 33559 23355 33593
rect 23389 33559 23401 33593
rect 23343 33525 23401 33559
rect 23343 33491 23355 33525
rect 23389 33491 23401 33525
rect 23343 33457 23401 33491
rect 23343 33423 23355 33457
rect 23389 33423 23401 33457
rect 23343 33389 23401 33423
rect 23343 33355 23355 33389
rect 23389 33355 23401 33389
rect 23343 33321 23401 33355
rect 23343 33287 23355 33321
rect 23389 33287 23401 33321
rect 23343 33253 23401 33287
rect 23343 33219 23355 33253
rect 23389 33219 23401 33253
rect 23343 33185 23401 33219
rect 23343 33151 23355 33185
rect 23389 33151 23401 33185
rect 23343 33117 23401 33151
rect 23343 33083 23355 33117
rect 23389 33083 23401 33117
rect 23343 33049 23401 33083
rect 23343 33015 23355 33049
rect 23389 33015 23401 33049
rect 23343 32981 23401 33015
rect 23343 32947 23355 32981
rect 23389 32947 23401 32981
rect 23343 32913 23401 32947
rect 23343 32879 23355 32913
rect 23389 32879 23401 32913
rect 23343 32845 23401 32879
rect 23343 32811 23355 32845
rect 23389 32811 23401 32845
rect 23343 32777 23401 32811
rect 23343 32743 23355 32777
rect 23389 32743 23401 32777
rect 23343 32709 23401 32743
rect 23343 32675 23355 32709
rect 23389 32675 23401 32709
rect 23343 32641 23401 32675
rect 23343 32607 23355 32641
rect 23389 32607 23401 32641
rect 23343 32573 23401 32607
rect 23343 32539 23355 32573
rect 23389 32539 23401 32573
rect 23343 32505 23401 32539
rect 23343 32471 23355 32505
rect 23389 32471 23401 32505
rect 23343 32437 23401 32471
rect 23343 32403 23355 32437
rect 23389 32403 23401 32437
rect 23343 32387 23401 32403
rect 23801 33661 23859 33677
rect 23801 33627 23813 33661
rect 23847 33627 23859 33661
rect 23801 33593 23859 33627
rect 23801 33559 23813 33593
rect 23847 33559 23859 33593
rect 23801 33525 23859 33559
rect 23801 33491 23813 33525
rect 23847 33491 23859 33525
rect 23801 33457 23859 33491
rect 23801 33423 23813 33457
rect 23847 33423 23859 33457
rect 23801 33389 23859 33423
rect 23801 33355 23813 33389
rect 23847 33355 23859 33389
rect 23801 33321 23859 33355
rect 23801 33287 23813 33321
rect 23847 33287 23859 33321
rect 23801 33253 23859 33287
rect 23801 33219 23813 33253
rect 23847 33219 23859 33253
rect 23801 33185 23859 33219
rect 23801 33151 23813 33185
rect 23847 33151 23859 33185
rect 23801 33117 23859 33151
rect 23801 33083 23813 33117
rect 23847 33083 23859 33117
rect 23801 33049 23859 33083
rect 23801 33015 23813 33049
rect 23847 33015 23859 33049
rect 23801 32981 23859 33015
rect 23801 32947 23813 32981
rect 23847 32947 23859 32981
rect 23801 32913 23859 32947
rect 23801 32879 23813 32913
rect 23847 32879 23859 32913
rect 23801 32845 23859 32879
rect 23801 32811 23813 32845
rect 23847 32811 23859 32845
rect 23801 32777 23859 32811
rect 23801 32743 23813 32777
rect 23847 32743 23859 32777
rect 23801 32709 23859 32743
rect 23801 32675 23813 32709
rect 23847 32675 23859 32709
rect 23801 32641 23859 32675
rect 23801 32607 23813 32641
rect 23847 32607 23859 32641
rect 23801 32573 23859 32607
rect 23801 32539 23813 32573
rect 23847 32539 23859 32573
rect 23801 32505 23859 32539
rect 23801 32471 23813 32505
rect 23847 32471 23859 32505
rect 23801 32437 23859 32471
rect 23801 32403 23813 32437
rect 23847 32403 23859 32437
rect 23801 32387 23859 32403
rect 24259 33661 24317 33677
rect 24259 33627 24271 33661
rect 24305 33627 24317 33661
rect 24259 33593 24317 33627
rect 24259 33559 24271 33593
rect 24305 33559 24317 33593
rect 24259 33525 24317 33559
rect 24259 33491 24271 33525
rect 24305 33491 24317 33525
rect 24259 33457 24317 33491
rect 24259 33423 24271 33457
rect 24305 33423 24317 33457
rect 24259 33389 24317 33423
rect 24259 33355 24271 33389
rect 24305 33355 24317 33389
rect 24259 33321 24317 33355
rect 24259 33287 24271 33321
rect 24305 33287 24317 33321
rect 24259 33253 24317 33287
rect 24259 33219 24271 33253
rect 24305 33219 24317 33253
rect 24259 33185 24317 33219
rect 24259 33151 24271 33185
rect 24305 33151 24317 33185
rect 24259 33117 24317 33151
rect 24259 33083 24271 33117
rect 24305 33083 24317 33117
rect 24259 33049 24317 33083
rect 24259 33015 24271 33049
rect 24305 33015 24317 33049
rect 24259 32981 24317 33015
rect 24259 32947 24271 32981
rect 24305 32947 24317 32981
rect 24259 32913 24317 32947
rect 24259 32879 24271 32913
rect 24305 32879 24317 32913
rect 24259 32845 24317 32879
rect 24259 32811 24271 32845
rect 24305 32811 24317 32845
rect 24259 32777 24317 32811
rect 24259 32743 24271 32777
rect 24305 32743 24317 32777
rect 24259 32709 24317 32743
rect 24259 32675 24271 32709
rect 24305 32675 24317 32709
rect 24259 32641 24317 32675
rect 24259 32607 24271 32641
rect 24305 32607 24317 32641
rect 24259 32573 24317 32607
rect 24259 32539 24271 32573
rect 24305 32539 24317 32573
rect 24259 32505 24317 32539
rect 24259 32471 24271 32505
rect 24305 32471 24317 32505
rect 24259 32437 24317 32471
rect 24259 32403 24271 32437
rect 24305 32403 24317 32437
rect 24259 32387 24317 32403
rect 24717 33661 24775 33677
rect 24717 33627 24729 33661
rect 24763 33627 24775 33661
rect 24717 33593 24775 33627
rect 24717 33559 24729 33593
rect 24763 33559 24775 33593
rect 24717 33525 24775 33559
rect 24717 33491 24729 33525
rect 24763 33491 24775 33525
rect 24717 33457 24775 33491
rect 24717 33423 24729 33457
rect 24763 33423 24775 33457
rect 24717 33389 24775 33423
rect 24717 33355 24729 33389
rect 24763 33355 24775 33389
rect 24717 33321 24775 33355
rect 24717 33287 24729 33321
rect 24763 33287 24775 33321
rect 24717 33253 24775 33287
rect 24717 33219 24729 33253
rect 24763 33219 24775 33253
rect 24717 33185 24775 33219
rect 24717 33151 24729 33185
rect 24763 33151 24775 33185
rect 24717 33117 24775 33151
rect 24717 33083 24729 33117
rect 24763 33083 24775 33117
rect 24717 33049 24775 33083
rect 24717 33015 24729 33049
rect 24763 33015 24775 33049
rect 24717 32981 24775 33015
rect 24717 32947 24729 32981
rect 24763 32947 24775 32981
rect 24717 32913 24775 32947
rect 24717 32879 24729 32913
rect 24763 32879 24775 32913
rect 24717 32845 24775 32879
rect 24717 32811 24729 32845
rect 24763 32811 24775 32845
rect 24717 32777 24775 32811
rect 24717 32743 24729 32777
rect 24763 32743 24775 32777
rect 24717 32709 24775 32743
rect 24717 32675 24729 32709
rect 24763 32675 24775 32709
rect 24717 32641 24775 32675
rect 24717 32607 24729 32641
rect 24763 32607 24775 32641
rect 24717 32573 24775 32607
rect 24717 32539 24729 32573
rect 24763 32539 24775 32573
rect 24717 32505 24775 32539
rect 24717 32471 24729 32505
rect 24763 32471 24775 32505
rect 24717 32437 24775 32471
rect 24717 32403 24729 32437
rect 24763 32403 24775 32437
rect 24717 32387 24775 32403
rect 25175 33661 25233 33677
rect 25175 33627 25187 33661
rect 25221 33627 25233 33661
rect 25175 33593 25233 33627
rect 25175 33559 25187 33593
rect 25221 33559 25233 33593
rect 25175 33525 25233 33559
rect 25175 33491 25187 33525
rect 25221 33491 25233 33525
rect 25175 33457 25233 33491
rect 25175 33423 25187 33457
rect 25221 33423 25233 33457
rect 25175 33389 25233 33423
rect 25175 33355 25187 33389
rect 25221 33355 25233 33389
rect 25175 33321 25233 33355
rect 25175 33287 25187 33321
rect 25221 33287 25233 33321
rect 25175 33253 25233 33287
rect 25175 33219 25187 33253
rect 25221 33219 25233 33253
rect 25175 33185 25233 33219
rect 25175 33151 25187 33185
rect 25221 33151 25233 33185
rect 25175 33117 25233 33151
rect 25175 33083 25187 33117
rect 25221 33083 25233 33117
rect 25175 33049 25233 33083
rect 25175 33015 25187 33049
rect 25221 33015 25233 33049
rect 25175 32981 25233 33015
rect 25175 32947 25187 32981
rect 25221 32947 25233 32981
rect 25175 32913 25233 32947
rect 25175 32879 25187 32913
rect 25221 32879 25233 32913
rect 25175 32845 25233 32879
rect 25175 32811 25187 32845
rect 25221 32811 25233 32845
rect 25175 32777 25233 32811
rect 25175 32743 25187 32777
rect 25221 32743 25233 32777
rect 25175 32709 25233 32743
rect 25175 32675 25187 32709
rect 25221 32675 25233 32709
rect 25175 32641 25233 32675
rect 25175 32607 25187 32641
rect 25221 32607 25233 32641
rect 25175 32573 25233 32607
rect 25175 32539 25187 32573
rect 25221 32539 25233 32573
rect 25175 32505 25233 32539
rect 25175 32471 25187 32505
rect 25221 32471 25233 32505
rect 25175 32437 25233 32471
rect 25175 32403 25187 32437
rect 25221 32403 25233 32437
rect 25175 32387 25233 32403
rect 25633 33661 25691 33677
rect 25633 33627 25645 33661
rect 25679 33627 25691 33661
rect 25633 33593 25691 33627
rect 25633 33559 25645 33593
rect 25679 33559 25691 33593
rect 25633 33525 25691 33559
rect 25633 33491 25645 33525
rect 25679 33491 25691 33525
rect 25633 33457 25691 33491
rect 25633 33423 25645 33457
rect 25679 33423 25691 33457
rect 25633 33389 25691 33423
rect 25633 33355 25645 33389
rect 25679 33355 25691 33389
rect 25633 33321 25691 33355
rect 25633 33287 25645 33321
rect 25679 33287 25691 33321
rect 25633 33253 25691 33287
rect 25633 33219 25645 33253
rect 25679 33219 25691 33253
rect 25633 33185 25691 33219
rect 25633 33151 25645 33185
rect 25679 33151 25691 33185
rect 25633 33117 25691 33151
rect 25633 33083 25645 33117
rect 25679 33083 25691 33117
rect 25633 33049 25691 33083
rect 25633 33015 25645 33049
rect 25679 33015 25691 33049
rect 25633 32981 25691 33015
rect 25633 32947 25645 32981
rect 25679 32947 25691 32981
rect 25633 32913 25691 32947
rect 25633 32879 25645 32913
rect 25679 32879 25691 32913
rect 25633 32845 25691 32879
rect 25633 32811 25645 32845
rect 25679 32811 25691 32845
rect 25633 32777 25691 32811
rect 25633 32743 25645 32777
rect 25679 32743 25691 32777
rect 25633 32709 25691 32743
rect 25633 32675 25645 32709
rect 25679 32675 25691 32709
rect 25633 32641 25691 32675
rect 25633 32607 25645 32641
rect 25679 32607 25691 32641
rect 25633 32573 25691 32607
rect 25633 32539 25645 32573
rect 25679 32539 25691 32573
rect 25633 32505 25691 32539
rect 25633 32471 25645 32505
rect 25679 32471 25691 32505
rect 25633 32437 25691 32471
rect 25633 32403 25645 32437
rect 25679 32403 25691 32437
rect 25633 32387 25691 32403
rect 26091 33661 26149 33677
rect 26091 33627 26103 33661
rect 26137 33627 26149 33661
rect 26091 33593 26149 33627
rect 26091 33559 26103 33593
rect 26137 33559 26149 33593
rect 26091 33525 26149 33559
rect 26091 33491 26103 33525
rect 26137 33491 26149 33525
rect 26091 33457 26149 33491
rect 26091 33423 26103 33457
rect 26137 33423 26149 33457
rect 26091 33389 26149 33423
rect 26091 33355 26103 33389
rect 26137 33355 26149 33389
rect 26091 33321 26149 33355
rect 26091 33287 26103 33321
rect 26137 33287 26149 33321
rect 26091 33253 26149 33287
rect 26091 33219 26103 33253
rect 26137 33219 26149 33253
rect 26091 33185 26149 33219
rect 26091 33151 26103 33185
rect 26137 33151 26149 33185
rect 26091 33117 26149 33151
rect 26091 33083 26103 33117
rect 26137 33083 26149 33117
rect 26091 33049 26149 33083
rect 26091 33015 26103 33049
rect 26137 33015 26149 33049
rect 26091 32981 26149 33015
rect 26091 32947 26103 32981
rect 26137 32947 26149 32981
rect 26091 32913 26149 32947
rect 26091 32879 26103 32913
rect 26137 32879 26149 32913
rect 26091 32845 26149 32879
rect 26091 32811 26103 32845
rect 26137 32811 26149 32845
rect 26091 32777 26149 32811
rect 26091 32743 26103 32777
rect 26137 32743 26149 32777
rect 26091 32709 26149 32743
rect 26091 32675 26103 32709
rect 26137 32675 26149 32709
rect 26091 32641 26149 32675
rect 26091 32607 26103 32641
rect 26137 32607 26149 32641
rect 26091 32573 26149 32607
rect 26091 32539 26103 32573
rect 26137 32539 26149 32573
rect 26091 32505 26149 32539
rect 26091 32471 26103 32505
rect 26137 32471 26149 32505
rect 26091 32437 26149 32471
rect 26091 32403 26103 32437
rect 26137 32403 26149 32437
rect 26091 32387 26149 32403
rect 26549 33661 26607 33677
rect 26549 33627 26561 33661
rect 26595 33627 26607 33661
rect 26549 33593 26607 33627
rect 26549 33559 26561 33593
rect 26595 33559 26607 33593
rect 26549 33525 26607 33559
rect 26549 33491 26561 33525
rect 26595 33491 26607 33525
rect 26549 33457 26607 33491
rect 26549 33423 26561 33457
rect 26595 33423 26607 33457
rect 26549 33389 26607 33423
rect 26549 33355 26561 33389
rect 26595 33355 26607 33389
rect 26549 33321 26607 33355
rect 26549 33287 26561 33321
rect 26595 33287 26607 33321
rect 26549 33253 26607 33287
rect 26549 33219 26561 33253
rect 26595 33219 26607 33253
rect 26549 33185 26607 33219
rect 26549 33151 26561 33185
rect 26595 33151 26607 33185
rect 26549 33117 26607 33151
rect 26549 33083 26561 33117
rect 26595 33083 26607 33117
rect 26549 33049 26607 33083
rect 26549 33015 26561 33049
rect 26595 33015 26607 33049
rect 26549 32981 26607 33015
rect 26549 32947 26561 32981
rect 26595 32947 26607 32981
rect 26549 32913 26607 32947
rect 26549 32879 26561 32913
rect 26595 32879 26607 32913
rect 26549 32845 26607 32879
rect 26549 32811 26561 32845
rect 26595 32811 26607 32845
rect 26549 32777 26607 32811
rect 26549 32743 26561 32777
rect 26595 32743 26607 32777
rect 26549 32709 26607 32743
rect 26549 32675 26561 32709
rect 26595 32675 26607 32709
rect 26549 32641 26607 32675
rect 26549 32607 26561 32641
rect 26595 32607 26607 32641
rect 26549 32573 26607 32607
rect 26549 32539 26561 32573
rect 26595 32539 26607 32573
rect 26549 32505 26607 32539
rect 26549 32471 26561 32505
rect 26595 32471 26607 32505
rect 26549 32437 26607 32471
rect 26549 32403 26561 32437
rect 26595 32403 26607 32437
rect 26549 32387 26607 32403
rect 27007 33661 27065 33677
rect 27007 33627 27019 33661
rect 27053 33627 27065 33661
rect 27007 33593 27065 33627
rect 27007 33559 27019 33593
rect 27053 33559 27065 33593
rect 27007 33525 27065 33559
rect 27007 33491 27019 33525
rect 27053 33491 27065 33525
rect 27007 33457 27065 33491
rect 27007 33423 27019 33457
rect 27053 33423 27065 33457
rect 27007 33389 27065 33423
rect 27007 33355 27019 33389
rect 27053 33355 27065 33389
rect 27007 33321 27065 33355
rect 27007 33287 27019 33321
rect 27053 33287 27065 33321
rect 27007 33253 27065 33287
rect 27007 33219 27019 33253
rect 27053 33219 27065 33253
rect 27007 33185 27065 33219
rect 27007 33151 27019 33185
rect 27053 33151 27065 33185
rect 27007 33117 27065 33151
rect 27007 33083 27019 33117
rect 27053 33083 27065 33117
rect 27007 33049 27065 33083
rect 27007 33015 27019 33049
rect 27053 33015 27065 33049
rect 27007 32981 27065 33015
rect 27007 32947 27019 32981
rect 27053 32947 27065 32981
rect 27007 32913 27065 32947
rect 27007 32879 27019 32913
rect 27053 32879 27065 32913
rect 27007 32845 27065 32879
rect 27007 32811 27019 32845
rect 27053 32811 27065 32845
rect 27007 32777 27065 32811
rect 27007 32743 27019 32777
rect 27053 32743 27065 32777
rect 27007 32709 27065 32743
rect 27007 32675 27019 32709
rect 27053 32675 27065 32709
rect 27007 32641 27065 32675
rect 27007 32607 27019 32641
rect 27053 32607 27065 32641
rect 27007 32573 27065 32607
rect 27007 32539 27019 32573
rect 27053 32539 27065 32573
rect 27007 32505 27065 32539
rect 27007 32471 27019 32505
rect 27053 32471 27065 32505
rect 27007 32437 27065 32471
rect 27007 32403 27019 32437
rect 27053 32403 27065 32437
rect 27007 32387 27065 32403
rect 27465 33661 27523 33677
rect 27465 33627 27477 33661
rect 27511 33627 27523 33661
rect 27465 33593 27523 33627
rect 27465 33559 27477 33593
rect 27511 33559 27523 33593
rect 27465 33525 27523 33559
rect 27465 33491 27477 33525
rect 27511 33491 27523 33525
rect 27465 33457 27523 33491
rect 27465 33423 27477 33457
rect 27511 33423 27523 33457
rect 27465 33389 27523 33423
rect 27465 33355 27477 33389
rect 27511 33355 27523 33389
rect 27465 33321 27523 33355
rect 27465 33287 27477 33321
rect 27511 33287 27523 33321
rect 27465 33253 27523 33287
rect 27465 33219 27477 33253
rect 27511 33219 27523 33253
rect 27465 33185 27523 33219
rect 27465 33151 27477 33185
rect 27511 33151 27523 33185
rect 27465 33117 27523 33151
rect 27465 33083 27477 33117
rect 27511 33083 27523 33117
rect 27465 33049 27523 33083
rect 27465 33015 27477 33049
rect 27511 33015 27523 33049
rect 27465 32981 27523 33015
rect 27465 32947 27477 32981
rect 27511 32947 27523 32981
rect 27465 32913 27523 32947
rect 27465 32879 27477 32913
rect 27511 32879 27523 32913
rect 27465 32845 27523 32879
rect 27465 32811 27477 32845
rect 27511 32811 27523 32845
rect 27465 32777 27523 32811
rect 27465 32743 27477 32777
rect 27511 32743 27523 32777
rect 27465 32709 27523 32743
rect 27465 32675 27477 32709
rect 27511 32675 27523 32709
rect 27465 32641 27523 32675
rect 27465 32607 27477 32641
rect 27511 32607 27523 32641
rect 27465 32573 27523 32607
rect 27465 32539 27477 32573
rect 27511 32539 27523 32573
rect 27465 32505 27523 32539
rect 27465 32471 27477 32505
rect 27511 32471 27523 32505
rect 27465 32437 27523 32471
rect 27465 32403 27477 32437
rect 27511 32403 27523 32437
rect 27465 32387 27523 32403
rect 27923 33661 27981 33677
rect 27923 33627 27935 33661
rect 27969 33627 27981 33661
rect 27923 33593 27981 33627
rect 27923 33559 27935 33593
rect 27969 33559 27981 33593
rect 27923 33525 27981 33559
rect 27923 33491 27935 33525
rect 27969 33491 27981 33525
rect 27923 33457 27981 33491
rect 27923 33423 27935 33457
rect 27969 33423 27981 33457
rect 27923 33389 27981 33423
rect 27923 33355 27935 33389
rect 27969 33355 27981 33389
rect 27923 33321 27981 33355
rect 27923 33287 27935 33321
rect 27969 33287 27981 33321
rect 27923 33253 27981 33287
rect 27923 33219 27935 33253
rect 27969 33219 27981 33253
rect 27923 33185 27981 33219
rect 27923 33151 27935 33185
rect 27969 33151 27981 33185
rect 27923 33117 27981 33151
rect 27923 33083 27935 33117
rect 27969 33083 27981 33117
rect 27923 33049 27981 33083
rect 27923 33015 27935 33049
rect 27969 33015 27981 33049
rect 27923 32981 27981 33015
rect 27923 32947 27935 32981
rect 27969 32947 27981 32981
rect 27923 32913 27981 32947
rect 27923 32879 27935 32913
rect 27969 32879 27981 32913
rect 27923 32845 27981 32879
rect 27923 32811 27935 32845
rect 27969 32811 27981 32845
rect 27923 32777 27981 32811
rect 27923 32743 27935 32777
rect 27969 32743 27981 32777
rect 27923 32709 27981 32743
rect 27923 32675 27935 32709
rect 27969 32675 27981 32709
rect 27923 32641 27981 32675
rect 27923 32607 27935 32641
rect 27969 32607 27981 32641
rect 27923 32573 27981 32607
rect 27923 32539 27935 32573
rect 27969 32539 27981 32573
rect 27923 32505 27981 32539
rect 27923 32471 27935 32505
rect 27969 32471 27981 32505
rect 27923 32437 27981 32471
rect 27923 32403 27935 32437
rect 27969 32403 27981 32437
rect 27923 32387 27981 32403
rect 28381 33661 28439 33677
rect 28381 33627 28393 33661
rect 28427 33627 28439 33661
rect 28381 33593 28439 33627
rect 28381 33559 28393 33593
rect 28427 33559 28439 33593
rect 28381 33525 28439 33559
rect 28381 33491 28393 33525
rect 28427 33491 28439 33525
rect 28381 33457 28439 33491
rect 28381 33423 28393 33457
rect 28427 33423 28439 33457
rect 28381 33389 28439 33423
rect 28381 33355 28393 33389
rect 28427 33355 28439 33389
rect 28381 33321 28439 33355
rect 28381 33287 28393 33321
rect 28427 33287 28439 33321
rect 28381 33253 28439 33287
rect 28381 33219 28393 33253
rect 28427 33219 28439 33253
rect 28381 33185 28439 33219
rect 28381 33151 28393 33185
rect 28427 33151 28439 33185
rect 28381 33117 28439 33151
rect 28381 33083 28393 33117
rect 28427 33083 28439 33117
rect 28381 33049 28439 33083
rect 28381 33015 28393 33049
rect 28427 33015 28439 33049
rect 28381 32981 28439 33015
rect 28381 32947 28393 32981
rect 28427 32947 28439 32981
rect 28381 32913 28439 32947
rect 28381 32879 28393 32913
rect 28427 32879 28439 32913
rect 28381 32845 28439 32879
rect 28381 32811 28393 32845
rect 28427 32811 28439 32845
rect 28381 32777 28439 32811
rect 28381 32743 28393 32777
rect 28427 32743 28439 32777
rect 28381 32709 28439 32743
rect 28381 32675 28393 32709
rect 28427 32675 28439 32709
rect 28381 32641 28439 32675
rect 28381 32607 28393 32641
rect 28427 32607 28439 32641
rect 28381 32573 28439 32607
rect 28381 32539 28393 32573
rect 28427 32539 28439 32573
rect 28381 32505 28439 32539
rect 28381 32471 28393 32505
rect 28427 32471 28439 32505
rect 28381 32437 28439 32471
rect 28381 32403 28393 32437
rect 28427 32403 28439 32437
rect 28381 32387 28439 32403
rect 28839 33661 28897 33677
rect 28839 33627 28851 33661
rect 28885 33627 28897 33661
rect 28839 33593 28897 33627
rect 28839 33559 28851 33593
rect 28885 33559 28897 33593
rect 28839 33525 28897 33559
rect 28839 33491 28851 33525
rect 28885 33491 28897 33525
rect 28839 33457 28897 33491
rect 28839 33423 28851 33457
rect 28885 33423 28897 33457
rect 28839 33389 28897 33423
rect 28839 33355 28851 33389
rect 28885 33355 28897 33389
rect 28839 33321 28897 33355
rect 28839 33287 28851 33321
rect 28885 33287 28897 33321
rect 28839 33253 28897 33287
rect 28839 33219 28851 33253
rect 28885 33219 28897 33253
rect 28839 33185 28897 33219
rect 28839 33151 28851 33185
rect 28885 33151 28897 33185
rect 28839 33117 28897 33151
rect 28839 33083 28851 33117
rect 28885 33083 28897 33117
rect 28839 33049 28897 33083
rect 28839 33015 28851 33049
rect 28885 33015 28897 33049
rect 28839 32981 28897 33015
rect 28839 32947 28851 32981
rect 28885 32947 28897 32981
rect 28839 32913 28897 32947
rect 28839 32879 28851 32913
rect 28885 32879 28897 32913
rect 28839 32845 28897 32879
rect 28839 32811 28851 32845
rect 28885 32811 28897 32845
rect 28839 32777 28897 32811
rect 28839 32743 28851 32777
rect 28885 32743 28897 32777
rect 28839 32709 28897 32743
rect 28839 32675 28851 32709
rect 28885 32675 28897 32709
rect 28839 32641 28897 32675
rect 28839 32607 28851 32641
rect 28885 32607 28897 32641
rect 28839 32573 28897 32607
rect 28839 32539 28851 32573
rect 28885 32539 28897 32573
rect 28839 32505 28897 32539
rect 28839 32471 28851 32505
rect 28885 32471 28897 32505
rect 28839 32437 28897 32471
rect 28839 32403 28851 32437
rect 28885 32403 28897 32437
rect 28839 32387 28897 32403
rect 29297 33661 29355 33677
rect 29297 33627 29309 33661
rect 29343 33627 29355 33661
rect 29297 33593 29355 33627
rect 29297 33559 29309 33593
rect 29343 33559 29355 33593
rect 29297 33525 29355 33559
rect 29297 33491 29309 33525
rect 29343 33491 29355 33525
rect 29297 33457 29355 33491
rect 29297 33423 29309 33457
rect 29343 33423 29355 33457
rect 29297 33389 29355 33423
rect 29297 33355 29309 33389
rect 29343 33355 29355 33389
rect 29297 33321 29355 33355
rect 29297 33287 29309 33321
rect 29343 33287 29355 33321
rect 29297 33253 29355 33287
rect 29297 33219 29309 33253
rect 29343 33219 29355 33253
rect 29297 33185 29355 33219
rect 29297 33151 29309 33185
rect 29343 33151 29355 33185
rect 29297 33117 29355 33151
rect 29297 33083 29309 33117
rect 29343 33083 29355 33117
rect 29297 33049 29355 33083
rect 29297 33015 29309 33049
rect 29343 33015 29355 33049
rect 29297 32981 29355 33015
rect 29297 32947 29309 32981
rect 29343 32947 29355 32981
rect 29297 32913 29355 32947
rect 29297 32879 29309 32913
rect 29343 32879 29355 32913
rect 29297 32845 29355 32879
rect 29297 32811 29309 32845
rect 29343 32811 29355 32845
rect 29297 32777 29355 32811
rect 29297 32743 29309 32777
rect 29343 32743 29355 32777
rect 29297 32709 29355 32743
rect 29297 32675 29309 32709
rect 29343 32675 29355 32709
rect 29297 32641 29355 32675
rect 29297 32607 29309 32641
rect 29343 32607 29355 32641
rect 29297 32573 29355 32607
rect 29297 32539 29309 32573
rect 29343 32539 29355 32573
rect 29297 32505 29355 32539
rect 29297 32471 29309 32505
rect 29343 32471 29355 32505
rect 29297 32437 29355 32471
rect 29297 32403 29309 32437
rect 29343 32403 29355 32437
rect 29297 32387 29355 32403
rect 29755 33661 29813 33677
rect 29755 33627 29767 33661
rect 29801 33627 29813 33661
rect 29755 33593 29813 33627
rect 29755 33559 29767 33593
rect 29801 33559 29813 33593
rect 29755 33525 29813 33559
rect 29755 33491 29767 33525
rect 29801 33491 29813 33525
rect 29755 33457 29813 33491
rect 29755 33423 29767 33457
rect 29801 33423 29813 33457
rect 29755 33389 29813 33423
rect 29755 33355 29767 33389
rect 29801 33355 29813 33389
rect 29755 33321 29813 33355
rect 29755 33287 29767 33321
rect 29801 33287 29813 33321
rect 29755 33253 29813 33287
rect 29755 33219 29767 33253
rect 29801 33219 29813 33253
rect 29755 33185 29813 33219
rect 29755 33151 29767 33185
rect 29801 33151 29813 33185
rect 29755 33117 29813 33151
rect 29755 33083 29767 33117
rect 29801 33083 29813 33117
rect 29755 33049 29813 33083
rect 29755 33015 29767 33049
rect 29801 33015 29813 33049
rect 29755 32981 29813 33015
rect 29755 32947 29767 32981
rect 29801 32947 29813 32981
rect 29755 32913 29813 32947
rect 29755 32879 29767 32913
rect 29801 32879 29813 32913
rect 29755 32845 29813 32879
rect 29755 32811 29767 32845
rect 29801 32811 29813 32845
rect 29755 32777 29813 32811
rect 29755 32743 29767 32777
rect 29801 32743 29813 32777
rect 29755 32709 29813 32743
rect 29755 32675 29767 32709
rect 29801 32675 29813 32709
rect 29755 32641 29813 32675
rect 29755 32607 29767 32641
rect 29801 32607 29813 32641
rect 29755 32573 29813 32607
rect 29755 32539 29767 32573
rect 29801 32539 29813 32573
rect 29755 32505 29813 32539
rect 29755 32471 29767 32505
rect 29801 32471 29813 32505
rect 29755 32437 29813 32471
rect 29755 32403 29767 32437
rect 29801 32403 29813 32437
rect 29755 32387 29813 32403
rect 30213 33661 30271 33677
rect 30213 33627 30225 33661
rect 30259 33627 30271 33661
rect 30213 33593 30271 33627
rect 30213 33559 30225 33593
rect 30259 33559 30271 33593
rect 30213 33525 30271 33559
rect 30213 33491 30225 33525
rect 30259 33491 30271 33525
rect 30213 33457 30271 33491
rect 30213 33423 30225 33457
rect 30259 33423 30271 33457
rect 30213 33389 30271 33423
rect 30213 33355 30225 33389
rect 30259 33355 30271 33389
rect 30213 33321 30271 33355
rect 30213 33287 30225 33321
rect 30259 33287 30271 33321
rect 30213 33253 30271 33287
rect 30213 33219 30225 33253
rect 30259 33219 30271 33253
rect 30213 33185 30271 33219
rect 30213 33151 30225 33185
rect 30259 33151 30271 33185
rect 30213 33117 30271 33151
rect 30213 33083 30225 33117
rect 30259 33083 30271 33117
rect 30213 33049 30271 33083
rect 30213 33015 30225 33049
rect 30259 33015 30271 33049
rect 30213 32981 30271 33015
rect 30213 32947 30225 32981
rect 30259 32947 30271 32981
rect 30213 32913 30271 32947
rect 30213 32879 30225 32913
rect 30259 32879 30271 32913
rect 30213 32845 30271 32879
rect 30213 32811 30225 32845
rect 30259 32811 30271 32845
rect 30213 32777 30271 32811
rect 30213 32743 30225 32777
rect 30259 32743 30271 32777
rect 30213 32709 30271 32743
rect 30213 32675 30225 32709
rect 30259 32675 30271 32709
rect 30213 32641 30271 32675
rect 30213 32607 30225 32641
rect 30259 32607 30271 32641
rect 30213 32573 30271 32607
rect 30213 32539 30225 32573
rect 30259 32539 30271 32573
rect 30213 32505 30271 32539
rect 30213 32471 30225 32505
rect 30259 32471 30271 32505
rect 30213 32437 30271 32471
rect 30213 32403 30225 32437
rect 30259 32403 30271 32437
rect 30213 32387 30271 32403
rect 30671 33661 30729 33677
rect 30671 33627 30683 33661
rect 30717 33627 30729 33661
rect 30671 33593 30729 33627
rect 30671 33559 30683 33593
rect 30717 33559 30729 33593
rect 30671 33525 30729 33559
rect 30671 33491 30683 33525
rect 30717 33491 30729 33525
rect 30671 33457 30729 33491
rect 30671 33423 30683 33457
rect 30717 33423 30729 33457
rect 30671 33389 30729 33423
rect 30671 33355 30683 33389
rect 30717 33355 30729 33389
rect 30671 33321 30729 33355
rect 30671 33287 30683 33321
rect 30717 33287 30729 33321
rect 30671 33253 30729 33287
rect 30671 33219 30683 33253
rect 30717 33219 30729 33253
rect 30671 33185 30729 33219
rect 30671 33151 30683 33185
rect 30717 33151 30729 33185
rect 30671 33117 30729 33151
rect 30671 33083 30683 33117
rect 30717 33083 30729 33117
rect 30671 33049 30729 33083
rect 30671 33015 30683 33049
rect 30717 33015 30729 33049
rect 30671 32981 30729 33015
rect 30671 32947 30683 32981
rect 30717 32947 30729 32981
rect 30671 32913 30729 32947
rect 30671 32879 30683 32913
rect 30717 32879 30729 32913
rect 30671 32845 30729 32879
rect 30671 32811 30683 32845
rect 30717 32811 30729 32845
rect 30671 32777 30729 32811
rect 30671 32743 30683 32777
rect 30717 32743 30729 32777
rect 30671 32709 30729 32743
rect 30671 32675 30683 32709
rect 30717 32675 30729 32709
rect 30671 32641 30729 32675
rect 30671 32607 30683 32641
rect 30717 32607 30729 32641
rect 30671 32573 30729 32607
rect 30671 32539 30683 32573
rect 30717 32539 30729 32573
rect 30671 32505 30729 32539
rect 30671 32471 30683 32505
rect 30717 32471 30729 32505
rect 30671 32437 30729 32471
rect 30671 32403 30683 32437
rect 30717 32403 30729 32437
rect 30671 32387 30729 32403
rect 31129 33661 31187 33677
rect 31129 33627 31141 33661
rect 31175 33627 31187 33661
rect 31129 33593 31187 33627
rect 31129 33559 31141 33593
rect 31175 33559 31187 33593
rect 31129 33525 31187 33559
rect 31129 33491 31141 33525
rect 31175 33491 31187 33525
rect 31129 33457 31187 33491
rect 31129 33423 31141 33457
rect 31175 33423 31187 33457
rect 31129 33389 31187 33423
rect 31129 33355 31141 33389
rect 31175 33355 31187 33389
rect 31129 33321 31187 33355
rect 31129 33287 31141 33321
rect 31175 33287 31187 33321
rect 31129 33253 31187 33287
rect 31129 33219 31141 33253
rect 31175 33219 31187 33253
rect 31129 33185 31187 33219
rect 31129 33151 31141 33185
rect 31175 33151 31187 33185
rect 31129 33117 31187 33151
rect 31129 33083 31141 33117
rect 31175 33083 31187 33117
rect 31129 33049 31187 33083
rect 31129 33015 31141 33049
rect 31175 33015 31187 33049
rect 31129 32981 31187 33015
rect 31129 32947 31141 32981
rect 31175 32947 31187 32981
rect 31129 32913 31187 32947
rect 31129 32879 31141 32913
rect 31175 32879 31187 32913
rect 31129 32845 31187 32879
rect 31129 32811 31141 32845
rect 31175 32811 31187 32845
rect 31129 32777 31187 32811
rect 31129 32743 31141 32777
rect 31175 32743 31187 32777
rect 31129 32709 31187 32743
rect 31129 32675 31141 32709
rect 31175 32675 31187 32709
rect 31129 32641 31187 32675
rect 31129 32607 31141 32641
rect 31175 32607 31187 32641
rect 31129 32573 31187 32607
rect 31129 32539 31141 32573
rect 31175 32539 31187 32573
rect 31129 32505 31187 32539
rect 31129 32471 31141 32505
rect 31175 32471 31187 32505
rect 31129 32437 31187 32471
rect 31129 32403 31141 32437
rect 31175 32403 31187 32437
rect 31129 32387 31187 32403
rect 31587 33661 31645 33677
rect 31587 33627 31599 33661
rect 31633 33627 31645 33661
rect 31587 33593 31645 33627
rect 31587 33559 31599 33593
rect 31633 33559 31645 33593
rect 31587 33525 31645 33559
rect 31587 33491 31599 33525
rect 31633 33491 31645 33525
rect 31587 33457 31645 33491
rect 31587 33423 31599 33457
rect 31633 33423 31645 33457
rect 31587 33389 31645 33423
rect 31587 33355 31599 33389
rect 31633 33355 31645 33389
rect 31587 33321 31645 33355
rect 31587 33287 31599 33321
rect 31633 33287 31645 33321
rect 31587 33253 31645 33287
rect 31587 33219 31599 33253
rect 31633 33219 31645 33253
rect 31587 33185 31645 33219
rect 31587 33151 31599 33185
rect 31633 33151 31645 33185
rect 31587 33117 31645 33151
rect 31587 33083 31599 33117
rect 31633 33083 31645 33117
rect 31587 33049 31645 33083
rect 31587 33015 31599 33049
rect 31633 33015 31645 33049
rect 31587 32981 31645 33015
rect 31587 32947 31599 32981
rect 31633 32947 31645 32981
rect 31587 32913 31645 32947
rect 31587 32879 31599 32913
rect 31633 32879 31645 32913
rect 31587 32845 31645 32879
rect 31587 32811 31599 32845
rect 31633 32811 31645 32845
rect 31587 32777 31645 32811
rect 31587 32743 31599 32777
rect 31633 32743 31645 32777
rect 31587 32709 31645 32743
rect 31587 32675 31599 32709
rect 31633 32675 31645 32709
rect 31587 32641 31645 32675
rect 31587 32607 31599 32641
rect 31633 32607 31645 32641
rect 31587 32573 31645 32607
rect 31587 32539 31599 32573
rect 31633 32539 31645 32573
rect 31587 32505 31645 32539
rect 31587 32471 31599 32505
rect 31633 32471 31645 32505
rect 31587 32437 31645 32471
rect 31587 32403 31599 32437
rect 31633 32403 31645 32437
rect 31587 32387 31645 32403
rect 32045 33661 32103 33677
rect 32045 33627 32057 33661
rect 32091 33627 32103 33661
rect 32045 33593 32103 33627
rect 32045 33559 32057 33593
rect 32091 33559 32103 33593
rect 32045 33525 32103 33559
rect 32045 33491 32057 33525
rect 32091 33491 32103 33525
rect 32045 33457 32103 33491
rect 32045 33423 32057 33457
rect 32091 33423 32103 33457
rect 32045 33389 32103 33423
rect 32045 33355 32057 33389
rect 32091 33355 32103 33389
rect 32045 33321 32103 33355
rect 32045 33287 32057 33321
rect 32091 33287 32103 33321
rect 32045 33253 32103 33287
rect 32045 33219 32057 33253
rect 32091 33219 32103 33253
rect 32045 33185 32103 33219
rect 32045 33151 32057 33185
rect 32091 33151 32103 33185
rect 32045 33117 32103 33151
rect 32045 33083 32057 33117
rect 32091 33083 32103 33117
rect 32045 33049 32103 33083
rect 32045 33015 32057 33049
rect 32091 33015 32103 33049
rect 32045 32981 32103 33015
rect 32045 32947 32057 32981
rect 32091 32947 32103 32981
rect 32045 32913 32103 32947
rect 32045 32879 32057 32913
rect 32091 32879 32103 32913
rect 32045 32845 32103 32879
rect 32045 32811 32057 32845
rect 32091 32811 32103 32845
rect 32045 32777 32103 32811
rect 32045 32743 32057 32777
rect 32091 32743 32103 32777
rect 32045 32709 32103 32743
rect 32045 32675 32057 32709
rect 32091 32675 32103 32709
rect 32045 32641 32103 32675
rect 32045 32607 32057 32641
rect 32091 32607 32103 32641
rect 32045 32573 32103 32607
rect 32045 32539 32057 32573
rect 32091 32539 32103 32573
rect 32045 32505 32103 32539
rect 32045 32471 32057 32505
rect 32091 32471 32103 32505
rect 32045 32437 32103 32471
rect 32045 32403 32057 32437
rect 32091 32403 32103 32437
rect 32045 32387 32103 32403
rect 32503 33661 32561 33677
rect 32503 33627 32515 33661
rect 32549 33627 32561 33661
rect 32503 33593 32561 33627
rect 32503 33559 32515 33593
rect 32549 33559 32561 33593
rect 32503 33525 32561 33559
rect 32503 33491 32515 33525
rect 32549 33491 32561 33525
rect 32503 33457 32561 33491
rect 32503 33423 32515 33457
rect 32549 33423 32561 33457
rect 32503 33389 32561 33423
rect 32503 33355 32515 33389
rect 32549 33355 32561 33389
rect 32503 33321 32561 33355
rect 32503 33287 32515 33321
rect 32549 33287 32561 33321
rect 32503 33253 32561 33287
rect 32503 33219 32515 33253
rect 32549 33219 32561 33253
rect 32503 33185 32561 33219
rect 32503 33151 32515 33185
rect 32549 33151 32561 33185
rect 32503 33117 32561 33151
rect 32503 33083 32515 33117
rect 32549 33083 32561 33117
rect 32503 33049 32561 33083
rect 32503 33015 32515 33049
rect 32549 33015 32561 33049
rect 32503 32981 32561 33015
rect 32503 32947 32515 32981
rect 32549 32947 32561 32981
rect 32503 32913 32561 32947
rect 32503 32879 32515 32913
rect 32549 32879 32561 32913
rect 32503 32845 32561 32879
rect 32503 32811 32515 32845
rect 32549 32811 32561 32845
rect 32503 32777 32561 32811
rect 32503 32743 32515 32777
rect 32549 32743 32561 32777
rect 32503 32709 32561 32743
rect 32503 32675 32515 32709
rect 32549 32675 32561 32709
rect 32503 32641 32561 32675
rect 32503 32607 32515 32641
rect 32549 32607 32561 32641
rect 32503 32573 32561 32607
rect 32503 32539 32515 32573
rect 32549 32539 32561 32573
rect 32503 32505 32561 32539
rect 32503 32471 32515 32505
rect 32549 32471 32561 32505
rect 32503 32437 32561 32471
rect 32503 32403 32515 32437
rect 32549 32403 32561 32437
rect 32503 32387 32561 32403
rect 32961 33661 33019 33677
rect 32961 33627 32973 33661
rect 33007 33627 33019 33661
rect 32961 33593 33019 33627
rect 32961 33559 32973 33593
rect 33007 33559 33019 33593
rect 32961 33525 33019 33559
rect 32961 33491 32973 33525
rect 33007 33491 33019 33525
rect 32961 33457 33019 33491
rect 32961 33423 32973 33457
rect 33007 33423 33019 33457
rect 32961 33389 33019 33423
rect 32961 33355 32973 33389
rect 33007 33355 33019 33389
rect 32961 33321 33019 33355
rect 32961 33287 32973 33321
rect 33007 33287 33019 33321
rect 32961 33253 33019 33287
rect 32961 33219 32973 33253
rect 33007 33219 33019 33253
rect 32961 33185 33019 33219
rect 32961 33151 32973 33185
rect 33007 33151 33019 33185
rect 32961 33117 33019 33151
rect 32961 33083 32973 33117
rect 33007 33083 33019 33117
rect 32961 33049 33019 33083
rect 32961 33015 32973 33049
rect 33007 33015 33019 33049
rect 32961 32981 33019 33015
rect 32961 32947 32973 32981
rect 33007 32947 33019 32981
rect 32961 32913 33019 32947
rect 32961 32879 32973 32913
rect 33007 32879 33019 32913
rect 32961 32845 33019 32879
rect 32961 32811 32973 32845
rect 33007 32811 33019 32845
rect 32961 32777 33019 32811
rect 32961 32743 32973 32777
rect 33007 32743 33019 32777
rect 32961 32709 33019 32743
rect 32961 32675 32973 32709
rect 33007 32675 33019 32709
rect 32961 32641 33019 32675
rect 32961 32607 32973 32641
rect 33007 32607 33019 32641
rect 32961 32573 33019 32607
rect 32961 32539 32973 32573
rect 33007 32539 33019 32573
rect 32961 32505 33019 32539
rect 32961 32471 32973 32505
rect 33007 32471 33019 32505
rect 32961 32437 33019 32471
rect 32961 32403 32973 32437
rect 33007 32403 33019 32437
rect 32961 32387 33019 32403
rect 33419 33661 33477 33677
rect 33419 33627 33431 33661
rect 33465 33627 33477 33661
rect 33419 33593 33477 33627
rect 33419 33559 33431 33593
rect 33465 33559 33477 33593
rect 33419 33525 33477 33559
rect 33419 33491 33431 33525
rect 33465 33491 33477 33525
rect 33419 33457 33477 33491
rect 33419 33423 33431 33457
rect 33465 33423 33477 33457
rect 33419 33389 33477 33423
rect 33419 33355 33431 33389
rect 33465 33355 33477 33389
rect 33419 33321 33477 33355
rect 33419 33287 33431 33321
rect 33465 33287 33477 33321
rect 33419 33253 33477 33287
rect 33419 33219 33431 33253
rect 33465 33219 33477 33253
rect 33419 33185 33477 33219
rect 33419 33151 33431 33185
rect 33465 33151 33477 33185
rect 33419 33117 33477 33151
rect 33419 33083 33431 33117
rect 33465 33083 33477 33117
rect 33419 33049 33477 33083
rect 33419 33015 33431 33049
rect 33465 33015 33477 33049
rect 33419 32981 33477 33015
rect 33419 32947 33431 32981
rect 33465 32947 33477 32981
rect 33419 32913 33477 32947
rect 33419 32879 33431 32913
rect 33465 32879 33477 32913
rect 33419 32845 33477 32879
rect 33419 32811 33431 32845
rect 33465 32811 33477 32845
rect 33419 32777 33477 32811
rect 33419 32743 33431 32777
rect 33465 32743 33477 32777
rect 33419 32709 33477 32743
rect 33419 32675 33431 32709
rect 33465 32675 33477 32709
rect 33419 32641 33477 32675
rect 33419 32607 33431 32641
rect 33465 32607 33477 32641
rect 33419 32573 33477 32607
rect 33419 32539 33431 32573
rect 33465 32539 33477 32573
rect 33419 32505 33477 32539
rect 33419 32471 33431 32505
rect 33465 32471 33477 32505
rect 33419 32437 33477 32471
rect 33419 32403 33431 32437
rect 33465 32403 33477 32437
rect 33419 32387 33477 32403
rect 33877 33661 33935 33677
rect 33877 33627 33889 33661
rect 33923 33627 33935 33661
rect 33877 33593 33935 33627
rect 33877 33559 33889 33593
rect 33923 33559 33935 33593
rect 33877 33525 33935 33559
rect 33877 33491 33889 33525
rect 33923 33491 33935 33525
rect 33877 33457 33935 33491
rect 33877 33423 33889 33457
rect 33923 33423 33935 33457
rect 33877 33389 33935 33423
rect 33877 33355 33889 33389
rect 33923 33355 33935 33389
rect 33877 33321 33935 33355
rect 33877 33287 33889 33321
rect 33923 33287 33935 33321
rect 33877 33253 33935 33287
rect 33877 33219 33889 33253
rect 33923 33219 33935 33253
rect 33877 33185 33935 33219
rect 33877 33151 33889 33185
rect 33923 33151 33935 33185
rect 33877 33117 33935 33151
rect 33877 33083 33889 33117
rect 33923 33083 33935 33117
rect 33877 33049 33935 33083
rect 33877 33015 33889 33049
rect 33923 33015 33935 33049
rect 33877 32981 33935 33015
rect 33877 32947 33889 32981
rect 33923 32947 33935 32981
rect 33877 32913 33935 32947
rect 33877 32879 33889 32913
rect 33923 32879 33935 32913
rect 33877 32845 33935 32879
rect 33877 32811 33889 32845
rect 33923 32811 33935 32845
rect 33877 32777 33935 32811
rect 33877 32743 33889 32777
rect 33923 32743 33935 32777
rect 33877 32709 33935 32743
rect 33877 32675 33889 32709
rect 33923 32675 33935 32709
rect 33877 32641 33935 32675
rect 33877 32607 33889 32641
rect 33923 32607 33935 32641
rect 33877 32573 33935 32607
rect 33877 32539 33889 32573
rect 33923 32539 33935 32573
rect 33877 32505 33935 32539
rect 33877 32471 33889 32505
rect 33923 32471 33935 32505
rect 33877 32437 33935 32471
rect 33877 32403 33889 32437
rect 33923 32403 33935 32437
rect 33877 32387 33935 32403
rect 34335 33661 34393 33677
rect 34335 33627 34347 33661
rect 34381 33627 34393 33661
rect 34335 33593 34393 33627
rect 34335 33559 34347 33593
rect 34381 33559 34393 33593
rect 34335 33525 34393 33559
rect 34335 33491 34347 33525
rect 34381 33491 34393 33525
rect 34335 33457 34393 33491
rect 34335 33423 34347 33457
rect 34381 33423 34393 33457
rect 34335 33389 34393 33423
rect 34335 33355 34347 33389
rect 34381 33355 34393 33389
rect 34335 33321 34393 33355
rect 34335 33287 34347 33321
rect 34381 33287 34393 33321
rect 34335 33253 34393 33287
rect 34335 33219 34347 33253
rect 34381 33219 34393 33253
rect 34335 33185 34393 33219
rect 34335 33151 34347 33185
rect 34381 33151 34393 33185
rect 34335 33117 34393 33151
rect 34335 33083 34347 33117
rect 34381 33083 34393 33117
rect 34335 33049 34393 33083
rect 34335 33015 34347 33049
rect 34381 33015 34393 33049
rect 34335 32981 34393 33015
rect 34335 32947 34347 32981
rect 34381 32947 34393 32981
rect 34335 32913 34393 32947
rect 34335 32879 34347 32913
rect 34381 32879 34393 32913
rect 34335 32845 34393 32879
rect 34335 32811 34347 32845
rect 34381 32811 34393 32845
rect 34335 32777 34393 32811
rect 34335 32743 34347 32777
rect 34381 32743 34393 32777
rect 34335 32709 34393 32743
rect 34335 32675 34347 32709
rect 34381 32675 34393 32709
rect 34335 32641 34393 32675
rect 34335 32607 34347 32641
rect 34381 32607 34393 32641
rect 34335 32573 34393 32607
rect 34335 32539 34347 32573
rect 34381 32539 34393 32573
rect 34335 32505 34393 32539
rect 34335 32471 34347 32505
rect 34381 32471 34393 32505
rect 34335 32437 34393 32471
rect 34335 32403 34347 32437
rect 34381 32403 34393 32437
rect 34335 32387 34393 32403
rect 34793 33661 34851 33677
rect 34793 33627 34805 33661
rect 34839 33627 34851 33661
rect 34793 33593 34851 33627
rect 34793 33559 34805 33593
rect 34839 33559 34851 33593
rect 34793 33525 34851 33559
rect 34793 33491 34805 33525
rect 34839 33491 34851 33525
rect 34793 33457 34851 33491
rect 34793 33423 34805 33457
rect 34839 33423 34851 33457
rect 34793 33389 34851 33423
rect 34793 33355 34805 33389
rect 34839 33355 34851 33389
rect 34793 33321 34851 33355
rect 34793 33287 34805 33321
rect 34839 33287 34851 33321
rect 34793 33253 34851 33287
rect 34793 33219 34805 33253
rect 34839 33219 34851 33253
rect 34793 33185 34851 33219
rect 34793 33151 34805 33185
rect 34839 33151 34851 33185
rect 34793 33117 34851 33151
rect 34793 33083 34805 33117
rect 34839 33083 34851 33117
rect 34793 33049 34851 33083
rect 34793 33015 34805 33049
rect 34839 33015 34851 33049
rect 34793 32981 34851 33015
rect 34793 32947 34805 32981
rect 34839 32947 34851 32981
rect 34793 32913 34851 32947
rect 34793 32879 34805 32913
rect 34839 32879 34851 32913
rect 34793 32845 34851 32879
rect 34793 32811 34805 32845
rect 34839 32811 34851 32845
rect 34793 32777 34851 32811
rect 34793 32743 34805 32777
rect 34839 32743 34851 32777
rect 34793 32709 34851 32743
rect 34793 32675 34805 32709
rect 34839 32675 34851 32709
rect 34793 32641 34851 32675
rect 34793 32607 34805 32641
rect 34839 32607 34851 32641
rect 34793 32573 34851 32607
rect 34793 32539 34805 32573
rect 34839 32539 34851 32573
rect 34793 32505 34851 32539
rect 34793 32471 34805 32505
rect 34839 32471 34851 32505
rect 34793 32437 34851 32471
rect 34793 32403 34805 32437
rect 34839 32403 34851 32437
rect 34793 32387 34851 32403
rect 35251 33661 35309 33677
rect 35251 33627 35263 33661
rect 35297 33627 35309 33661
rect 35251 33593 35309 33627
rect 35251 33559 35263 33593
rect 35297 33559 35309 33593
rect 35251 33525 35309 33559
rect 35251 33491 35263 33525
rect 35297 33491 35309 33525
rect 35251 33457 35309 33491
rect 35251 33423 35263 33457
rect 35297 33423 35309 33457
rect 35251 33389 35309 33423
rect 35251 33355 35263 33389
rect 35297 33355 35309 33389
rect 35251 33321 35309 33355
rect 35251 33287 35263 33321
rect 35297 33287 35309 33321
rect 35251 33253 35309 33287
rect 35251 33219 35263 33253
rect 35297 33219 35309 33253
rect 35251 33185 35309 33219
rect 35251 33151 35263 33185
rect 35297 33151 35309 33185
rect 35251 33117 35309 33151
rect 35251 33083 35263 33117
rect 35297 33083 35309 33117
rect 35251 33049 35309 33083
rect 35251 33015 35263 33049
rect 35297 33015 35309 33049
rect 35251 32981 35309 33015
rect 35251 32947 35263 32981
rect 35297 32947 35309 32981
rect 35251 32913 35309 32947
rect 35251 32879 35263 32913
rect 35297 32879 35309 32913
rect 35251 32845 35309 32879
rect 35251 32811 35263 32845
rect 35297 32811 35309 32845
rect 35251 32777 35309 32811
rect 35251 32743 35263 32777
rect 35297 32743 35309 32777
rect 35251 32709 35309 32743
rect 35251 32675 35263 32709
rect 35297 32675 35309 32709
rect 35251 32641 35309 32675
rect 35251 32607 35263 32641
rect 35297 32607 35309 32641
rect 35251 32573 35309 32607
rect 35251 32539 35263 32573
rect 35297 32539 35309 32573
rect 35251 32505 35309 32539
rect 35251 32471 35263 32505
rect 35297 32471 35309 32505
rect 35251 32437 35309 32471
rect 35251 32403 35263 32437
rect 35297 32403 35309 32437
rect 35251 32387 35309 32403
rect 35709 33661 35767 33677
rect 35709 33627 35721 33661
rect 35755 33627 35767 33661
rect 35709 33593 35767 33627
rect 35709 33559 35721 33593
rect 35755 33559 35767 33593
rect 35709 33525 35767 33559
rect 35709 33491 35721 33525
rect 35755 33491 35767 33525
rect 35709 33457 35767 33491
rect 35709 33423 35721 33457
rect 35755 33423 35767 33457
rect 35709 33389 35767 33423
rect 35709 33355 35721 33389
rect 35755 33355 35767 33389
rect 35709 33321 35767 33355
rect 35709 33287 35721 33321
rect 35755 33287 35767 33321
rect 35709 33253 35767 33287
rect 35709 33219 35721 33253
rect 35755 33219 35767 33253
rect 35709 33185 35767 33219
rect 35709 33151 35721 33185
rect 35755 33151 35767 33185
rect 35709 33117 35767 33151
rect 35709 33083 35721 33117
rect 35755 33083 35767 33117
rect 35709 33049 35767 33083
rect 35709 33015 35721 33049
rect 35755 33015 35767 33049
rect 35709 32981 35767 33015
rect 35709 32947 35721 32981
rect 35755 32947 35767 32981
rect 35709 32913 35767 32947
rect 35709 32879 35721 32913
rect 35755 32879 35767 32913
rect 35709 32845 35767 32879
rect 35709 32811 35721 32845
rect 35755 32811 35767 32845
rect 35709 32777 35767 32811
rect 35709 32743 35721 32777
rect 35755 32743 35767 32777
rect 35709 32709 35767 32743
rect 35709 32675 35721 32709
rect 35755 32675 35767 32709
rect 35709 32641 35767 32675
rect 35709 32607 35721 32641
rect 35755 32607 35767 32641
rect 35709 32573 35767 32607
rect 35709 32539 35721 32573
rect 35755 32539 35767 32573
rect 35709 32505 35767 32539
rect 35709 32471 35721 32505
rect 35755 32471 35767 32505
rect 35709 32437 35767 32471
rect 35709 32403 35721 32437
rect 35755 32403 35767 32437
rect 35709 32387 35767 32403
rect 36167 33661 36225 33677
rect 36167 33627 36179 33661
rect 36213 33627 36225 33661
rect 36167 33593 36225 33627
rect 36167 33559 36179 33593
rect 36213 33559 36225 33593
rect 36167 33525 36225 33559
rect 36167 33491 36179 33525
rect 36213 33491 36225 33525
rect 36167 33457 36225 33491
rect 36167 33423 36179 33457
rect 36213 33423 36225 33457
rect 36167 33389 36225 33423
rect 36167 33355 36179 33389
rect 36213 33355 36225 33389
rect 36167 33321 36225 33355
rect 36167 33287 36179 33321
rect 36213 33287 36225 33321
rect 36167 33253 36225 33287
rect 36167 33219 36179 33253
rect 36213 33219 36225 33253
rect 36167 33185 36225 33219
rect 36167 33151 36179 33185
rect 36213 33151 36225 33185
rect 36167 33117 36225 33151
rect 36167 33083 36179 33117
rect 36213 33083 36225 33117
rect 36167 33049 36225 33083
rect 36167 33015 36179 33049
rect 36213 33015 36225 33049
rect 36167 32981 36225 33015
rect 36167 32947 36179 32981
rect 36213 32947 36225 32981
rect 36167 32913 36225 32947
rect 36167 32879 36179 32913
rect 36213 32879 36225 32913
rect 36167 32845 36225 32879
rect 36167 32811 36179 32845
rect 36213 32811 36225 32845
rect 36167 32777 36225 32811
rect 36167 32743 36179 32777
rect 36213 32743 36225 32777
rect 36167 32709 36225 32743
rect 36167 32675 36179 32709
rect 36213 32675 36225 32709
rect 36167 32641 36225 32675
rect 36167 32607 36179 32641
rect 36213 32607 36225 32641
rect 36167 32573 36225 32607
rect 36167 32539 36179 32573
rect 36213 32539 36225 32573
rect 36167 32505 36225 32539
rect 36167 32471 36179 32505
rect 36213 32471 36225 32505
rect 36167 32437 36225 32471
rect 36167 32403 36179 32437
rect 36213 32403 36225 32437
rect 36167 32387 36225 32403
rect 36625 33661 36683 33677
rect 36625 33627 36637 33661
rect 36671 33627 36683 33661
rect 36625 33593 36683 33627
rect 36625 33559 36637 33593
rect 36671 33559 36683 33593
rect 36625 33525 36683 33559
rect 36625 33491 36637 33525
rect 36671 33491 36683 33525
rect 36625 33457 36683 33491
rect 36625 33423 36637 33457
rect 36671 33423 36683 33457
rect 36625 33389 36683 33423
rect 36625 33355 36637 33389
rect 36671 33355 36683 33389
rect 36625 33321 36683 33355
rect 36625 33287 36637 33321
rect 36671 33287 36683 33321
rect 36625 33253 36683 33287
rect 36625 33219 36637 33253
rect 36671 33219 36683 33253
rect 36625 33185 36683 33219
rect 36625 33151 36637 33185
rect 36671 33151 36683 33185
rect 36625 33117 36683 33151
rect 36625 33083 36637 33117
rect 36671 33083 36683 33117
rect 36625 33049 36683 33083
rect 36625 33015 36637 33049
rect 36671 33015 36683 33049
rect 36625 32981 36683 33015
rect 36625 32947 36637 32981
rect 36671 32947 36683 32981
rect 36625 32913 36683 32947
rect 36625 32879 36637 32913
rect 36671 32879 36683 32913
rect 36625 32845 36683 32879
rect 36625 32811 36637 32845
rect 36671 32811 36683 32845
rect 36625 32777 36683 32811
rect 36625 32743 36637 32777
rect 36671 32743 36683 32777
rect 36625 32709 36683 32743
rect 36625 32675 36637 32709
rect 36671 32675 36683 32709
rect 36625 32641 36683 32675
rect 36625 32607 36637 32641
rect 36671 32607 36683 32641
rect 36625 32573 36683 32607
rect 36625 32539 36637 32573
rect 36671 32539 36683 32573
rect 36625 32505 36683 32539
rect 36625 32471 36637 32505
rect 36671 32471 36683 32505
rect 36625 32437 36683 32471
rect 36625 32403 36637 32437
rect 36671 32403 36683 32437
rect 36625 32387 36683 32403
rect 37083 33661 37141 33677
rect 37083 33627 37095 33661
rect 37129 33627 37141 33661
rect 37083 33593 37141 33627
rect 37083 33559 37095 33593
rect 37129 33559 37141 33593
rect 37083 33525 37141 33559
rect 37083 33491 37095 33525
rect 37129 33491 37141 33525
rect 37083 33457 37141 33491
rect 37083 33423 37095 33457
rect 37129 33423 37141 33457
rect 37083 33389 37141 33423
rect 37083 33355 37095 33389
rect 37129 33355 37141 33389
rect 37083 33321 37141 33355
rect 37083 33287 37095 33321
rect 37129 33287 37141 33321
rect 37083 33253 37141 33287
rect 37083 33219 37095 33253
rect 37129 33219 37141 33253
rect 37083 33185 37141 33219
rect 37083 33151 37095 33185
rect 37129 33151 37141 33185
rect 37083 33117 37141 33151
rect 37083 33083 37095 33117
rect 37129 33083 37141 33117
rect 37083 33049 37141 33083
rect 37083 33015 37095 33049
rect 37129 33015 37141 33049
rect 37083 32981 37141 33015
rect 37083 32947 37095 32981
rect 37129 32947 37141 32981
rect 37083 32913 37141 32947
rect 37083 32879 37095 32913
rect 37129 32879 37141 32913
rect 37083 32845 37141 32879
rect 37083 32811 37095 32845
rect 37129 32811 37141 32845
rect 37083 32777 37141 32811
rect 37083 32743 37095 32777
rect 37129 32743 37141 32777
rect 37083 32709 37141 32743
rect 37083 32675 37095 32709
rect 37129 32675 37141 32709
rect 37083 32641 37141 32675
rect 37083 32607 37095 32641
rect 37129 32607 37141 32641
rect 37083 32573 37141 32607
rect 37083 32539 37095 32573
rect 37129 32539 37141 32573
rect 37083 32505 37141 32539
rect 37083 32471 37095 32505
rect 37129 32471 37141 32505
rect 37083 32437 37141 32471
rect 37083 32403 37095 32437
rect 37129 32403 37141 32437
rect 37083 32387 37141 32403
rect 37541 33661 37599 33677
rect 37541 33627 37553 33661
rect 37587 33627 37599 33661
rect 37541 33593 37599 33627
rect 37541 33559 37553 33593
rect 37587 33559 37599 33593
rect 37541 33525 37599 33559
rect 37541 33491 37553 33525
rect 37587 33491 37599 33525
rect 37541 33457 37599 33491
rect 37541 33423 37553 33457
rect 37587 33423 37599 33457
rect 37541 33389 37599 33423
rect 37541 33355 37553 33389
rect 37587 33355 37599 33389
rect 37541 33321 37599 33355
rect 37541 33287 37553 33321
rect 37587 33287 37599 33321
rect 37541 33253 37599 33287
rect 37541 33219 37553 33253
rect 37587 33219 37599 33253
rect 37541 33185 37599 33219
rect 37541 33151 37553 33185
rect 37587 33151 37599 33185
rect 37541 33117 37599 33151
rect 37541 33083 37553 33117
rect 37587 33083 37599 33117
rect 37541 33049 37599 33083
rect 37541 33015 37553 33049
rect 37587 33015 37599 33049
rect 37541 32981 37599 33015
rect 37541 32947 37553 32981
rect 37587 32947 37599 32981
rect 37541 32913 37599 32947
rect 37541 32879 37553 32913
rect 37587 32879 37599 32913
rect 37541 32845 37599 32879
rect 37541 32811 37553 32845
rect 37587 32811 37599 32845
rect 37541 32777 37599 32811
rect 37541 32743 37553 32777
rect 37587 32743 37599 32777
rect 37541 32709 37599 32743
rect 37541 32675 37553 32709
rect 37587 32675 37599 32709
rect 37541 32641 37599 32675
rect 37541 32607 37553 32641
rect 37587 32607 37599 32641
rect 37541 32573 37599 32607
rect 37541 32539 37553 32573
rect 37587 32539 37599 32573
rect 37541 32505 37599 32539
rect 37541 32471 37553 32505
rect 37587 32471 37599 32505
rect 37541 32437 37599 32471
rect 37541 32403 37553 32437
rect 37587 32403 37599 32437
rect 37541 32387 37599 32403
rect 37999 33661 38057 33677
rect 37999 33627 38011 33661
rect 38045 33627 38057 33661
rect 37999 33593 38057 33627
rect 37999 33559 38011 33593
rect 38045 33559 38057 33593
rect 37999 33525 38057 33559
rect 37999 33491 38011 33525
rect 38045 33491 38057 33525
rect 37999 33457 38057 33491
rect 37999 33423 38011 33457
rect 38045 33423 38057 33457
rect 37999 33389 38057 33423
rect 37999 33355 38011 33389
rect 38045 33355 38057 33389
rect 37999 33321 38057 33355
rect 37999 33287 38011 33321
rect 38045 33287 38057 33321
rect 37999 33253 38057 33287
rect 37999 33219 38011 33253
rect 38045 33219 38057 33253
rect 37999 33185 38057 33219
rect 37999 33151 38011 33185
rect 38045 33151 38057 33185
rect 37999 33117 38057 33151
rect 37999 33083 38011 33117
rect 38045 33083 38057 33117
rect 37999 33049 38057 33083
rect 37999 33015 38011 33049
rect 38045 33015 38057 33049
rect 37999 32981 38057 33015
rect 37999 32947 38011 32981
rect 38045 32947 38057 32981
rect 37999 32913 38057 32947
rect 37999 32879 38011 32913
rect 38045 32879 38057 32913
rect 37999 32845 38057 32879
rect 37999 32811 38011 32845
rect 38045 32811 38057 32845
rect 37999 32777 38057 32811
rect 37999 32743 38011 32777
rect 38045 32743 38057 32777
rect 37999 32709 38057 32743
rect 37999 32675 38011 32709
rect 38045 32675 38057 32709
rect 37999 32641 38057 32675
rect 37999 32607 38011 32641
rect 38045 32607 38057 32641
rect 37999 32573 38057 32607
rect 37999 32539 38011 32573
rect 38045 32539 38057 32573
rect 37999 32505 38057 32539
rect 37999 32471 38011 32505
rect 38045 32471 38057 32505
rect 37999 32437 38057 32471
rect 37999 32403 38011 32437
rect 38045 32403 38057 32437
rect 37999 32387 38057 32403
rect 38457 33661 38515 33677
rect 38457 33627 38469 33661
rect 38503 33627 38515 33661
rect 38457 33593 38515 33627
rect 38457 33559 38469 33593
rect 38503 33559 38515 33593
rect 38457 33525 38515 33559
rect 38457 33491 38469 33525
rect 38503 33491 38515 33525
rect 38457 33457 38515 33491
rect 38457 33423 38469 33457
rect 38503 33423 38515 33457
rect 38457 33389 38515 33423
rect 38457 33355 38469 33389
rect 38503 33355 38515 33389
rect 38457 33321 38515 33355
rect 38457 33287 38469 33321
rect 38503 33287 38515 33321
rect 38457 33253 38515 33287
rect 38457 33219 38469 33253
rect 38503 33219 38515 33253
rect 38457 33185 38515 33219
rect 38457 33151 38469 33185
rect 38503 33151 38515 33185
rect 38457 33117 38515 33151
rect 38457 33083 38469 33117
rect 38503 33083 38515 33117
rect 38457 33049 38515 33083
rect 38457 33015 38469 33049
rect 38503 33015 38515 33049
rect 38457 32981 38515 33015
rect 38457 32947 38469 32981
rect 38503 32947 38515 32981
rect 38457 32913 38515 32947
rect 38457 32879 38469 32913
rect 38503 32879 38515 32913
rect 38457 32845 38515 32879
rect 38457 32811 38469 32845
rect 38503 32811 38515 32845
rect 38457 32777 38515 32811
rect 38457 32743 38469 32777
rect 38503 32743 38515 32777
rect 38457 32709 38515 32743
rect 38457 32675 38469 32709
rect 38503 32675 38515 32709
rect 38457 32641 38515 32675
rect 38457 32607 38469 32641
rect 38503 32607 38515 32641
rect 38457 32573 38515 32607
rect 38457 32539 38469 32573
rect 38503 32539 38515 32573
rect 38457 32505 38515 32539
rect 38457 32471 38469 32505
rect 38503 32471 38515 32505
rect 38457 32437 38515 32471
rect 38457 32403 38469 32437
rect 38503 32403 38515 32437
rect 38457 32387 38515 32403
rect 38915 33661 38973 33677
rect 38915 33627 38927 33661
rect 38961 33627 38973 33661
rect 38915 33593 38973 33627
rect 38915 33559 38927 33593
rect 38961 33559 38973 33593
rect 38915 33525 38973 33559
rect 38915 33491 38927 33525
rect 38961 33491 38973 33525
rect 38915 33457 38973 33491
rect 38915 33423 38927 33457
rect 38961 33423 38973 33457
rect 38915 33389 38973 33423
rect 38915 33355 38927 33389
rect 38961 33355 38973 33389
rect 38915 33321 38973 33355
rect 38915 33287 38927 33321
rect 38961 33287 38973 33321
rect 38915 33253 38973 33287
rect 38915 33219 38927 33253
rect 38961 33219 38973 33253
rect 38915 33185 38973 33219
rect 38915 33151 38927 33185
rect 38961 33151 38973 33185
rect 38915 33117 38973 33151
rect 38915 33083 38927 33117
rect 38961 33083 38973 33117
rect 38915 33049 38973 33083
rect 38915 33015 38927 33049
rect 38961 33015 38973 33049
rect 38915 32981 38973 33015
rect 38915 32947 38927 32981
rect 38961 32947 38973 32981
rect 38915 32913 38973 32947
rect 38915 32879 38927 32913
rect 38961 32879 38973 32913
rect 38915 32845 38973 32879
rect 38915 32811 38927 32845
rect 38961 32811 38973 32845
rect 38915 32777 38973 32811
rect 38915 32743 38927 32777
rect 38961 32743 38973 32777
rect 38915 32709 38973 32743
rect 38915 32675 38927 32709
rect 38961 32675 38973 32709
rect 38915 32641 38973 32675
rect 38915 32607 38927 32641
rect 38961 32607 38973 32641
rect 38915 32573 38973 32607
rect 38915 32539 38927 32573
rect 38961 32539 38973 32573
rect 38915 32505 38973 32539
rect 38915 32471 38927 32505
rect 38961 32471 38973 32505
rect 38915 32437 38973 32471
rect 38915 32403 38927 32437
rect 38961 32403 38973 32437
rect 38915 32387 38973 32403
rect 39373 33661 39431 33677
rect 39373 33627 39385 33661
rect 39419 33627 39431 33661
rect 39373 33593 39431 33627
rect 39373 33559 39385 33593
rect 39419 33559 39431 33593
rect 39373 33525 39431 33559
rect 39373 33491 39385 33525
rect 39419 33491 39431 33525
rect 39373 33457 39431 33491
rect 39373 33423 39385 33457
rect 39419 33423 39431 33457
rect 39373 33389 39431 33423
rect 39373 33355 39385 33389
rect 39419 33355 39431 33389
rect 39373 33321 39431 33355
rect 39373 33287 39385 33321
rect 39419 33287 39431 33321
rect 39373 33253 39431 33287
rect 39373 33219 39385 33253
rect 39419 33219 39431 33253
rect 39373 33185 39431 33219
rect 39373 33151 39385 33185
rect 39419 33151 39431 33185
rect 39373 33117 39431 33151
rect 39373 33083 39385 33117
rect 39419 33083 39431 33117
rect 39373 33049 39431 33083
rect 39373 33015 39385 33049
rect 39419 33015 39431 33049
rect 39373 32981 39431 33015
rect 39373 32947 39385 32981
rect 39419 32947 39431 32981
rect 39373 32913 39431 32947
rect 39373 32879 39385 32913
rect 39419 32879 39431 32913
rect 39373 32845 39431 32879
rect 39373 32811 39385 32845
rect 39419 32811 39431 32845
rect 39373 32777 39431 32811
rect 39373 32743 39385 32777
rect 39419 32743 39431 32777
rect 39373 32709 39431 32743
rect 39373 32675 39385 32709
rect 39419 32675 39431 32709
rect 39373 32641 39431 32675
rect 39373 32607 39385 32641
rect 39419 32607 39431 32641
rect 39373 32573 39431 32607
rect 39373 32539 39385 32573
rect 39419 32539 39431 32573
rect 39373 32505 39431 32539
rect 39373 32471 39385 32505
rect 39419 32471 39431 32505
rect 39373 32437 39431 32471
rect 39373 32403 39385 32437
rect 39419 32403 39431 32437
rect 39373 32387 39431 32403
rect 39831 33661 39889 33677
rect 39831 33627 39843 33661
rect 39877 33627 39889 33661
rect 39831 33593 39889 33627
rect 39831 33559 39843 33593
rect 39877 33559 39889 33593
rect 39831 33525 39889 33559
rect 39831 33491 39843 33525
rect 39877 33491 39889 33525
rect 39831 33457 39889 33491
rect 39831 33423 39843 33457
rect 39877 33423 39889 33457
rect 39831 33389 39889 33423
rect 39831 33355 39843 33389
rect 39877 33355 39889 33389
rect 39831 33321 39889 33355
rect 39831 33287 39843 33321
rect 39877 33287 39889 33321
rect 39831 33253 39889 33287
rect 39831 33219 39843 33253
rect 39877 33219 39889 33253
rect 39831 33185 39889 33219
rect 39831 33151 39843 33185
rect 39877 33151 39889 33185
rect 39831 33117 39889 33151
rect 39831 33083 39843 33117
rect 39877 33083 39889 33117
rect 39831 33049 39889 33083
rect 39831 33015 39843 33049
rect 39877 33015 39889 33049
rect 39831 32981 39889 33015
rect 39831 32947 39843 32981
rect 39877 32947 39889 32981
rect 39831 32913 39889 32947
rect 39831 32879 39843 32913
rect 39877 32879 39889 32913
rect 39831 32845 39889 32879
rect 39831 32811 39843 32845
rect 39877 32811 39889 32845
rect 39831 32777 39889 32811
rect 39831 32743 39843 32777
rect 39877 32743 39889 32777
rect 39831 32709 39889 32743
rect 39831 32675 39843 32709
rect 39877 32675 39889 32709
rect 39831 32641 39889 32675
rect 39831 32607 39843 32641
rect 39877 32607 39889 32641
rect 39831 32573 39889 32607
rect 39831 32539 39843 32573
rect 39877 32539 39889 32573
rect 39831 32505 39889 32539
rect 39831 32471 39843 32505
rect 39877 32471 39889 32505
rect 39831 32437 39889 32471
rect 39831 32403 39843 32437
rect 39877 32403 39889 32437
rect 39831 32387 39889 32403
rect 40289 33661 40347 33677
rect 40289 33627 40301 33661
rect 40335 33627 40347 33661
rect 40289 33593 40347 33627
rect 40289 33559 40301 33593
rect 40335 33559 40347 33593
rect 40289 33525 40347 33559
rect 40289 33491 40301 33525
rect 40335 33491 40347 33525
rect 40289 33457 40347 33491
rect 40289 33423 40301 33457
rect 40335 33423 40347 33457
rect 40289 33389 40347 33423
rect 40289 33355 40301 33389
rect 40335 33355 40347 33389
rect 40289 33321 40347 33355
rect 40289 33287 40301 33321
rect 40335 33287 40347 33321
rect 40289 33253 40347 33287
rect 40289 33219 40301 33253
rect 40335 33219 40347 33253
rect 40289 33185 40347 33219
rect 40289 33151 40301 33185
rect 40335 33151 40347 33185
rect 40289 33117 40347 33151
rect 40289 33083 40301 33117
rect 40335 33083 40347 33117
rect 40289 33049 40347 33083
rect 40289 33015 40301 33049
rect 40335 33015 40347 33049
rect 40289 32981 40347 33015
rect 40289 32947 40301 32981
rect 40335 32947 40347 32981
rect 40289 32913 40347 32947
rect 40289 32879 40301 32913
rect 40335 32879 40347 32913
rect 40289 32845 40347 32879
rect 40289 32811 40301 32845
rect 40335 32811 40347 32845
rect 40289 32777 40347 32811
rect 40289 32743 40301 32777
rect 40335 32743 40347 32777
rect 40289 32709 40347 32743
rect 40289 32675 40301 32709
rect 40335 32675 40347 32709
rect 40289 32641 40347 32675
rect 40289 32607 40301 32641
rect 40335 32607 40347 32641
rect 40289 32573 40347 32607
rect 40289 32539 40301 32573
rect 40335 32539 40347 32573
rect 40289 32505 40347 32539
rect 40289 32471 40301 32505
rect 40335 32471 40347 32505
rect 40289 32437 40347 32471
rect 40289 32403 40301 32437
rect 40335 32403 40347 32437
rect 40289 32387 40347 32403
rect 40747 33661 40805 33677
rect 40747 33627 40759 33661
rect 40793 33627 40805 33661
rect 40747 33593 40805 33627
rect 40747 33559 40759 33593
rect 40793 33559 40805 33593
rect 40747 33525 40805 33559
rect 40747 33491 40759 33525
rect 40793 33491 40805 33525
rect 40747 33457 40805 33491
rect 40747 33423 40759 33457
rect 40793 33423 40805 33457
rect 40747 33389 40805 33423
rect 40747 33355 40759 33389
rect 40793 33355 40805 33389
rect 40747 33321 40805 33355
rect 40747 33287 40759 33321
rect 40793 33287 40805 33321
rect 40747 33253 40805 33287
rect 40747 33219 40759 33253
rect 40793 33219 40805 33253
rect 40747 33185 40805 33219
rect 40747 33151 40759 33185
rect 40793 33151 40805 33185
rect 40747 33117 40805 33151
rect 40747 33083 40759 33117
rect 40793 33083 40805 33117
rect 40747 33049 40805 33083
rect 40747 33015 40759 33049
rect 40793 33015 40805 33049
rect 40747 32981 40805 33015
rect 40747 32947 40759 32981
rect 40793 32947 40805 32981
rect 40747 32913 40805 32947
rect 40747 32879 40759 32913
rect 40793 32879 40805 32913
rect 40747 32845 40805 32879
rect 40747 32811 40759 32845
rect 40793 32811 40805 32845
rect 40747 32777 40805 32811
rect 40747 32743 40759 32777
rect 40793 32743 40805 32777
rect 40747 32709 40805 32743
rect 40747 32675 40759 32709
rect 40793 32675 40805 32709
rect 40747 32641 40805 32675
rect 40747 32607 40759 32641
rect 40793 32607 40805 32641
rect 40747 32573 40805 32607
rect 40747 32539 40759 32573
rect 40793 32539 40805 32573
rect 40747 32505 40805 32539
rect 40747 32471 40759 32505
rect 40793 32471 40805 32505
rect 40747 32437 40805 32471
rect 40747 32403 40759 32437
rect 40793 32403 40805 32437
rect 40747 32387 40805 32403
rect 41205 33661 41263 33677
rect 41205 33627 41217 33661
rect 41251 33627 41263 33661
rect 41205 33593 41263 33627
rect 41205 33559 41217 33593
rect 41251 33559 41263 33593
rect 41205 33525 41263 33559
rect 41205 33491 41217 33525
rect 41251 33491 41263 33525
rect 41205 33457 41263 33491
rect 41205 33423 41217 33457
rect 41251 33423 41263 33457
rect 41205 33389 41263 33423
rect 41205 33355 41217 33389
rect 41251 33355 41263 33389
rect 41205 33321 41263 33355
rect 41205 33287 41217 33321
rect 41251 33287 41263 33321
rect 41205 33253 41263 33287
rect 41205 33219 41217 33253
rect 41251 33219 41263 33253
rect 41205 33185 41263 33219
rect 41205 33151 41217 33185
rect 41251 33151 41263 33185
rect 41205 33117 41263 33151
rect 41205 33083 41217 33117
rect 41251 33083 41263 33117
rect 41205 33049 41263 33083
rect 41205 33015 41217 33049
rect 41251 33015 41263 33049
rect 41205 32981 41263 33015
rect 41205 32947 41217 32981
rect 41251 32947 41263 32981
rect 41205 32913 41263 32947
rect 41205 32879 41217 32913
rect 41251 32879 41263 32913
rect 41205 32845 41263 32879
rect 41205 32811 41217 32845
rect 41251 32811 41263 32845
rect 41205 32777 41263 32811
rect 41205 32743 41217 32777
rect 41251 32743 41263 32777
rect 41205 32709 41263 32743
rect 41205 32675 41217 32709
rect 41251 32675 41263 32709
rect 41205 32641 41263 32675
rect 41205 32607 41217 32641
rect 41251 32607 41263 32641
rect 41205 32573 41263 32607
rect 41205 32539 41217 32573
rect 41251 32539 41263 32573
rect 41205 32505 41263 32539
rect 41205 32471 41217 32505
rect 41251 32471 41263 32505
rect 41205 32437 41263 32471
rect 41205 32403 41217 32437
rect 41251 32403 41263 32437
rect 41205 32387 41263 32403
rect 41663 33661 41721 33677
rect 41663 33627 41675 33661
rect 41709 33627 41721 33661
rect 41663 33593 41721 33627
rect 41663 33559 41675 33593
rect 41709 33559 41721 33593
rect 41663 33525 41721 33559
rect 41663 33491 41675 33525
rect 41709 33491 41721 33525
rect 41663 33457 41721 33491
rect 41663 33423 41675 33457
rect 41709 33423 41721 33457
rect 41663 33389 41721 33423
rect 41663 33355 41675 33389
rect 41709 33355 41721 33389
rect 41663 33321 41721 33355
rect 41663 33287 41675 33321
rect 41709 33287 41721 33321
rect 41663 33253 41721 33287
rect 41663 33219 41675 33253
rect 41709 33219 41721 33253
rect 41663 33185 41721 33219
rect 41663 33151 41675 33185
rect 41709 33151 41721 33185
rect 41663 33117 41721 33151
rect 41663 33083 41675 33117
rect 41709 33083 41721 33117
rect 41663 33049 41721 33083
rect 41663 33015 41675 33049
rect 41709 33015 41721 33049
rect 41663 32981 41721 33015
rect 41663 32947 41675 32981
rect 41709 32947 41721 32981
rect 41663 32913 41721 32947
rect 41663 32879 41675 32913
rect 41709 32879 41721 32913
rect 41663 32845 41721 32879
rect 41663 32811 41675 32845
rect 41709 32811 41721 32845
rect 41663 32777 41721 32811
rect 41663 32743 41675 32777
rect 41709 32743 41721 32777
rect 41663 32709 41721 32743
rect 41663 32675 41675 32709
rect 41709 32675 41721 32709
rect 41663 32641 41721 32675
rect 41663 32607 41675 32641
rect 41709 32607 41721 32641
rect 41663 32573 41721 32607
rect 41663 32539 41675 32573
rect 41709 32539 41721 32573
rect 41663 32505 41721 32539
rect 41663 32471 41675 32505
rect 41709 32471 41721 32505
rect 41663 32437 41721 32471
rect 41663 32403 41675 32437
rect 41709 32403 41721 32437
rect 41663 32387 41721 32403
rect 6049 29901 6107 29917
rect 6049 29867 6061 29901
rect 6095 29867 6107 29901
rect 6049 29833 6107 29867
rect 6049 29799 6061 29833
rect 6095 29799 6107 29833
rect 6049 29765 6107 29799
rect 6049 29731 6061 29765
rect 6095 29731 6107 29765
rect 6049 29697 6107 29731
rect 6049 29663 6061 29697
rect 6095 29663 6107 29697
rect 6049 29629 6107 29663
rect 6049 29595 6061 29629
rect 6095 29595 6107 29629
rect 6049 29561 6107 29595
rect 6049 29527 6061 29561
rect 6095 29527 6107 29561
rect 6049 29493 6107 29527
rect 6049 29459 6061 29493
rect 6095 29459 6107 29493
rect 6049 29425 6107 29459
rect 6049 29391 6061 29425
rect 6095 29391 6107 29425
rect 6049 29357 6107 29391
rect 6049 29323 6061 29357
rect 6095 29323 6107 29357
rect 6049 29289 6107 29323
rect 6049 29255 6061 29289
rect 6095 29255 6107 29289
rect 6049 29221 6107 29255
rect 6049 29187 6061 29221
rect 6095 29187 6107 29221
rect 6049 29153 6107 29187
rect 6049 29119 6061 29153
rect 6095 29119 6107 29153
rect 6049 29085 6107 29119
rect 6049 29051 6061 29085
rect 6095 29051 6107 29085
rect 6049 29017 6107 29051
rect 6049 28983 6061 29017
rect 6095 28983 6107 29017
rect 6049 28949 6107 28983
rect 6049 28915 6061 28949
rect 6095 28915 6107 28949
rect 6049 28881 6107 28915
rect 6049 28847 6061 28881
rect 6095 28847 6107 28881
rect 6049 28813 6107 28847
rect 6049 28779 6061 28813
rect 6095 28779 6107 28813
rect 6049 28745 6107 28779
rect 6049 28711 6061 28745
rect 6095 28711 6107 28745
rect 6049 28677 6107 28711
rect 6049 28643 6061 28677
rect 6095 28643 6107 28677
rect 6049 28627 6107 28643
rect 6507 29901 6565 29917
rect 6507 29867 6519 29901
rect 6553 29867 6565 29901
rect 6507 29833 6565 29867
rect 6507 29799 6519 29833
rect 6553 29799 6565 29833
rect 6507 29765 6565 29799
rect 6507 29731 6519 29765
rect 6553 29731 6565 29765
rect 6507 29697 6565 29731
rect 6507 29663 6519 29697
rect 6553 29663 6565 29697
rect 6507 29629 6565 29663
rect 6507 29595 6519 29629
rect 6553 29595 6565 29629
rect 6507 29561 6565 29595
rect 6507 29527 6519 29561
rect 6553 29527 6565 29561
rect 6507 29493 6565 29527
rect 6507 29459 6519 29493
rect 6553 29459 6565 29493
rect 6507 29425 6565 29459
rect 6507 29391 6519 29425
rect 6553 29391 6565 29425
rect 6507 29357 6565 29391
rect 6507 29323 6519 29357
rect 6553 29323 6565 29357
rect 6507 29289 6565 29323
rect 6507 29255 6519 29289
rect 6553 29255 6565 29289
rect 6507 29221 6565 29255
rect 6507 29187 6519 29221
rect 6553 29187 6565 29221
rect 6507 29153 6565 29187
rect 6507 29119 6519 29153
rect 6553 29119 6565 29153
rect 6507 29085 6565 29119
rect 6507 29051 6519 29085
rect 6553 29051 6565 29085
rect 6507 29017 6565 29051
rect 6507 28983 6519 29017
rect 6553 28983 6565 29017
rect 6507 28949 6565 28983
rect 6507 28915 6519 28949
rect 6553 28915 6565 28949
rect 6507 28881 6565 28915
rect 6507 28847 6519 28881
rect 6553 28847 6565 28881
rect 6507 28813 6565 28847
rect 6507 28779 6519 28813
rect 6553 28779 6565 28813
rect 6507 28745 6565 28779
rect 6507 28711 6519 28745
rect 6553 28711 6565 28745
rect 6507 28677 6565 28711
rect 6507 28643 6519 28677
rect 6553 28643 6565 28677
rect 6507 28627 6565 28643
rect 6965 29901 7023 29917
rect 6965 29867 6977 29901
rect 7011 29867 7023 29901
rect 6965 29833 7023 29867
rect 6965 29799 6977 29833
rect 7011 29799 7023 29833
rect 6965 29765 7023 29799
rect 6965 29731 6977 29765
rect 7011 29731 7023 29765
rect 6965 29697 7023 29731
rect 6965 29663 6977 29697
rect 7011 29663 7023 29697
rect 6965 29629 7023 29663
rect 6965 29595 6977 29629
rect 7011 29595 7023 29629
rect 6965 29561 7023 29595
rect 6965 29527 6977 29561
rect 7011 29527 7023 29561
rect 6965 29493 7023 29527
rect 6965 29459 6977 29493
rect 7011 29459 7023 29493
rect 6965 29425 7023 29459
rect 6965 29391 6977 29425
rect 7011 29391 7023 29425
rect 6965 29357 7023 29391
rect 6965 29323 6977 29357
rect 7011 29323 7023 29357
rect 6965 29289 7023 29323
rect 6965 29255 6977 29289
rect 7011 29255 7023 29289
rect 6965 29221 7023 29255
rect 6965 29187 6977 29221
rect 7011 29187 7023 29221
rect 6965 29153 7023 29187
rect 6965 29119 6977 29153
rect 7011 29119 7023 29153
rect 6965 29085 7023 29119
rect 6965 29051 6977 29085
rect 7011 29051 7023 29085
rect 6965 29017 7023 29051
rect 6965 28983 6977 29017
rect 7011 28983 7023 29017
rect 6965 28949 7023 28983
rect 6965 28915 6977 28949
rect 7011 28915 7023 28949
rect 6965 28881 7023 28915
rect 6965 28847 6977 28881
rect 7011 28847 7023 28881
rect 6965 28813 7023 28847
rect 6965 28779 6977 28813
rect 7011 28779 7023 28813
rect 6965 28745 7023 28779
rect 6965 28711 6977 28745
rect 7011 28711 7023 28745
rect 6965 28677 7023 28711
rect 6965 28643 6977 28677
rect 7011 28643 7023 28677
rect 6965 28627 7023 28643
rect 7423 29901 7481 29917
rect 7423 29867 7435 29901
rect 7469 29867 7481 29901
rect 7423 29833 7481 29867
rect 7423 29799 7435 29833
rect 7469 29799 7481 29833
rect 7423 29765 7481 29799
rect 7423 29731 7435 29765
rect 7469 29731 7481 29765
rect 7423 29697 7481 29731
rect 7423 29663 7435 29697
rect 7469 29663 7481 29697
rect 7423 29629 7481 29663
rect 7423 29595 7435 29629
rect 7469 29595 7481 29629
rect 7423 29561 7481 29595
rect 7423 29527 7435 29561
rect 7469 29527 7481 29561
rect 7423 29493 7481 29527
rect 7423 29459 7435 29493
rect 7469 29459 7481 29493
rect 7423 29425 7481 29459
rect 7423 29391 7435 29425
rect 7469 29391 7481 29425
rect 7423 29357 7481 29391
rect 7423 29323 7435 29357
rect 7469 29323 7481 29357
rect 7423 29289 7481 29323
rect 7423 29255 7435 29289
rect 7469 29255 7481 29289
rect 7423 29221 7481 29255
rect 7423 29187 7435 29221
rect 7469 29187 7481 29221
rect 7423 29153 7481 29187
rect 7423 29119 7435 29153
rect 7469 29119 7481 29153
rect 7423 29085 7481 29119
rect 7423 29051 7435 29085
rect 7469 29051 7481 29085
rect 7423 29017 7481 29051
rect 7423 28983 7435 29017
rect 7469 28983 7481 29017
rect 7423 28949 7481 28983
rect 7423 28915 7435 28949
rect 7469 28915 7481 28949
rect 7423 28881 7481 28915
rect 7423 28847 7435 28881
rect 7469 28847 7481 28881
rect 7423 28813 7481 28847
rect 7423 28779 7435 28813
rect 7469 28779 7481 28813
rect 7423 28745 7481 28779
rect 7423 28711 7435 28745
rect 7469 28711 7481 28745
rect 7423 28677 7481 28711
rect 7423 28643 7435 28677
rect 7469 28643 7481 28677
rect 7423 28627 7481 28643
rect 7881 29901 7939 29917
rect 7881 29867 7893 29901
rect 7927 29867 7939 29901
rect 7881 29833 7939 29867
rect 7881 29799 7893 29833
rect 7927 29799 7939 29833
rect 7881 29765 7939 29799
rect 7881 29731 7893 29765
rect 7927 29731 7939 29765
rect 7881 29697 7939 29731
rect 7881 29663 7893 29697
rect 7927 29663 7939 29697
rect 7881 29629 7939 29663
rect 7881 29595 7893 29629
rect 7927 29595 7939 29629
rect 7881 29561 7939 29595
rect 7881 29527 7893 29561
rect 7927 29527 7939 29561
rect 7881 29493 7939 29527
rect 7881 29459 7893 29493
rect 7927 29459 7939 29493
rect 7881 29425 7939 29459
rect 7881 29391 7893 29425
rect 7927 29391 7939 29425
rect 7881 29357 7939 29391
rect 7881 29323 7893 29357
rect 7927 29323 7939 29357
rect 7881 29289 7939 29323
rect 7881 29255 7893 29289
rect 7927 29255 7939 29289
rect 7881 29221 7939 29255
rect 7881 29187 7893 29221
rect 7927 29187 7939 29221
rect 7881 29153 7939 29187
rect 7881 29119 7893 29153
rect 7927 29119 7939 29153
rect 7881 29085 7939 29119
rect 7881 29051 7893 29085
rect 7927 29051 7939 29085
rect 7881 29017 7939 29051
rect 7881 28983 7893 29017
rect 7927 28983 7939 29017
rect 7881 28949 7939 28983
rect 7881 28915 7893 28949
rect 7927 28915 7939 28949
rect 7881 28881 7939 28915
rect 7881 28847 7893 28881
rect 7927 28847 7939 28881
rect 7881 28813 7939 28847
rect 7881 28779 7893 28813
rect 7927 28779 7939 28813
rect 7881 28745 7939 28779
rect 7881 28711 7893 28745
rect 7927 28711 7939 28745
rect 7881 28677 7939 28711
rect 7881 28643 7893 28677
rect 7927 28643 7939 28677
rect 7881 28627 7939 28643
rect 8339 29901 8397 29917
rect 8339 29867 8351 29901
rect 8385 29867 8397 29901
rect 8339 29833 8397 29867
rect 8339 29799 8351 29833
rect 8385 29799 8397 29833
rect 8339 29765 8397 29799
rect 8339 29731 8351 29765
rect 8385 29731 8397 29765
rect 8339 29697 8397 29731
rect 8339 29663 8351 29697
rect 8385 29663 8397 29697
rect 8339 29629 8397 29663
rect 8339 29595 8351 29629
rect 8385 29595 8397 29629
rect 8339 29561 8397 29595
rect 8339 29527 8351 29561
rect 8385 29527 8397 29561
rect 8339 29493 8397 29527
rect 8339 29459 8351 29493
rect 8385 29459 8397 29493
rect 8339 29425 8397 29459
rect 8339 29391 8351 29425
rect 8385 29391 8397 29425
rect 8339 29357 8397 29391
rect 8339 29323 8351 29357
rect 8385 29323 8397 29357
rect 8339 29289 8397 29323
rect 8339 29255 8351 29289
rect 8385 29255 8397 29289
rect 8339 29221 8397 29255
rect 8339 29187 8351 29221
rect 8385 29187 8397 29221
rect 8339 29153 8397 29187
rect 8339 29119 8351 29153
rect 8385 29119 8397 29153
rect 8339 29085 8397 29119
rect 8339 29051 8351 29085
rect 8385 29051 8397 29085
rect 8339 29017 8397 29051
rect 8339 28983 8351 29017
rect 8385 28983 8397 29017
rect 8339 28949 8397 28983
rect 8339 28915 8351 28949
rect 8385 28915 8397 28949
rect 8339 28881 8397 28915
rect 8339 28847 8351 28881
rect 8385 28847 8397 28881
rect 8339 28813 8397 28847
rect 8339 28779 8351 28813
rect 8385 28779 8397 28813
rect 8339 28745 8397 28779
rect 8339 28711 8351 28745
rect 8385 28711 8397 28745
rect 8339 28677 8397 28711
rect 8339 28643 8351 28677
rect 8385 28643 8397 28677
rect 8339 28627 8397 28643
rect 8797 29901 8855 29917
rect 8797 29867 8809 29901
rect 8843 29867 8855 29901
rect 8797 29833 8855 29867
rect 8797 29799 8809 29833
rect 8843 29799 8855 29833
rect 8797 29765 8855 29799
rect 8797 29731 8809 29765
rect 8843 29731 8855 29765
rect 8797 29697 8855 29731
rect 8797 29663 8809 29697
rect 8843 29663 8855 29697
rect 8797 29629 8855 29663
rect 8797 29595 8809 29629
rect 8843 29595 8855 29629
rect 8797 29561 8855 29595
rect 8797 29527 8809 29561
rect 8843 29527 8855 29561
rect 8797 29493 8855 29527
rect 8797 29459 8809 29493
rect 8843 29459 8855 29493
rect 8797 29425 8855 29459
rect 8797 29391 8809 29425
rect 8843 29391 8855 29425
rect 8797 29357 8855 29391
rect 8797 29323 8809 29357
rect 8843 29323 8855 29357
rect 8797 29289 8855 29323
rect 8797 29255 8809 29289
rect 8843 29255 8855 29289
rect 8797 29221 8855 29255
rect 8797 29187 8809 29221
rect 8843 29187 8855 29221
rect 8797 29153 8855 29187
rect 8797 29119 8809 29153
rect 8843 29119 8855 29153
rect 8797 29085 8855 29119
rect 8797 29051 8809 29085
rect 8843 29051 8855 29085
rect 8797 29017 8855 29051
rect 8797 28983 8809 29017
rect 8843 28983 8855 29017
rect 8797 28949 8855 28983
rect 8797 28915 8809 28949
rect 8843 28915 8855 28949
rect 8797 28881 8855 28915
rect 8797 28847 8809 28881
rect 8843 28847 8855 28881
rect 8797 28813 8855 28847
rect 8797 28779 8809 28813
rect 8843 28779 8855 28813
rect 8797 28745 8855 28779
rect 8797 28711 8809 28745
rect 8843 28711 8855 28745
rect 8797 28677 8855 28711
rect 8797 28643 8809 28677
rect 8843 28643 8855 28677
rect 8797 28627 8855 28643
rect 9255 29901 9313 29917
rect 9255 29867 9267 29901
rect 9301 29867 9313 29901
rect 9255 29833 9313 29867
rect 9255 29799 9267 29833
rect 9301 29799 9313 29833
rect 9255 29765 9313 29799
rect 9255 29731 9267 29765
rect 9301 29731 9313 29765
rect 9255 29697 9313 29731
rect 9255 29663 9267 29697
rect 9301 29663 9313 29697
rect 9255 29629 9313 29663
rect 9255 29595 9267 29629
rect 9301 29595 9313 29629
rect 9255 29561 9313 29595
rect 9255 29527 9267 29561
rect 9301 29527 9313 29561
rect 9255 29493 9313 29527
rect 9255 29459 9267 29493
rect 9301 29459 9313 29493
rect 9255 29425 9313 29459
rect 9255 29391 9267 29425
rect 9301 29391 9313 29425
rect 9255 29357 9313 29391
rect 9255 29323 9267 29357
rect 9301 29323 9313 29357
rect 9255 29289 9313 29323
rect 9255 29255 9267 29289
rect 9301 29255 9313 29289
rect 9255 29221 9313 29255
rect 9255 29187 9267 29221
rect 9301 29187 9313 29221
rect 9255 29153 9313 29187
rect 9255 29119 9267 29153
rect 9301 29119 9313 29153
rect 9255 29085 9313 29119
rect 9255 29051 9267 29085
rect 9301 29051 9313 29085
rect 9255 29017 9313 29051
rect 9255 28983 9267 29017
rect 9301 28983 9313 29017
rect 9255 28949 9313 28983
rect 9255 28915 9267 28949
rect 9301 28915 9313 28949
rect 9255 28881 9313 28915
rect 9255 28847 9267 28881
rect 9301 28847 9313 28881
rect 9255 28813 9313 28847
rect 9255 28779 9267 28813
rect 9301 28779 9313 28813
rect 9255 28745 9313 28779
rect 9255 28711 9267 28745
rect 9301 28711 9313 28745
rect 9255 28677 9313 28711
rect 9255 28643 9267 28677
rect 9301 28643 9313 28677
rect 9255 28627 9313 28643
rect 9713 29901 9771 29917
rect 9713 29867 9725 29901
rect 9759 29867 9771 29901
rect 9713 29833 9771 29867
rect 9713 29799 9725 29833
rect 9759 29799 9771 29833
rect 9713 29765 9771 29799
rect 9713 29731 9725 29765
rect 9759 29731 9771 29765
rect 9713 29697 9771 29731
rect 9713 29663 9725 29697
rect 9759 29663 9771 29697
rect 9713 29629 9771 29663
rect 9713 29595 9725 29629
rect 9759 29595 9771 29629
rect 9713 29561 9771 29595
rect 9713 29527 9725 29561
rect 9759 29527 9771 29561
rect 9713 29493 9771 29527
rect 9713 29459 9725 29493
rect 9759 29459 9771 29493
rect 9713 29425 9771 29459
rect 9713 29391 9725 29425
rect 9759 29391 9771 29425
rect 9713 29357 9771 29391
rect 9713 29323 9725 29357
rect 9759 29323 9771 29357
rect 9713 29289 9771 29323
rect 9713 29255 9725 29289
rect 9759 29255 9771 29289
rect 9713 29221 9771 29255
rect 9713 29187 9725 29221
rect 9759 29187 9771 29221
rect 9713 29153 9771 29187
rect 9713 29119 9725 29153
rect 9759 29119 9771 29153
rect 9713 29085 9771 29119
rect 9713 29051 9725 29085
rect 9759 29051 9771 29085
rect 9713 29017 9771 29051
rect 9713 28983 9725 29017
rect 9759 28983 9771 29017
rect 9713 28949 9771 28983
rect 9713 28915 9725 28949
rect 9759 28915 9771 28949
rect 9713 28881 9771 28915
rect 9713 28847 9725 28881
rect 9759 28847 9771 28881
rect 9713 28813 9771 28847
rect 9713 28779 9725 28813
rect 9759 28779 9771 28813
rect 9713 28745 9771 28779
rect 9713 28711 9725 28745
rect 9759 28711 9771 28745
rect 9713 28677 9771 28711
rect 9713 28643 9725 28677
rect 9759 28643 9771 28677
rect 9713 28627 9771 28643
rect 10171 29901 10229 29917
rect 10171 29867 10183 29901
rect 10217 29867 10229 29901
rect 10171 29833 10229 29867
rect 10171 29799 10183 29833
rect 10217 29799 10229 29833
rect 10171 29765 10229 29799
rect 10171 29731 10183 29765
rect 10217 29731 10229 29765
rect 10171 29697 10229 29731
rect 10171 29663 10183 29697
rect 10217 29663 10229 29697
rect 10171 29629 10229 29663
rect 10171 29595 10183 29629
rect 10217 29595 10229 29629
rect 10171 29561 10229 29595
rect 10171 29527 10183 29561
rect 10217 29527 10229 29561
rect 10171 29493 10229 29527
rect 10171 29459 10183 29493
rect 10217 29459 10229 29493
rect 10171 29425 10229 29459
rect 10171 29391 10183 29425
rect 10217 29391 10229 29425
rect 10171 29357 10229 29391
rect 10171 29323 10183 29357
rect 10217 29323 10229 29357
rect 10171 29289 10229 29323
rect 10171 29255 10183 29289
rect 10217 29255 10229 29289
rect 10171 29221 10229 29255
rect 10171 29187 10183 29221
rect 10217 29187 10229 29221
rect 10171 29153 10229 29187
rect 10171 29119 10183 29153
rect 10217 29119 10229 29153
rect 10171 29085 10229 29119
rect 10171 29051 10183 29085
rect 10217 29051 10229 29085
rect 10171 29017 10229 29051
rect 10171 28983 10183 29017
rect 10217 28983 10229 29017
rect 10171 28949 10229 28983
rect 10171 28915 10183 28949
rect 10217 28915 10229 28949
rect 10171 28881 10229 28915
rect 10171 28847 10183 28881
rect 10217 28847 10229 28881
rect 10171 28813 10229 28847
rect 10171 28779 10183 28813
rect 10217 28779 10229 28813
rect 10171 28745 10229 28779
rect 10171 28711 10183 28745
rect 10217 28711 10229 28745
rect 10171 28677 10229 28711
rect 10171 28643 10183 28677
rect 10217 28643 10229 28677
rect 10171 28627 10229 28643
rect 10629 29901 10687 29917
rect 10629 29867 10641 29901
rect 10675 29867 10687 29901
rect 10629 29833 10687 29867
rect 10629 29799 10641 29833
rect 10675 29799 10687 29833
rect 10629 29765 10687 29799
rect 10629 29731 10641 29765
rect 10675 29731 10687 29765
rect 10629 29697 10687 29731
rect 10629 29663 10641 29697
rect 10675 29663 10687 29697
rect 10629 29629 10687 29663
rect 10629 29595 10641 29629
rect 10675 29595 10687 29629
rect 10629 29561 10687 29595
rect 10629 29527 10641 29561
rect 10675 29527 10687 29561
rect 10629 29493 10687 29527
rect 10629 29459 10641 29493
rect 10675 29459 10687 29493
rect 10629 29425 10687 29459
rect 10629 29391 10641 29425
rect 10675 29391 10687 29425
rect 10629 29357 10687 29391
rect 10629 29323 10641 29357
rect 10675 29323 10687 29357
rect 10629 29289 10687 29323
rect 10629 29255 10641 29289
rect 10675 29255 10687 29289
rect 10629 29221 10687 29255
rect 10629 29187 10641 29221
rect 10675 29187 10687 29221
rect 10629 29153 10687 29187
rect 10629 29119 10641 29153
rect 10675 29119 10687 29153
rect 10629 29085 10687 29119
rect 10629 29051 10641 29085
rect 10675 29051 10687 29085
rect 10629 29017 10687 29051
rect 10629 28983 10641 29017
rect 10675 28983 10687 29017
rect 10629 28949 10687 28983
rect 10629 28915 10641 28949
rect 10675 28915 10687 28949
rect 10629 28881 10687 28915
rect 10629 28847 10641 28881
rect 10675 28847 10687 28881
rect 10629 28813 10687 28847
rect 10629 28779 10641 28813
rect 10675 28779 10687 28813
rect 10629 28745 10687 28779
rect 10629 28711 10641 28745
rect 10675 28711 10687 28745
rect 10629 28677 10687 28711
rect 10629 28643 10641 28677
rect 10675 28643 10687 28677
rect 10629 28627 10687 28643
rect 11087 29901 11145 29917
rect 11087 29867 11099 29901
rect 11133 29867 11145 29901
rect 11087 29833 11145 29867
rect 11087 29799 11099 29833
rect 11133 29799 11145 29833
rect 11087 29765 11145 29799
rect 11087 29731 11099 29765
rect 11133 29731 11145 29765
rect 11087 29697 11145 29731
rect 11087 29663 11099 29697
rect 11133 29663 11145 29697
rect 11087 29629 11145 29663
rect 11087 29595 11099 29629
rect 11133 29595 11145 29629
rect 11087 29561 11145 29595
rect 11087 29527 11099 29561
rect 11133 29527 11145 29561
rect 11087 29493 11145 29527
rect 11087 29459 11099 29493
rect 11133 29459 11145 29493
rect 11087 29425 11145 29459
rect 11087 29391 11099 29425
rect 11133 29391 11145 29425
rect 11087 29357 11145 29391
rect 11087 29323 11099 29357
rect 11133 29323 11145 29357
rect 11087 29289 11145 29323
rect 11087 29255 11099 29289
rect 11133 29255 11145 29289
rect 11087 29221 11145 29255
rect 11087 29187 11099 29221
rect 11133 29187 11145 29221
rect 11087 29153 11145 29187
rect 11087 29119 11099 29153
rect 11133 29119 11145 29153
rect 11087 29085 11145 29119
rect 11087 29051 11099 29085
rect 11133 29051 11145 29085
rect 11087 29017 11145 29051
rect 11087 28983 11099 29017
rect 11133 28983 11145 29017
rect 11087 28949 11145 28983
rect 11087 28915 11099 28949
rect 11133 28915 11145 28949
rect 11087 28881 11145 28915
rect 11087 28847 11099 28881
rect 11133 28847 11145 28881
rect 11087 28813 11145 28847
rect 11087 28779 11099 28813
rect 11133 28779 11145 28813
rect 11087 28745 11145 28779
rect 11087 28711 11099 28745
rect 11133 28711 11145 28745
rect 11087 28677 11145 28711
rect 11087 28643 11099 28677
rect 11133 28643 11145 28677
rect 11087 28627 11145 28643
rect 11545 29901 11603 29917
rect 11545 29867 11557 29901
rect 11591 29867 11603 29901
rect 11545 29833 11603 29867
rect 11545 29799 11557 29833
rect 11591 29799 11603 29833
rect 11545 29765 11603 29799
rect 11545 29731 11557 29765
rect 11591 29731 11603 29765
rect 11545 29697 11603 29731
rect 11545 29663 11557 29697
rect 11591 29663 11603 29697
rect 11545 29629 11603 29663
rect 11545 29595 11557 29629
rect 11591 29595 11603 29629
rect 11545 29561 11603 29595
rect 11545 29527 11557 29561
rect 11591 29527 11603 29561
rect 11545 29493 11603 29527
rect 11545 29459 11557 29493
rect 11591 29459 11603 29493
rect 11545 29425 11603 29459
rect 11545 29391 11557 29425
rect 11591 29391 11603 29425
rect 11545 29357 11603 29391
rect 11545 29323 11557 29357
rect 11591 29323 11603 29357
rect 11545 29289 11603 29323
rect 11545 29255 11557 29289
rect 11591 29255 11603 29289
rect 11545 29221 11603 29255
rect 11545 29187 11557 29221
rect 11591 29187 11603 29221
rect 11545 29153 11603 29187
rect 11545 29119 11557 29153
rect 11591 29119 11603 29153
rect 11545 29085 11603 29119
rect 11545 29051 11557 29085
rect 11591 29051 11603 29085
rect 11545 29017 11603 29051
rect 11545 28983 11557 29017
rect 11591 28983 11603 29017
rect 11545 28949 11603 28983
rect 11545 28915 11557 28949
rect 11591 28915 11603 28949
rect 11545 28881 11603 28915
rect 11545 28847 11557 28881
rect 11591 28847 11603 28881
rect 11545 28813 11603 28847
rect 11545 28779 11557 28813
rect 11591 28779 11603 28813
rect 11545 28745 11603 28779
rect 11545 28711 11557 28745
rect 11591 28711 11603 28745
rect 11545 28677 11603 28711
rect 11545 28643 11557 28677
rect 11591 28643 11603 28677
rect 11545 28627 11603 28643
rect 12003 29901 12061 29917
rect 12003 29867 12015 29901
rect 12049 29867 12061 29901
rect 12003 29833 12061 29867
rect 12003 29799 12015 29833
rect 12049 29799 12061 29833
rect 12003 29765 12061 29799
rect 12003 29731 12015 29765
rect 12049 29731 12061 29765
rect 12003 29697 12061 29731
rect 12003 29663 12015 29697
rect 12049 29663 12061 29697
rect 12003 29629 12061 29663
rect 12003 29595 12015 29629
rect 12049 29595 12061 29629
rect 12003 29561 12061 29595
rect 12003 29527 12015 29561
rect 12049 29527 12061 29561
rect 12003 29493 12061 29527
rect 12003 29459 12015 29493
rect 12049 29459 12061 29493
rect 12003 29425 12061 29459
rect 12003 29391 12015 29425
rect 12049 29391 12061 29425
rect 12003 29357 12061 29391
rect 12003 29323 12015 29357
rect 12049 29323 12061 29357
rect 12003 29289 12061 29323
rect 12003 29255 12015 29289
rect 12049 29255 12061 29289
rect 12003 29221 12061 29255
rect 12003 29187 12015 29221
rect 12049 29187 12061 29221
rect 12003 29153 12061 29187
rect 12003 29119 12015 29153
rect 12049 29119 12061 29153
rect 12003 29085 12061 29119
rect 12003 29051 12015 29085
rect 12049 29051 12061 29085
rect 12003 29017 12061 29051
rect 12003 28983 12015 29017
rect 12049 28983 12061 29017
rect 12003 28949 12061 28983
rect 12003 28915 12015 28949
rect 12049 28915 12061 28949
rect 12003 28881 12061 28915
rect 12003 28847 12015 28881
rect 12049 28847 12061 28881
rect 12003 28813 12061 28847
rect 12003 28779 12015 28813
rect 12049 28779 12061 28813
rect 12003 28745 12061 28779
rect 12003 28711 12015 28745
rect 12049 28711 12061 28745
rect 12003 28677 12061 28711
rect 12003 28643 12015 28677
rect 12049 28643 12061 28677
rect 12003 28627 12061 28643
rect 12461 29901 12519 29917
rect 12461 29867 12473 29901
rect 12507 29867 12519 29901
rect 12461 29833 12519 29867
rect 12461 29799 12473 29833
rect 12507 29799 12519 29833
rect 12461 29765 12519 29799
rect 12461 29731 12473 29765
rect 12507 29731 12519 29765
rect 12461 29697 12519 29731
rect 12461 29663 12473 29697
rect 12507 29663 12519 29697
rect 12461 29629 12519 29663
rect 12461 29595 12473 29629
rect 12507 29595 12519 29629
rect 12461 29561 12519 29595
rect 12461 29527 12473 29561
rect 12507 29527 12519 29561
rect 12461 29493 12519 29527
rect 12461 29459 12473 29493
rect 12507 29459 12519 29493
rect 12461 29425 12519 29459
rect 12461 29391 12473 29425
rect 12507 29391 12519 29425
rect 12461 29357 12519 29391
rect 12461 29323 12473 29357
rect 12507 29323 12519 29357
rect 12461 29289 12519 29323
rect 12461 29255 12473 29289
rect 12507 29255 12519 29289
rect 12461 29221 12519 29255
rect 12461 29187 12473 29221
rect 12507 29187 12519 29221
rect 12461 29153 12519 29187
rect 12461 29119 12473 29153
rect 12507 29119 12519 29153
rect 12461 29085 12519 29119
rect 12461 29051 12473 29085
rect 12507 29051 12519 29085
rect 12461 29017 12519 29051
rect 12461 28983 12473 29017
rect 12507 28983 12519 29017
rect 12461 28949 12519 28983
rect 12461 28915 12473 28949
rect 12507 28915 12519 28949
rect 12461 28881 12519 28915
rect 12461 28847 12473 28881
rect 12507 28847 12519 28881
rect 12461 28813 12519 28847
rect 12461 28779 12473 28813
rect 12507 28779 12519 28813
rect 12461 28745 12519 28779
rect 12461 28711 12473 28745
rect 12507 28711 12519 28745
rect 12461 28677 12519 28711
rect 12461 28643 12473 28677
rect 12507 28643 12519 28677
rect 12461 28627 12519 28643
rect 12919 29901 12977 29917
rect 12919 29867 12931 29901
rect 12965 29867 12977 29901
rect 12919 29833 12977 29867
rect 12919 29799 12931 29833
rect 12965 29799 12977 29833
rect 12919 29765 12977 29799
rect 12919 29731 12931 29765
rect 12965 29731 12977 29765
rect 12919 29697 12977 29731
rect 12919 29663 12931 29697
rect 12965 29663 12977 29697
rect 12919 29629 12977 29663
rect 12919 29595 12931 29629
rect 12965 29595 12977 29629
rect 12919 29561 12977 29595
rect 12919 29527 12931 29561
rect 12965 29527 12977 29561
rect 12919 29493 12977 29527
rect 12919 29459 12931 29493
rect 12965 29459 12977 29493
rect 12919 29425 12977 29459
rect 12919 29391 12931 29425
rect 12965 29391 12977 29425
rect 12919 29357 12977 29391
rect 12919 29323 12931 29357
rect 12965 29323 12977 29357
rect 12919 29289 12977 29323
rect 12919 29255 12931 29289
rect 12965 29255 12977 29289
rect 12919 29221 12977 29255
rect 12919 29187 12931 29221
rect 12965 29187 12977 29221
rect 12919 29153 12977 29187
rect 12919 29119 12931 29153
rect 12965 29119 12977 29153
rect 12919 29085 12977 29119
rect 12919 29051 12931 29085
rect 12965 29051 12977 29085
rect 12919 29017 12977 29051
rect 12919 28983 12931 29017
rect 12965 28983 12977 29017
rect 12919 28949 12977 28983
rect 12919 28915 12931 28949
rect 12965 28915 12977 28949
rect 12919 28881 12977 28915
rect 12919 28847 12931 28881
rect 12965 28847 12977 28881
rect 12919 28813 12977 28847
rect 12919 28779 12931 28813
rect 12965 28779 12977 28813
rect 12919 28745 12977 28779
rect 12919 28711 12931 28745
rect 12965 28711 12977 28745
rect 12919 28677 12977 28711
rect 12919 28643 12931 28677
rect 12965 28643 12977 28677
rect 12919 28627 12977 28643
rect 13377 29901 13435 29917
rect 13377 29867 13389 29901
rect 13423 29867 13435 29901
rect 13377 29833 13435 29867
rect 13377 29799 13389 29833
rect 13423 29799 13435 29833
rect 13377 29765 13435 29799
rect 13377 29731 13389 29765
rect 13423 29731 13435 29765
rect 13377 29697 13435 29731
rect 13377 29663 13389 29697
rect 13423 29663 13435 29697
rect 13377 29629 13435 29663
rect 13377 29595 13389 29629
rect 13423 29595 13435 29629
rect 13377 29561 13435 29595
rect 13377 29527 13389 29561
rect 13423 29527 13435 29561
rect 13377 29493 13435 29527
rect 13377 29459 13389 29493
rect 13423 29459 13435 29493
rect 13377 29425 13435 29459
rect 13377 29391 13389 29425
rect 13423 29391 13435 29425
rect 13377 29357 13435 29391
rect 13377 29323 13389 29357
rect 13423 29323 13435 29357
rect 13377 29289 13435 29323
rect 13377 29255 13389 29289
rect 13423 29255 13435 29289
rect 13377 29221 13435 29255
rect 13377 29187 13389 29221
rect 13423 29187 13435 29221
rect 13377 29153 13435 29187
rect 13377 29119 13389 29153
rect 13423 29119 13435 29153
rect 13377 29085 13435 29119
rect 13377 29051 13389 29085
rect 13423 29051 13435 29085
rect 13377 29017 13435 29051
rect 13377 28983 13389 29017
rect 13423 28983 13435 29017
rect 13377 28949 13435 28983
rect 13377 28915 13389 28949
rect 13423 28915 13435 28949
rect 13377 28881 13435 28915
rect 13377 28847 13389 28881
rect 13423 28847 13435 28881
rect 13377 28813 13435 28847
rect 13377 28779 13389 28813
rect 13423 28779 13435 28813
rect 13377 28745 13435 28779
rect 13377 28711 13389 28745
rect 13423 28711 13435 28745
rect 13377 28677 13435 28711
rect 13377 28643 13389 28677
rect 13423 28643 13435 28677
rect 13377 28627 13435 28643
rect 13835 29901 13893 29917
rect 13835 29867 13847 29901
rect 13881 29867 13893 29901
rect 13835 29833 13893 29867
rect 13835 29799 13847 29833
rect 13881 29799 13893 29833
rect 13835 29765 13893 29799
rect 13835 29731 13847 29765
rect 13881 29731 13893 29765
rect 13835 29697 13893 29731
rect 13835 29663 13847 29697
rect 13881 29663 13893 29697
rect 13835 29629 13893 29663
rect 13835 29595 13847 29629
rect 13881 29595 13893 29629
rect 13835 29561 13893 29595
rect 13835 29527 13847 29561
rect 13881 29527 13893 29561
rect 13835 29493 13893 29527
rect 13835 29459 13847 29493
rect 13881 29459 13893 29493
rect 13835 29425 13893 29459
rect 13835 29391 13847 29425
rect 13881 29391 13893 29425
rect 13835 29357 13893 29391
rect 13835 29323 13847 29357
rect 13881 29323 13893 29357
rect 13835 29289 13893 29323
rect 13835 29255 13847 29289
rect 13881 29255 13893 29289
rect 13835 29221 13893 29255
rect 13835 29187 13847 29221
rect 13881 29187 13893 29221
rect 13835 29153 13893 29187
rect 13835 29119 13847 29153
rect 13881 29119 13893 29153
rect 13835 29085 13893 29119
rect 13835 29051 13847 29085
rect 13881 29051 13893 29085
rect 13835 29017 13893 29051
rect 13835 28983 13847 29017
rect 13881 28983 13893 29017
rect 13835 28949 13893 28983
rect 13835 28915 13847 28949
rect 13881 28915 13893 28949
rect 13835 28881 13893 28915
rect 13835 28847 13847 28881
rect 13881 28847 13893 28881
rect 13835 28813 13893 28847
rect 13835 28779 13847 28813
rect 13881 28779 13893 28813
rect 13835 28745 13893 28779
rect 13835 28711 13847 28745
rect 13881 28711 13893 28745
rect 13835 28677 13893 28711
rect 13835 28643 13847 28677
rect 13881 28643 13893 28677
rect 13835 28627 13893 28643
rect 14293 29901 14351 29917
rect 14293 29867 14305 29901
rect 14339 29867 14351 29901
rect 14293 29833 14351 29867
rect 14293 29799 14305 29833
rect 14339 29799 14351 29833
rect 14293 29765 14351 29799
rect 14293 29731 14305 29765
rect 14339 29731 14351 29765
rect 14293 29697 14351 29731
rect 14293 29663 14305 29697
rect 14339 29663 14351 29697
rect 14293 29629 14351 29663
rect 14293 29595 14305 29629
rect 14339 29595 14351 29629
rect 14293 29561 14351 29595
rect 14293 29527 14305 29561
rect 14339 29527 14351 29561
rect 14293 29493 14351 29527
rect 14293 29459 14305 29493
rect 14339 29459 14351 29493
rect 14293 29425 14351 29459
rect 14293 29391 14305 29425
rect 14339 29391 14351 29425
rect 14293 29357 14351 29391
rect 14293 29323 14305 29357
rect 14339 29323 14351 29357
rect 14293 29289 14351 29323
rect 14293 29255 14305 29289
rect 14339 29255 14351 29289
rect 14293 29221 14351 29255
rect 14293 29187 14305 29221
rect 14339 29187 14351 29221
rect 14293 29153 14351 29187
rect 14293 29119 14305 29153
rect 14339 29119 14351 29153
rect 14293 29085 14351 29119
rect 14293 29051 14305 29085
rect 14339 29051 14351 29085
rect 14293 29017 14351 29051
rect 14293 28983 14305 29017
rect 14339 28983 14351 29017
rect 14293 28949 14351 28983
rect 14293 28915 14305 28949
rect 14339 28915 14351 28949
rect 14293 28881 14351 28915
rect 14293 28847 14305 28881
rect 14339 28847 14351 28881
rect 14293 28813 14351 28847
rect 14293 28779 14305 28813
rect 14339 28779 14351 28813
rect 14293 28745 14351 28779
rect 14293 28711 14305 28745
rect 14339 28711 14351 28745
rect 14293 28677 14351 28711
rect 14293 28643 14305 28677
rect 14339 28643 14351 28677
rect 14293 28627 14351 28643
rect 14751 29901 14809 29917
rect 14751 29867 14763 29901
rect 14797 29867 14809 29901
rect 14751 29833 14809 29867
rect 14751 29799 14763 29833
rect 14797 29799 14809 29833
rect 14751 29765 14809 29799
rect 14751 29731 14763 29765
rect 14797 29731 14809 29765
rect 14751 29697 14809 29731
rect 14751 29663 14763 29697
rect 14797 29663 14809 29697
rect 14751 29629 14809 29663
rect 14751 29595 14763 29629
rect 14797 29595 14809 29629
rect 14751 29561 14809 29595
rect 14751 29527 14763 29561
rect 14797 29527 14809 29561
rect 14751 29493 14809 29527
rect 14751 29459 14763 29493
rect 14797 29459 14809 29493
rect 14751 29425 14809 29459
rect 14751 29391 14763 29425
rect 14797 29391 14809 29425
rect 14751 29357 14809 29391
rect 14751 29323 14763 29357
rect 14797 29323 14809 29357
rect 14751 29289 14809 29323
rect 14751 29255 14763 29289
rect 14797 29255 14809 29289
rect 14751 29221 14809 29255
rect 14751 29187 14763 29221
rect 14797 29187 14809 29221
rect 14751 29153 14809 29187
rect 14751 29119 14763 29153
rect 14797 29119 14809 29153
rect 14751 29085 14809 29119
rect 14751 29051 14763 29085
rect 14797 29051 14809 29085
rect 14751 29017 14809 29051
rect 14751 28983 14763 29017
rect 14797 28983 14809 29017
rect 14751 28949 14809 28983
rect 14751 28915 14763 28949
rect 14797 28915 14809 28949
rect 14751 28881 14809 28915
rect 14751 28847 14763 28881
rect 14797 28847 14809 28881
rect 14751 28813 14809 28847
rect 14751 28779 14763 28813
rect 14797 28779 14809 28813
rect 14751 28745 14809 28779
rect 14751 28711 14763 28745
rect 14797 28711 14809 28745
rect 14751 28677 14809 28711
rect 14751 28643 14763 28677
rect 14797 28643 14809 28677
rect 14751 28627 14809 28643
rect 15209 29901 15267 29917
rect 15209 29867 15221 29901
rect 15255 29867 15267 29901
rect 15209 29833 15267 29867
rect 15209 29799 15221 29833
rect 15255 29799 15267 29833
rect 15209 29765 15267 29799
rect 15209 29731 15221 29765
rect 15255 29731 15267 29765
rect 15209 29697 15267 29731
rect 15209 29663 15221 29697
rect 15255 29663 15267 29697
rect 15209 29629 15267 29663
rect 15209 29595 15221 29629
rect 15255 29595 15267 29629
rect 15209 29561 15267 29595
rect 15209 29527 15221 29561
rect 15255 29527 15267 29561
rect 15209 29493 15267 29527
rect 15209 29459 15221 29493
rect 15255 29459 15267 29493
rect 15209 29425 15267 29459
rect 15209 29391 15221 29425
rect 15255 29391 15267 29425
rect 15209 29357 15267 29391
rect 15209 29323 15221 29357
rect 15255 29323 15267 29357
rect 15209 29289 15267 29323
rect 15209 29255 15221 29289
rect 15255 29255 15267 29289
rect 15209 29221 15267 29255
rect 15209 29187 15221 29221
rect 15255 29187 15267 29221
rect 15209 29153 15267 29187
rect 15209 29119 15221 29153
rect 15255 29119 15267 29153
rect 15209 29085 15267 29119
rect 15209 29051 15221 29085
rect 15255 29051 15267 29085
rect 15209 29017 15267 29051
rect 15209 28983 15221 29017
rect 15255 28983 15267 29017
rect 15209 28949 15267 28983
rect 15209 28915 15221 28949
rect 15255 28915 15267 28949
rect 15209 28881 15267 28915
rect 15209 28847 15221 28881
rect 15255 28847 15267 28881
rect 15209 28813 15267 28847
rect 15209 28779 15221 28813
rect 15255 28779 15267 28813
rect 15209 28745 15267 28779
rect 15209 28711 15221 28745
rect 15255 28711 15267 28745
rect 15209 28677 15267 28711
rect 15209 28643 15221 28677
rect 15255 28643 15267 28677
rect 15209 28627 15267 28643
rect 15667 29901 15725 29917
rect 15667 29867 15679 29901
rect 15713 29867 15725 29901
rect 15667 29833 15725 29867
rect 15667 29799 15679 29833
rect 15713 29799 15725 29833
rect 15667 29765 15725 29799
rect 15667 29731 15679 29765
rect 15713 29731 15725 29765
rect 15667 29697 15725 29731
rect 15667 29663 15679 29697
rect 15713 29663 15725 29697
rect 15667 29629 15725 29663
rect 15667 29595 15679 29629
rect 15713 29595 15725 29629
rect 15667 29561 15725 29595
rect 15667 29527 15679 29561
rect 15713 29527 15725 29561
rect 15667 29493 15725 29527
rect 15667 29459 15679 29493
rect 15713 29459 15725 29493
rect 15667 29425 15725 29459
rect 15667 29391 15679 29425
rect 15713 29391 15725 29425
rect 15667 29357 15725 29391
rect 15667 29323 15679 29357
rect 15713 29323 15725 29357
rect 15667 29289 15725 29323
rect 15667 29255 15679 29289
rect 15713 29255 15725 29289
rect 15667 29221 15725 29255
rect 15667 29187 15679 29221
rect 15713 29187 15725 29221
rect 15667 29153 15725 29187
rect 15667 29119 15679 29153
rect 15713 29119 15725 29153
rect 15667 29085 15725 29119
rect 15667 29051 15679 29085
rect 15713 29051 15725 29085
rect 15667 29017 15725 29051
rect 15667 28983 15679 29017
rect 15713 28983 15725 29017
rect 15667 28949 15725 28983
rect 15667 28915 15679 28949
rect 15713 28915 15725 28949
rect 15667 28881 15725 28915
rect 15667 28847 15679 28881
rect 15713 28847 15725 28881
rect 15667 28813 15725 28847
rect 15667 28779 15679 28813
rect 15713 28779 15725 28813
rect 15667 28745 15725 28779
rect 15667 28711 15679 28745
rect 15713 28711 15725 28745
rect 15667 28677 15725 28711
rect 15667 28643 15679 28677
rect 15713 28643 15725 28677
rect 15667 28627 15725 28643
rect 16125 29901 16183 29917
rect 16125 29867 16137 29901
rect 16171 29867 16183 29901
rect 16125 29833 16183 29867
rect 16125 29799 16137 29833
rect 16171 29799 16183 29833
rect 16125 29765 16183 29799
rect 16125 29731 16137 29765
rect 16171 29731 16183 29765
rect 16125 29697 16183 29731
rect 16125 29663 16137 29697
rect 16171 29663 16183 29697
rect 16125 29629 16183 29663
rect 16125 29595 16137 29629
rect 16171 29595 16183 29629
rect 16125 29561 16183 29595
rect 16125 29527 16137 29561
rect 16171 29527 16183 29561
rect 16125 29493 16183 29527
rect 16125 29459 16137 29493
rect 16171 29459 16183 29493
rect 16125 29425 16183 29459
rect 16125 29391 16137 29425
rect 16171 29391 16183 29425
rect 16125 29357 16183 29391
rect 16125 29323 16137 29357
rect 16171 29323 16183 29357
rect 16125 29289 16183 29323
rect 16125 29255 16137 29289
rect 16171 29255 16183 29289
rect 16125 29221 16183 29255
rect 16125 29187 16137 29221
rect 16171 29187 16183 29221
rect 16125 29153 16183 29187
rect 16125 29119 16137 29153
rect 16171 29119 16183 29153
rect 16125 29085 16183 29119
rect 16125 29051 16137 29085
rect 16171 29051 16183 29085
rect 16125 29017 16183 29051
rect 16125 28983 16137 29017
rect 16171 28983 16183 29017
rect 16125 28949 16183 28983
rect 16125 28915 16137 28949
rect 16171 28915 16183 28949
rect 16125 28881 16183 28915
rect 16125 28847 16137 28881
rect 16171 28847 16183 28881
rect 16125 28813 16183 28847
rect 16125 28779 16137 28813
rect 16171 28779 16183 28813
rect 16125 28745 16183 28779
rect 16125 28711 16137 28745
rect 16171 28711 16183 28745
rect 16125 28677 16183 28711
rect 16125 28643 16137 28677
rect 16171 28643 16183 28677
rect 16125 28627 16183 28643
rect 16583 29901 16641 29917
rect 16583 29867 16595 29901
rect 16629 29867 16641 29901
rect 16583 29833 16641 29867
rect 16583 29799 16595 29833
rect 16629 29799 16641 29833
rect 16583 29765 16641 29799
rect 16583 29731 16595 29765
rect 16629 29731 16641 29765
rect 16583 29697 16641 29731
rect 16583 29663 16595 29697
rect 16629 29663 16641 29697
rect 16583 29629 16641 29663
rect 16583 29595 16595 29629
rect 16629 29595 16641 29629
rect 16583 29561 16641 29595
rect 16583 29527 16595 29561
rect 16629 29527 16641 29561
rect 16583 29493 16641 29527
rect 16583 29459 16595 29493
rect 16629 29459 16641 29493
rect 16583 29425 16641 29459
rect 16583 29391 16595 29425
rect 16629 29391 16641 29425
rect 16583 29357 16641 29391
rect 16583 29323 16595 29357
rect 16629 29323 16641 29357
rect 16583 29289 16641 29323
rect 16583 29255 16595 29289
rect 16629 29255 16641 29289
rect 16583 29221 16641 29255
rect 16583 29187 16595 29221
rect 16629 29187 16641 29221
rect 16583 29153 16641 29187
rect 16583 29119 16595 29153
rect 16629 29119 16641 29153
rect 16583 29085 16641 29119
rect 16583 29051 16595 29085
rect 16629 29051 16641 29085
rect 16583 29017 16641 29051
rect 16583 28983 16595 29017
rect 16629 28983 16641 29017
rect 16583 28949 16641 28983
rect 16583 28915 16595 28949
rect 16629 28915 16641 28949
rect 16583 28881 16641 28915
rect 16583 28847 16595 28881
rect 16629 28847 16641 28881
rect 16583 28813 16641 28847
rect 16583 28779 16595 28813
rect 16629 28779 16641 28813
rect 16583 28745 16641 28779
rect 16583 28711 16595 28745
rect 16629 28711 16641 28745
rect 16583 28677 16641 28711
rect 16583 28643 16595 28677
rect 16629 28643 16641 28677
rect 16583 28627 16641 28643
rect 17041 29901 17099 29917
rect 17041 29867 17053 29901
rect 17087 29867 17099 29901
rect 17041 29833 17099 29867
rect 17041 29799 17053 29833
rect 17087 29799 17099 29833
rect 17041 29765 17099 29799
rect 17041 29731 17053 29765
rect 17087 29731 17099 29765
rect 17041 29697 17099 29731
rect 17041 29663 17053 29697
rect 17087 29663 17099 29697
rect 17041 29629 17099 29663
rect 17041 29595 17053 29629
rect 17087 29595 17099 29629
rect 17041 29561 17099 29595
rect 17041 29527 17053 29561
rect 17087 29527 17099 29561
rect 17041 29493 17099 29527
rect 17041 29459 17053 29493
rect 17087 29459 17099 29493
rect 17041 29425 17099 29459
rect 17041 29391 17053 29425
rect 17087 29391 17099 29425
rect 17041 29357 17099 29391
rect 17041 29323 17053 29357
rect 17087 29323 17099 29357
rect 17041 29289 17099 29323
rect 17041 29255 17053 29289
rect 17087 29255 17099 29289
rect 17041 29221 17099 29255
rect 17041 29187 17053 29221
rect 17087 29187 17099 29221
rect 17041 29153 17099 29187
rect 17041 29119 17053 29153
rect 17087 29119 17099 29153
rect 17041 29085 17099 29119
rect 17041 29051 17053 29085
rect 17087 29051 17099 29085
rect 17041 29017 17099 29051
rect 17041 28983 17053 29017
rect 17087 28983 17099 29017
rect 17041 28949 17099 28983
rect 17041 28915 17053 28949
rect 17087 28915 17099 28949
rect 17041 28881 17099 28915
rect 17041 28847 17053 28881
rect 17087 28847 17099 28881
rect 17041 28813 17099 28847
rect 17041 28779 17053 28813
rect 17087 28779 17099 28813
rect 17041 28745 17099 28779
rect 17041 28711 17053 28745
rect 17087 28711 17099 28745
rect 17041 28677 17099 28711
rect 17041 28643 17053 28677
rect 17087 28643 17099 28677
rect 17041 28627 17099 28643
rect 17499 29901 17557 29917
rect 17499 29867 17511 29901
rect 17545 29867 17557 29901
rect 17499 29833 17557 29867
rect 17499 29799 17511 29833
rect 17545 29799 17557 29833
rect 17499 29765 17557 29799
rect 17499 29731 17511 29765
rect 17545 29731 17557 29765
rect 17499 29697 17557 29731
rect 17499 29663 17511 29697
rect 17545 29663 17557 29697
rect 17499 29629 17557 29663
rect 17499 29595 17511 29629
rect 17545 29595 17557 29629
rect 17499 29561 17557 29595
rect 17499 29527 17511 29561
rect 17545 29527 17557 29561
rect 17499 29493 17557 29527
rect 17499 29459 17511 29493
rect 17545 29459 17557 29493
rect 17499 29425 17557 29459
rect 17499 29391 17511 29425
rect 17545 29391 17557 29425
rect 17499 29357 17557 29391
rect 17499 29323 17511 29357
rect 17545 29323 17557 29357
rect 17499 29289 17557 29323
rect 17499 29255 17511 29289
rect 17545 29255 17557 29289
rect 17499 29221 17557 29255
rect 17499 29187 17511 29221
rect 17545 29187 17557 29221
rect 17499 29153 17557 29187
rect 17499 29119 17511 29153
rect 17545 29119 17557 29153
rect 17499 29085 17557 29119
rect 17499 29051 17511 29085
rect 17545 29051 17557 29085
rect 17499 29017 17557 29051
rect 17499 28983 17511 29017
rect 17545 28983 17557 29017
rect 17499 28949 17557 28983
rect 17499 28915 17511 28949
rect 17545 28915 17557 28949
rect 17499 28881 17557 28915
rect 17499 28847 17511 28881
rect 17545 28847 17557 28881
rect 17499 28813 17557 28847
rect 17499 28779 17511 28813
rect 17545 28779 17557 28813
rect 17499 28745 17557 28779
rect 17499 28711 17511 28745
rect 17545 28711 17557 28745
rect 17499 28677 17557 28711
rect 17499 28643 17511 28677
rect 17545 28643 17557 28677
rect 17499 28627 17557 28643
rect 17957 29901 18015 29917
rect 17957 29867 17969 29901
rect 18003 29867 18015 29901
rect 17957 29833 18015 29867
rect 17957 29799 17969 29833
rect 18003 29799 18015 29833
rect 17957 29765 18015 29799
rect 17957 29731 17969 29765
rect 18003 29731 18015 29765
rect 17957 29697 18015 29731
rect 17957 29663 17969 29697
rect 18003 29663 18015 29697
rect 17957 29629 18015 29663
rect 17957 29595 17969 29629
rect 18003 29595 18015 29629
rect 17957 29561 18015 29595
rect 17957 29527 17969 29561
rect 18003 29527 18015 29561
rect 17957 29493 18015 29527
rect 17957 29459 17969 29493
rect 18003 29459 18015 29493
rect 17957 29425 18015 29459
rect 17957 29391 17969 29425
rect 18003 29391 18015 29425
rect 17957 29357 18015 29391
rect 17957 29323 17969 29357
rect 18003 29323 18015 29357
rect 17957 29289 18015 29323
rect 17957 29255 17969 29289
rect 18003 29255 18015 29289
rect 17957 29221 18015 29255
rect 17957 29187 17969 29221
rect 18003 29187 18015 29221
rect 17957 29153 18015 29187
rect 17957 29119 17969 29153
rect 18003 29119 18015 29153
rect 17957 29085 18015 29119
rect 17957 29051 17969 29085
rect 18003 29051 18015 29085
rect 17957 29017 18015 29051
rect 17957 28983 17969 29017
rect 18003 28983 18015 29017
rect 17957 28949 18015 28983
rect 17957 28915 17969 28949
rect 18003 28915 18015 28949
rect 17957 28881 18015 28915
rect 17957 28847 17969 28881
rect 18003 28847 18015 28881
rect 17957 28813 18015 28847
rect 17957 28779 17969 28813
rect 18003 28779 18015 28813
rect 17957 28745 18015 28779
rect 17957 28711 17969 28745
rect 18003 28711 18015 28745
rect 17957 28677 18015 28711
rect 17957 28643 17969 28677
rect 18003 28643 18015 28677
rect 17957 28627 18015 28643
rect 18415 29901 18473 29917
rect 18415 29867 18427 29901
rect 18461 29867 18473 29901
rect 18415 29833 18473 29867
rect 18415 29799 18427 29833
rect 18461 29799 18473 29833
rect 18415 29765 18473 29799
rect 18415 29731 18427 29765
rect 18461 29731 18473 29765
rect 18415 29697 18473 29731
rect 18415 29663 18427 29697
rect 18461 29663 18473 29697
rect 18415 29629 18473 29663
rect 18415 29595 18427 29629
rect 18461 29595 18473 29629
rect 18415 29561 18473 29595
rect 18415 29527 18427 29561
rect 18461 29527 18473 29561
rect 18415 29493 18473 29527
rect 18415 29459 18427 29493
rect 18461 29459 18473 29493
rect 18415 29425 18473 29459
rect 18415 29391 18427 29425
rect 18461 29391 18473 29425
rect 18415 29357 18473 29391
rect 18415 29323 18427 29357
rect 18461 29323 18473 29357
rect 18415 29289 18473 29323
rect 18415 29255 18427 29289
rect 18461 29255 18473 29289
rect 18415 29221 18473 29255
rect 18415 29187 18427 29221
rect 18461 29187 18473 29221
rect 18415 29153 18473 29187
rect 18415 29119 18427 29153
rect 18461 29119 18473 29153
rect 18415 29085 18473 29119
rect 18415 29051 18427 29085
rect 18461 29051 18473 29085
rect 18415 29017 18473 29051
rect 18415 28983 18427 29017
rect 18461 28983 18473 29017
rect 18415 28949 18473 28983
rect 18415 28915 18427 28949
rect 18461 28915 18473 28949
rect 18415 28881 18473 28915
rect 18415 28847 18427 28881
rect 18461 28847 18473 28881
rect 18415 28813 18473 28847
rect 18415 28779 18427 28813
rect 18461 28779 18473 28813
rect 18415 28745 18473 28779
rect 18415 28711 18427 28745
rect 18461 28711 18473 28745
rect 18415 28677 18473 28711
rect 18415 28643 18427 28677
rect 18461 28643 18473 28677
rect 18415 28627 18473 28643
rect 18873 29901 18931 29917
rect 18873 29867 18885 29901
rect 18919 29867 18931 29901
rect 18873 29833 18931 29867
rect 18873 29799 18885 29833
rect 18919 29799 18931 29833
rect 18873 29765 18931 29799
rect 18873 29731 18885 29765
rect 18919 29731 18931 29765
rect 18873 29697 18931 29731
rect 18873 29663 18885 29697
rect 18919 29663 18931 29697
rect 18873 29629 18931 29663
rect 18873 29595 18885 29629
rect 18919 29595 18931 29629
rect 18873 29561 18931 29595
rect 18873 29527 18885 29561
rect 18919 29527 18931 29561
rect 18873 29493 18931 29527
rect 18873 29459 18885 29493
rect 18919 29459 18931 29493
rect 18873 29425 18931 29459
rect 18873 29391 18885 29425
rect 18919 29391 18931 29425
rect 18873 29357 18931 29391
rect 18873 29323 18885 29357
rect 18919 29323 18931 29357
rect 18873 29289 18931 29323
rect 18873 29255 18885 29289
rect 18919 29255 18931 29289
rect 18873 29221 18931 29255
rect 18873 29187 18885 29221
rect 18919 29187 18931 29221
rect 18873 29153 18931 29187
rect 18873 29119 18885 29153
rect 18919 29119 18931 29153
rect 18873 29085 18931 29119
rect 18873 29051 18885 29085
rect 18919 29051 18931 29085
rect 18873 29017 18931 29051
rect 18873 28983 18885 29017
rect 18919 28983 18931 29017
rect 18873 28949 18931 28983
rect 18873 28915 18885 28949
rect 18919 28915 18931 28949
rect 18873 28881 18931 28915
rect 18873 28847 18885 28881
rect 18919 28847 18931 28881
rect 18873 28813 18931 28847
rect 18873 28779 18885 28813
rect 18919 28779 18931 28813
rect 18873 28745 18931 28779
rect 18873 28711 18885 28745
rect 18919 28711 18931 28745
rect 18873 28677 18931 28711
rect 18873 28643 18885 28677
rect 18919 28643 18931 28677
rect 18873 28627 18931 28643
rect 19331 29901 19389 29917
rect 19331 29867 19343 29901
rect 19377 29867 19389 29901
rect 19331 29833 19389 29867
rect 19331 29799 19343 29833
rect 19377 29799 19389 29833
rect 19331 29765 19389 29799
rect 19331 29731 19343 29765
rect 19377 29731 19389 29765
rect 19331 29697 19389 29731
rect 19331 29663 19343 29697
rect 19377 29663 19389 29697
rect 19331 29629 19389 29663
rect 19331 29595 19343 29629
rect 19377 29595 19389 29629
rect 19331 29561 19389 29595
rect 19331 29527 19343 29561
rect 19377 29527 19389 29561
rect 19331 29493 19389 29527
rect 19331 29459 19343 29493
rect 19377 29459 19389 29493
rect 19331 29425 19389 29459
rect 19331 29391 19343 29425
rect 19377 29391 19389 29425
rect 19331 29357 19389 29391
rect 19331 29323 19343 29357
rect 19377 29323 19389 29357
rect 19331 29289 19389 29323
rect 19331 29255 19343 29289
rect 19377 29255 19389 29289
rect 19331 29221 19389 29255
rect 19331 29187 19343 29221
rect 19377 29187 19389 29221
rect 19331 29153 19389 29187
rect 19331 29119 19343 29153
rect 19377 29119 19389 29153
rect 19331 29085 19389 29119
rect 19331 29051 19343 29085
rect 19377 29051 19389 29085
rect 19331 29017 19389 29051
rect 19331 28983 19343 29017
rect 19377 28983 19389 29017
rect 19331 28949 19389 28983
rect 19331 28915 19343 28949
rect 19377 28915 19389 28949
rect 19331 28881 19389 28915
rect 19331 28847 19343 28881
rect 19377 28847 19389 28881
rect 19331 28813 19389 28847
rect 19331 28779 19343 28813
rect 19377 28779 19389 28813
rect 19331 28745 19389 28779
rect 19331 28711 19343 28745
rect 19377 28711 19389 28745
rect 19331 28677 19389 28711
rect 19331 28643 19343 28677
rect 19377 28643 19389 28677
rect 19331 28627 19389 28643
rect 19789 29901 19847 29917
rect 19789 29867 19801 29901
rect 19835 29867 19847 29901
rect 19789 29833 19847 29867
rect 19789 29799 19801 29833
rect 19835 29799 19847 29833
rect 19789 29765 19847 29799
rect 19789 29731 19801 29765
rect 19835 29731 19847 29765
rect 19789 29697 19847 29731
rect 19789 29663 19801 29697
rect 19835 29663 19847 29697
rect 19789 29629 19847 29663
rect 19789 29595 19801 29629
rect 19835 29595 19847 29629
rect 19789 29561 19847 29595
rect 19789 29527 19801 29561
rect 19835 29527 19847 29561
rect 19789 29493 19847 29527
rect 19789 29459 19801 29493
rect 19835 29459 19847 29493
rect 19789 29425 19847 29459
rect 19789 29391 19801 29425
rect 19835 29391 19847 29425
rect 19789 29357 19847 29391
rect 19789 29323 19801 29357
rect 19835 29323 19847 29357
rect 19789 29289 19847 29323
rect 19789 29255 19801 29289
rect 19835 29255 19847 29289
rect 19789 29221 19847 29255
rect 19789 29187 19801 29221
rect 19835 29187 19847 29221
rect 19789 29153 19847 29187
rect 19789 29119 19801 29153
rect 19835 29119 19847 29153
rect 19789 29085 19847 29119
rect 19789 29051 19801 29085
rect 19835 29051 19847 29085
rect 19789 29017 19847 29051
rect 19789 28983 19801 29017
rect 19835 28983 19847 29017
rect 19789 28949 19847 28983
rect 19789 28915 19801 28949
rect 19835 28915 19847 28949
rect 19789 28881 19847 28915
rect 19789 28847 19801 28881
rect 19835 28847 19847 28881
rect 19789 28813 19847 28847
rect 19789 28779 19801 28813
rect 19835 28779 19847 28813
rect 19789 28745 19847 28779
rect 19789 28711 19801 28745
rect 19835 28711 19847 28745
rect 19789 28677 19847 28711
rect 19789 28643 19801 28677
rect 19835 28643 19847 28677
rect 19789 28627 19847 28643
rect 20247 29901 20305 29917
rect 20247 29867 20259 29901
rect 20293 29867 20305 29901
rect 20247 29833 20305 29867
rect 20247 29799 20259 29833
rect 20293 29799 20305 29833
rect 20247 29765 20305 29799
rect 20247 29731 20259 29765
rect 20293 29731 20305 29765
rect 20247 29697 20305 29731
rect 20247 29663 20259 29697
rect 20293 29663 20305 29697
rect 20247 29629 20305 29663
rect 20247 29595 20259 29629
rect 20293 29595 20305 29629
rect 20247 29561 20305 29595
rect 20247 29527 20259 29561
rect 20293 29527 20305 29561
rect 20247 29493 20305 29527
rect 20247 29459 20259 29493
rect 20293 29459 20305 29493
rect 20247 29425 20305 29459
rect 20247 29391 20259 29425
rect 20293 29391 20305 29425
rect 20247 29357 20305 29391
rect 20247 29323 20259 29357
rect 20293 29323 20305 29357
rect 20247 29289 20305 29323
rect 20247 29255 20259 29289
rect 20293 29255 20305 29289
rect 20247 29221 20305 29255
rect 20247 29187 20259 29221
rect 20293 29187 20305 29221
rect 20247 29153 20305 29187
rect 20247 29119 20259 29153
rect 20293 29119 20305 29153
rect 20247 29085 20305 29119
rect 20247 29051 20259 29085
rect 20293 29051 20305 29085
rect 20247 29017 20305 29051
rect 20247 28983 20259 29017
rect 20293 28983 20305 29017
rect 20247 28949 20305 28983
rect 20247 28915 20259 28949
rect 20293 28915 20305 28949
rect 20247 28881 20305 28915
rect 20247 28847 20259 28881
rect 20293 28847 20305 28881
rect 20247 28813 20305 28847
rect 20247 28779 20259 28813
rect 20293 28779 20305 28813
rect 20247 28745 20305 28779
rect 20247 28711 20259 28745
rect 20293 28711 20305 28745
rect 20247 28677 20305 28711
rect 20247 28643 20259 28677
rect 20293 28643 20305 28677
rect 20247 28627 20305 28643
rect 20705 29901 20763 29917
rect 20705 29867 20717 29901
rect 20751 29867 20763 29901
rect 20705 29833 20763 29867
rect 20705 29799 20717 29833
rect 20751 29799 20763 29833
rect 20705 29765 20763 29799
rect 20705 29731 20717 29765
rect 20751 29731 20763 29765
rect 20705 29697 20763 29731
rect 20705 29663 20717 29697
rect 20751 29663 20763 29697
rect 20705 29629 20763 29663
rect 20705 29595 20717 29629
rect 20751 29595 20763 29629
rect 20705 29561 20763 29595
rect 20705 29527 20717 29561
rect 20751 29527 20763 29561
rect 20705 29493 20763 29527
rect 20705 29459 20717 29493
rect 20751 29459 20763 29493
rect 20705 29425 20763 29459
rect 20705 29391 20717 29425
rect 20751 29391 20763 29425
rect 20705 29357 20763 29391
rect 20705 29323 20717 29357
rect 20751 29323 20763 29357
rect 20705 29289 20763 29323
rect 20705 29255 20717 29289
rect 20751 29255 20763 29289
rect 20705 29221 20763 29255
rect 20705 29187 20717 29221
rect 20751 29187 20763 29221
rect 20705 29153 20763 29187
rect 20705 29119 20717 29153
rect 20751 29119 20763 29153
rect 20705 29085 20763 29119
rect 20705 29051 20717 29085
rect 20751 29051 20763 29085
rect 20705 29017 20763 29051
rect 20705 28983 20717 29017
rect 20751 28983 20763 29017
rect 20705 28949 20763 28983
rect 20705 28915 20717 28949
rect 20751 28915 20763 28949
rect 20705 28881 20763 28915
rect 20705 28847 20717 28881
rect 20751 28847 20763 28881
rect 20705 28813 20763 28847
rect 20705 28779 20717 28813
rect 20751 28779 20763 28813
rect 20705 28745 20763 28779
rect 20705 28711 20717 28745
rect 20751 28711 20763 28745
rect 20705 28677 20763 28711
rect 20705 28643 20717 28677
rect 20751 28643 20763 28677
rect 20705 28627 20763 28643
rect 21163 29901 21221 29917
rect 21163 29867 21175 29901
rect 21209 29867 21221 29901
rect 21163 29833 21221 29867
rect 21163 29799 21175 29833
rect 21209 29799 21221 29833
rect 21163 29765 21221 29799
rect 21163 29731 21175 29765
rect 21209 29731 21221 29765
rect 21163 29697 21221 29731
rect 21163 29663 21175 29697
rect 21209 29663 21221 29697
rect 21163 29629 21221 29663
rect 21163 29595 21175 29629
rect 21209 29595 21221 29629
rect 21163 29561 21221 29595
rect 21163 29527 21175 29561
rect 21209 29527 21221 29561
rect 21163 29493 21221 29527
rect 21163 29459 21175 29493
rect 21209 29459 21221 29493
rect 21163 29425 21221 29459
rect 21163 29391 21175 29425
rect 21209 29391 21221 29425
rect 21163 29357 21221 29391
rect 21163 29323 21175 29357
rect 21209 29323 21221 29357
rect 21163 29289 21221 29323
rect 21163 29255 21175 29289
rect 21209 29255 21221 29289
rect 21163 29221 21221 29255
rect 21163 29187 21175 29221
rect 21209 29187 21221 29221
rect 21163 29153 21221 29187
rect 21163 29119 21175 29153
rect 21209 29119 21221 29153
rect 21163 29085 21221 29119
rect 21163 29051 21175 29085
rect 21209 29051 21221 29085
rect 21163 29017 21221 29051
rect 21163 28983 21175 29017
rect 21209 28983 21221 29017
rect 21163 28949 21221 28983
rect 21163 28915 21175 28949
rect 21209 28915 21221 28949
rect 21163 28881 21221 28915
rect 21163 28847 21175 28881
rect 21209 28847 21221 28881
rect 21163 28813 21221 28847
rect 21163 28779 21175 28813
rect 21209 28779 21221 28813
rect 21163 28745 21221 28779
rect 21163 28711 21175 28745
rect 21209 28711 21221 28745
rect 21163 28677 21221 28711
rect 21163 28643 21175 28677
rect 21209 28643 21221 28677
rect 21163 28627 21221 28643
rect 21621 29901 21679 29917
rect 21621 29867 21633 29901
rect 21667 29867 21679 29901
rect 21621 29833 21679 29867
rect 21621 29799 21633 29833
rect 21667 29799 21679 29833
rect 21621 29765 21679 29799
rect 21621 29731 21633 29765
rect 21667 29731 21679 29765
rect 21621 29697 21679 29731
rect 21621 29663 21633 29697
rect 21667 29663 21679 29697
rect 21621 29629 21679 29663
rect 21621 29595 21633 29629
rect 21667 29595 21679 29629
rect 21621 29561 21679 29595
rect 21621 29527 21633 29561
rect 21667 29527 21679 29561
rect 21621 29493 21679 29527
rect 21621 29459 21633 29493
rect 21667 29459 21679 29493
rect 21621 29425 21679 29459
rect 21621 29391 21633 29425
rect 21667 29391 21679 29425
rect 21621 29357 21679 29391
rect 21621 29323 21633 29357
rect 21667 29323 21679 29357
rect 21621 29289 21679 29323
rect 21621 29255 21633 29289
rect 21667 29255 21679 29289
rect 21621 29221 21679 29255
rect 21621 29187 21633 29221
rect 21667 29187 21679 29221
rect 21621 29153 21679 29187
rect 21621 29119 21633 29153
rect 21667 29119 21679 29153
rect 21621 29085 21679 29119
rect 21621 29051 21633 29085
rect 21667 29051 21679 29085
rect 21621 29017 21679 29051
rect 21621 28983 21633 29017
rect 21667 28983 21679 29017
rect 21621 28949 21679 28983
rect 21621 28915 21633 28949
rect 21667 28915 21679 28949
rect 21621 28881 21679 28915
rect 21621 28847 21633 28881
rect 21667 28847 21679 28881
rect 21621 28813 21679 28847
rect 21621 28779 21633 28813
rect 21667 28779 21679 28813
rect 21621 28745 21679 28779
rect 21621 28711 21633 28745
rect 21667 28711 21679 28745
rect 21621 28677 21679 28711
rect 21621 28643 21633 28677
rect 21667 28643 21679 28677
rect 21621 28627 21679 28643
rect 22079 29901 22137 29917
rect 22079 29867 22091 29901
rect 22125 29867 22137 29901
rect 22079 29833 22137 29867
rect 22079 29799 22091 29833
rect 22125 29799 22137 29833
rect 22079 29765 22137 29799
rect 22079 29731 22091 29765
rect 22125 29731 22137 29765
rect 22079 29697 22137 29731
rect 22079 29663 22091 29697
rect 22125 29663 22137 29697
rect 22079 29629 22137 29663
rect 22079 29595 22091 29629
rect 22125 29595 22137 29629
rect 22079 29561 22137 29595
rect 22079 29527 22091 29561
rect 22125 29527 22137 29561
rect 22079 29493 22137 29527
rect 22079 29459 22091 29493
rect 22125 29459 22137 29493
rect 22079 29425 22137 29459
rect 22079 29391 22091 29425
rect 22125 29391 22137 29425
rect 22079 29357 22137 29391
rect 22079 29323 22091 29357
rect 22125 29323 22137 29357
rect 22079 29289 22137 29323
rect 22079 29255 22091 29289
rect 22125 29255 22137 29289
rect 22079 29221 22137 29255
rect 22079 29187 22091 29221
rect 22125 29187 22137 29221
rect 22079 29153 22137 29187
rect 22079 29119 22091 29153
rect 22125 29119 22137 29153
rect 22079 29085 22137 29119
rect 22079 29051 22091 29085
rect 22125 29051 22137 29085
rect 22079 29017 22137 29051
rect 22079 28983 22091 29017
rect 22125 28983 22137 29017
rect 22079 28949 22137 28983
rect 22079 28915 22091 28949
rect 22125 28915 22137 28949
rect 22079 28881 22137 28915
rect 22079 28847 22091 28881
rect 22125 28847 22137 28881
rect 22079 28813 22137 28847
rect 22079 28779 22091 28813
rect 22125 28779 22137 28813
rect 22079 28745 22137 28779
rect 22079 28711 22091 28745
rect 22125 28711 22137 28745
rect 22079 28677 22137 28711
rect 22079 28643 22091 28677
rect 22125 28643 22137 28677
rect 22079 28627 22137 28643
rect 22537 29901 22595 29917
rect 22537 29867 22549 29901
rect 22583 29867 22595 29901
rect 22537 29833 22595 29867
rect 22537 29799 22549 29833
rect 22583 29799 22595 29833
rect 22537 29765 22595 29799
rect 22537 29731 22549 29765
rect 22583 29731 22595 29765
rect 22537 29697 22595 29731
rect 22537 29663 22549 29697
rect 22583 29663 22595 29697
rect 22537 29629 22595 29663
rect 22537 29595 22549 29629
rect 22583 29595 22595 29629
rect 22537 29561 22595 29595
rect 22537 29527 22549 29561
rect 22583 29527 22595 29561
rect 22537 29493 22595 29527
rect 22537 29459 22549 29493
rect 22583 29459 22595 29493
rect 22537 29425 22595 29459
rect 22537 29391 22549 29425
rect 22583 29391 22595 29425
rect 22537 29357 22595 29391
rect 22537 29323 22549 29357
rect 22583 29323 22595 29357
rect 22537 29289 22595 29323
rect 22537 29255 22549 29289
rect 22583 29255 22595 29289
rect 22537 29221 22595 29255
rect 22537 29187 22549 29221
rect 22583 29187 22595 29221
rect 22537 29153 22595 29187
rect 22537 29119 22549 29153
rect 22583 29119 22595 29153
rect 22537 29085 22595 29119
rect 22537 29051 22549 29085
rect 22583 29051 22595 29085
rect 22537 29017 22595 29051
rect 22537 28983 22549 29017
rect 22583 28983 22595 29017
rect 22537 28949 22595 28983
rect 22537 28915 22549 28949
rect 22583 28915 22595 28949
rect 22537 28881 22595 28915
rect 22537 28847 22549 28881
rect 22583 28847 22595 28881
rect 22537 28813 22595 28847
rect 22537 28779 22549 28813
rect 22583 28779 22595 28813
rect 22537 28745 22595 28779
rect 22537 28711 22549 28745
rect 22583 28711 22595 28745
rect 22537 28677 22595 28711
rect 22537 28643 22549 28677
rect 22583 28643 22595 28677
rect 22537 28627 22595 28643
rect 22995 29901 23053 29917
rect 22995 29867 23007 29901
rect 23041 29867 23053 29901
rect 22995 29833 23053 29867
rect 22995 29799 23007 29833
rect 23041 29799 23053 29833
rect 22995 29765 23053 29799
rect 22995 29731 23007 29765
rect 23041 29731 23053 29765
rect 22995 29697 23053 29731
rect 22995 29663 23007 29697
rect 23041 29663 23053 29697
rect 22995 29629 23053 29663
rect 22995 29595 23007 29629
rect 23041 29595 23053 29629
rect 22995 29561 23053 29595
rect 22995 29527 23007 29561
rect 23041 29527 23053 29561
rect 22995 29493 23053 29527
rect 22995 29459 23007 29493
rect 23041 29459 23053 29493
rect 22995 29425 23053 29459
rect 22995 29391 23007 29425
rect 23041 29391 23053 29425
rect 22995 29357 23053 29391
rect 22995 29323 23007 29357
rect 23041 29323 23053 29357
rect 22995 29289 23053 29323
rect 22995 29255 23007 29289
rect 23041 29255 23053 29289
rect 22995 29221 23053 29255
rect 22995 29187 23007 29221
rect 23041 29187 23053 29221
rect 22995 29153 23053 29187
rect 22995 29119 23007 29153
rect 23041 29119 23053 29153
rect 22995 29085 23053 29119
rect 22995 29051 23007 29085
rect 23041 29051 23053 29085
rect 22995 29017 23053 29051
rect 22995 28983 23007 29017
rect 23041 28983 23053 29017
rect 22995 28949 23053 28983
rect 22995 28915 23007 28949
rect 23041 28915 23053 28949
rect 22995 28881 23053 28915
rect 22995 28847 23007 28881
rect 23041 28847 23053 28881
rect 22995 28813 23053 28847
rect 22995 28779 23007 28813
rect 23041 28779 23053 28813
rect 22995 28745 23053 28779
rect 22995 28711 23007 28745
rect 23041 28711 23053 28745
rect 22995 28677 23053 28711
rect 22995 28643 23007 28677
rect 23041 28643 23053 28677
rect 22995 28627 23053 28643
rect 23453 29901 23511 29917
rect 23453 29867 23465 29901
rect 23499 29867 23511 29901
rect 23453 29833 23511 29867
rect 23453 29799 23465 29833
rect 23499 29799 23511 29833
rect 23453 29765 23511 29799
rect 23453 29731 23465 29765
rect 23499 29731 23511 29765
rect 23453 29697 23511 29731
rect 23453 29663 23465 29697
rect 23499 29663 23511 29697
rect 23453 29629 23511 29663
rect 23453 29595 23465 29629
rect 23499 29595 23511 29629
rect 23453 29561 23511 29595
rect 23453 29527 23465 29561
rect 23499 29527 23511 29561
rect 23453 29493 23511 29527
rect 23453 29459 23465 29493
rect 23499 29459 23511 29493
rect 23453 29425 23511 29459
rect 23453 29391 23465 29425
rect 23499 29391 23511 29425
rect 23453 29357 23511 29391
rect 23453 29323 23465 29357
rect 23499 29323 23511 29357
rect 23453 29289 23511 29323
rect 23453 29255 23465 29289
rect 23499 29255 23511 29289
rect 23453 29221 23511 29255
rect 23453 29187 23465 29221
rect 23499 29187 23511 29221
rect 23453 29153 23511 29187
rect 23453 29119 23465 29153
rect 23499 29119 23511 29153
rect 23453 29085 23511 29119
rect 23453 29051 23465 29085
rect 23499 29051 23511 29085
rect 23453 29017 23511 29051
rect 23453 28983 23465 29017
rect 23499 28983 23511 29017
rect 23453 28949 23511 28983
rect 23453 28915 23465 28949
rect 23499 28915 23511 28949
rect 23453 28881 23511 28915
rect 23453 28847 23465 28881
rect 23499 28847 23511 28881
rect 23453 28813 23511 28847
rect 23453 28779 23465 28813
rect 23499 28779 23511 28813
rect 23453 28745 23511 28779
rect 23453 28711 23465 28745
rect 23499 28711 23511 28745
rect 23453 28677 23511 28711
rect 23453 28643 23465 28677
rect 23499 28643 23511 28677
rect 23453 28627 23511 28643
rect 23911 29901 23969 29917
rect 23911 29867 23923 29901
rect 23957 29867 23969 29901
rect 23911 29833 23969 29867
rect 23911 29799 23923 29833
rect 23957 29799 23969 29833
rect 23911 29765 23969 29799
rect 23911 29731 23923 29765
rect 23957 29731 23969 29765
rect 23911 29697 23969 29731
rect 23911 29663 23923 29697
rect 23957 29663 23969 29697
rect 23911 29629 23969 29663
rect 23911 29595 23923 29629
rect 23957 29595 23969 29629
rect 23911 29561 23969 29595
rect 23911 29527 23923 29561
rect 23957 29527 23969 29561
rect 23911 29493 23969 29527
rect 23911 29459 23923 29493
rect 23957 29459 23969 29493
rect 23911 29425 23969 29459
rect 23911 29391 23923 29425
rect 23957 29391 23969 29425
rect 23911 29357 23969 29391
rect 23911 29323 23923 29357
rect 23957 29323 23969 29357
rect 23911 29289 23969 29323
rect 23911 29255 23923 29289
rect 23957 29255 23969 29289
rect 23911 29221 23969 29255
rect 23911 29187 23923 29221
rect 23957 29187 23969 29221
rect 23911 29153 23969 29187
rect 23911 29119 23923 29153
rect 23957 29119 23969 29153
rect 23911 29085 23969 29119
rect 23911 29051 23923 29085
rect 23957 29051 23969 29085
rect 23911 29017 23969 29051
rect 23911 28983 23923 29017
rect 23957 28983 23969 29017
rect 23911 28949 23969 28983
rect 23911 28915 23923 28949
rect 23957 28915 23969 28949
rect 23911 28881 23969 28915
rect 23911 28847 23923 28881
rect 23957 28847 23969 28881
rect 23911 28813 23969 28847
rect 23911 28779 23923 28813
rect 23957 28779 23969 28813
rect 23911 28745 23969 28779
rect 23911 28711 23923 28745
rect 23957 28711 23969 28745
rect 23911 28677 23969 28711
rect 23911 28643 23923 28677
rect 23957 28643 23969 28677
rect 23911 28627 23969 28643
rect 24369 29901 24427 29917
rect 24369 29867 24381 29901
rect 24415 29867 24427 29901
rect 24369 29833 24427 29867
rect 24369 29799 24381 29833
rect 24415 29799 24427 29833
rect 24369 29765 24427 29799
rect 24369 29731 24381 29765
rect 24415 29731 24427 29765
rect 24369 29697 24427 29731
rect 24369 29663 24381 29697
rect 24415 29663 24427 29697
rect 24369 29629 24427 29663
rect 24369 29595 24381 29629
rect 24415 29595 24427 29629
rect 24369 29561 24427 29595
rect 24369 29527 24381 29561
rect 24415 29527 24427 29561
rect 24369 29493 24427 29527
rect 24369 29459 24381 29493
rect 24415 29459 24427 29493
rect 24369 29425 24427 29459
rect 24369 29391 24381 29425
rect 24415 29391 24427 29425
rect 24369 29357 24427 29391
rect 24369 29323 24381 29357
rect 24415 29323 24427 29357
rect 24369 29289 24427 29323
rect 24369 29255 24381 29289
rect 24415 29255 24427 29289
rect 24369 29221 24427 29255
rect 24369 29187 24381 29221
rect 24415 29187 24427 29221
rect 24369 29153 24427 29187
rect 24369 29119 24381 29153
rect 24415 29119 24427 29153
rect 24369 29085 24427 29119
rect 24369 29051 24381 29085
rect 24415 29051 24427 29085
rect 24369 29017 24427 29051
rect 24369 28983 24381 29017
rect 24415 28983 24427 29017
rect 24369 28949 24427 28983
rect 24369 28915 24381 28949
rect 24415 28915 24427 28949
rect 24369 28881 24427 28915
rect 24369 28847 24381 28881
rect 24415 28847 24427 28881
rect 24369 28813 24427 28847
rect 24369 28779 24381 28813
rect 24415 28779 24427 28813
rect 24369 28745 24427 28779
rect 24369 28711 24381 28745
rect 24415 28711 24427 28745
rect 24369 28677 24427 28711
rect 24369 28643 24381 28677
rect 24415 28643 24427 28677
rect 24369 28627 24427 28643
rect 24827 29901 24885 29917
rect 24827 29867 24839 29901
rect 24873 29867 24885 29901
rect 24827 29833 24885 29867
rect 24827 29799 24839 29833
rect 24873 29799 24885 29833
rect 24827 29765 24885 29799
rect 24827 29731 24839 29765
rect 24873 29731 24885 29765
rect 24827 29697 24885 29731
rect 24827 29663 24839 29697
rect 24873 29663 24885 29697
rect 24827 29629 24885 29663
rect 24827 29595 24839 29629
rect 24873 29595 24885 29629
rect 24827 29561 24885 29595
rect 24827 29527 24839 29561
rect 24873 29527 24885 29561
rect 24827 29493 24885 29527
rect 24827 29459 24839 29493
rect 24873 29459 24885 29493
rect 24827 29425 24885 29459
rect 24827 29391 24839 29425
rect 24873 29391 24885 29425
rect 24827 29357 24885 29391
rect 24827 29323 24839 29357
rect 24873 29323 24885 29357
rect 24827 29289 24885 29323
rect 24827 29255 24839 29289
rect 24873 29255 24885 29289
rect 24827 29221 24885 29255
rect 24827 29187 24839 29221
rect 24873 29187 24885 29221
rect 24827 29153 24885 29187
rect 24827 29119 24839 29153
rect 24873 29119 24885 29153
rect 24827 29085 24885 29119
rect 24827 29051 24839 29085
rect 24873 29051 24885 29085
rect 24827 29017 24885 29051
rect 24827 28983 24839 29017
rect 24873 28983 24885 29017
rect 24827 28949 24885 28983
rect 24827 28915 24839 28949
rect 24873 28915 24885 28949
rect 24827 28881 24885 28915
rect 24827 28847 24839 28881
rect 24873 28847 24885 28881
rect 24827 28813 24885 28847
rect 24827 28779 24839 28813
rect 24873 28779 24885 28813
rect 24827 28745 24885 28779
rect 24827 28711 24839 28745
rect 24873 28711 24885 28745
rect 24827 28677 24885 28711
rect 24827 28643 24839 28677
rect 24873 28643 24885 28677
rect 24827 28627 24885 28643
rect 25285 29901 25343 29917
rect 25285 29867 25297 29901
rect 25331 29867 25343 29901
rect 25285 29833 25343 29867
rect 25285 29799 25297 29833
rect 25331 29799 25343 29833
rect 25285 29765 25343 29799
rect 25285 29731 25297 29765
rect 25331 29731 25343 29765
rect 25285 29697 25343 29731
rect 25285 29663 25297 29697
rect 25331 29663 25343 29697
rect 25285 29629 25343 29663
rect 25285 29595 25297 29629
rect 25331 29595 25343 29629
rect 25285 29561 25343 29595
rect 25285 29527 25297 29561
rect 25331 29527 25343 29561
rect 25285 29493 25343 29527
rect 25285 29459 25297 29493
rect 25331 29459 25343 29493
rect 25285 29425 25343 29459
rect 25285 29391 25297 29425
rect 25331 29391 25343 29425
rect 25285 29357 25343 29391
rect 25285 29323 25297 29357
rect 25331 29323 25343 29357
rect 25285 29289 25343 29323
rect 25285 29255 25297 29289
rect 25331 29255 25343 29289
rect 25285 29221 25343 29255
rect 25285 29187 25297 29221
rect 25331 29187 25343 29221
rect 25285 29153 25343 29187
rect 25285 29119 25297 29153
rect 25331 29119 25343 29153
rect 25285 29085 25343 29119
rect 25285 29051 25297 29085
rect 25331 29051 25343 29085
rect 25285 29017 25343 29051
rect 25285 28983 25297 29017
rect 25331 28983 25343 29017
rect 25285 28949 25343 28983
rect 25285 28915 25297 28949
rect 25331 28915 25343 28949
rect 25285 28881 25343 28915
rect 25285 28847 25297 28881
rect 25331 28847 25343 28881
rect 25285 28813 25343 28847
rect 25285 28779 25297 28813
rect 25331 28779 25343 28813
rect 25285 28745 25343 28779
rect 25285 28711 25297 28745
rect 25331 28711 25343 28745
rect 25285 28677 25343 28711
rect 25285 28643 25297 28677
rect 25331 28643 25343 28677
rect 25285 28627 25343 28643
rect 25743 29901 25801 29917
rect 25743 29867 25755 29901
rect 25789 29867 25801 29901
rect 25743 29833 25801 29867
rect 25743 29799 25755 29833
rect 25789 29799 25801 29833
rect 25743 29765 25801 29799
rect 25743 29731 25755 29765
rect 25789 29731 25801 29765
rect 25743 29697 25801 29731
rect 25743 29663 25755 29697
rect 25789 29663 25801 29697
rect 25743 29629 25801 29663
rect 25743 29595 25755 29629
rect 25789 29595 25801 29629
rect 25743 29561 25801 29595
rect 25743 29527 25755 29561
rect 25789 29527 25801 29561
rect 25743 29493 25801 29527
rect 25743 29459 25755 29493
rect 25789 29459 25801 29493
rect 25743 29425 25801 29459
rect 25743 29391 25755 29425
rect 25789 29391 25801 29425
rect 25743 29357 25801 29391
rect 25743 29323 25755 29357
rect 25789 29323 25801 29357
rect 25743 29289 25801 29323
rect 25743 29255 25755 29289
rect 25789 29255 25801 29289
rect 25743 29221 25801 29255
rect 25743 29187 25755 29221
rect 25789 29187 25801 29221
rect 25743 29153 25801 29187
rect 25743 29119 25755 29153
rect 25789 29119 25801 29153
rect 25743 29085 25801 29119
rect 25743 29051 25755 29085
rect 25789 29051 25801 29085
rect 25743 29017 25801 29051
rect 25743 28983 25755 29017
rect 25789 28983 25801 29017
rect 25743 28949 25801 28983
rect 25743 28915 25755 28949
rect 25789 28915 25801 28949
rect 25743 28881 25801 28915
rect 25743 28847 25755 28881
rect 25789 28847 25801 28881
rect 25743 28813 25801 28847
rect 25743 28779 25755 28813
rect 25789 28779 25801 28813
rect 25743 28745 25801 28779
rect 25743 28711 25755 28745
rect 25789 28711 25801 28745
rect 25743 28677 25801 28711
rect 25743 28643 25755 28677
rect 25789 28643 25801 28677
rect 25743 28627 25801 28643
rect 26201 29901 26259 29917
rect 26201 29867 26213 29901
rect 26247 29867 26259 29901
rect 26201 29833 26259 29867
rect 26201 29799 26213 29833
rect 26247 29799 26259 29833
rect 26201 29765 26259 29799
rect 26201 29731 26213 29765
rect 26247 29731 26259 29765
rect 26201 29697 26259 29731
rect 26201 29663 26213 29697
rect 26247 29663 26259 29697
rect 26201 29629 26259 29663
rect 26201 29595 26213 29629
rect 26247 29595 26259 29629
rect 26201 29561 26259 29595
rect 26201 29527 26213 29561
rect 26247 29527 26259 29561
rect 26201 29493 26259 29527
rect 26201 29459 26213 29493
rect 26247 29459 26259 29493
rect 26201 29425 26259 29459
rect 26201 29391 26213 29425
rect 26247 29391 26259 29425
rect 26201 29357 26259 29391
rect 26201 29323 26213 29357
rect 26247 29323 26259 29357
rect 26201 29289 26259 29323
rect 26201 29255 26213 29289
rect 26247 29255 26259 29289
rect 26201 29221 26259 29255
rect 26201 29187 26213 29221
rect 26247 29187 26259 29221
rect 26201 29153 26259 29187
rect 26201 29119 26213 29153
rect 26247 29119 26259 29153
rect 26201 29085 26259 29119
rect 26201 29051 26213 29085
rect 26247 29051 26259 29085
rect 26201 29017 26259 29051
rect 26201 28983 26213 29017
rect 26247 28983 26259 29017
rect 26201 28949 26259 28983
rect 26201 28915 26213 28949
rect 26247 28915 26259 28949
rect 26201 28881 26259 28915
rect 26201 28847 26213 28881
rect 26247 28847 26259 28881
rect 26201 28813 26259 28847
rect 26201 28779 26213 28813
rect 26247 28779 26259 28813
rect 26201 28745 26259 28779
rect 26201 28711 26213 28745
rect 26247 28711 26259 28745
rect 26201 28677 26259 28711
rect 26201 28643 26213 28677
rect 26247 28643 26259 28677
rect 26201 28627 26259 28643
rect 26659 29901 26717 29917
rect 26659 29867 26671 29901
rect 26705 29867 26717 29901
rect 26659 29833 26717 29867
rect 26659 29799 26671 29833
rect 26705 29799 26717 29833
rect 26659 29765 26717 29799
rect 26659 29731 26671 29765
rect 26705 29731 26717 29765
rect 26659 29697 26717 29731
rect 26659 29663 26671 29697
rect 26705 29663 26717 29697
rect 26659 29629 26717 29663
rect 26659 29595 26671 29629
rect 26705 29595 26717 29629
rect 26659 29561 26717 29595
rect 26659 29527 26671 29561
rect 26705 29527 26717 29561
rect 26659 29493 26717 29527
rect 26659 29459 26671 29493
rect 26705 29459 26717 29493
rect 26659 29425 26717 29459
rect 26659 29391 26671 29425
rect 26705 29391 26717 29425
rect 26659 29357 26717 29391
rect 26659 29323 26671 29357
rect 26705 29323 26717 29357
rect 26659 29289 26717 29323
rect 26659 29255 26671 29289
rect 26705 29255 26717 29289
rect 26659 29221 26717 29255
rect 26659 29187 26671 29221
rect 26705 29187 26717 29221
rect 26659 29153 26717 29187
rect 26659 29119 26671 29153
rect 26705 29119 26717 29153
rect 26659 29085 26717 29119
rect 26659 29051 26671 29085
rect 26705 29051 26717 29085
rect 26659 29017 26717 29051
rect 26659 28983 26671 29017
rect 26705 28983 26717 29017
rect 26659 28949 26717 28983
rect 26659 28915 26671 28949
rect 26705 28915 26717 28949
rect 26659 28881 26717 28915
rect 26659 28847 26671 28881
rect 26705 28847 26717 28881
rect 26659 28813 26717 28847
rect 26659 28779 26671 28813
rect 26705 28779 26717 28813
rect 26659 28745 26717 28779
rect 26659 28711 26671 28745
rect 26705 28711 26717 28745
rect 26659 28677 26717 28711
rect 26659 28643 26671 28677
rect 26705 28643 26717 28677
rect 26659 28627 26717 28643
rect 27117 29901 27175 29917
rect 27117 29867 27129 29901
rect 27163 29867 27175 29901
rect 27117 29833 27175 29867
rect 27117 29799 27129 29833
rect 27163 29799 27175 29833
rect 27117 29765 27175 29799
rect 27117 29731 27129 29765
rect 27163 29731 27175 29765
rect 27117 29697 27175 29731
rect 27117 29663 27129 29697
rect 27163 29663 27175 29697
rect 27117 29629 27175 29663
rect 27117 29595 27129 29629
rect 27163 29595 27175 29629
rect 27117 29561 27175 29595
rect 27117 29527 27129 29561
rect 27163 29527 27175 29561
rect 27117 29493 27175 29527
rect 27117 29459 27129 29493
rect 27163 29459 27175 29493
rect 27117 29425 27175 29459
rect 27117 29391 27129 29425
rect 27163 29391 27175 29425
rect 27117 29357 27175 29391
rect 27117 29323 27129 29357
rect 27163 29323 27175 29357
rect 27117 29289 27175 29323
rect 27117 29255 27129 29289
rect 27163 29255 27175 29289
rect 27117 29221 27175 29255
rect 27117 29187 27129 29221
rect 27163 29187 27175 29221
rect 27117 29153 27175 29187
rect 27117 29119 27129 29153
rect 27163 29119 27175 29153
rect 27117 29085 27175 29119
rect 27117 29051 27129 29085
rect 27163 29051 27175 29085
rect 27117 29017 27175 29051
rect 27117 28983 27129 29017
rect 27163 28983 27175 29017
rect 27117 28949 27175 28983
rect 27117 28915 27129 28949
rect 27163 28915 27175 28949
rect 27117 28881 27175 28915
rect 27117 28847 27129 28881
rect 27163 28847 27175 28881
rect 27117 28813 27175 28847
rect 27117 28779 27129 28813
rect 27163 28779 27175 28813
rect 27117 28745 27175 28779
rect 27117 28711 27129 28745
rect 27163 28711 27175 28745
rect 27117 28677 27175 28711
rect 27117 28643 27129 28677
rect 27163 28643 27175 28677
rect 27117 28627 27175 28643
rect 27575 29901 27633 29917
rect 27575 29867 27587 29901
rect 27621 29867 27633 29901
rect 27575 29833 27633 29867
rect 27575 29799 27587 29833
rect 27621 29799 27633 29833
rect 27575 29765 27633 29799
rect 27575 29731 27587 29765
rect 27621 29731 27633 29765
rect 27575 29697 27633 29731
rect 27575 29663 27587 29697
rect 27621 29663 27633 29697
rect 27575 29629 27633 29663
rect 27575 29595 27587 29629
rect 27621 29595 27633 29629
rect 27575 29561 27633 29595
rect 27575 29527 27587 29561
rect 27621 29527 27633 29561
rect 27575 29493 27633 29527
rect 27575 29459 27587 29493
rect 27621 29459 27633 29493
rect 27575 29425 27633 29459
rect 27575 29391 27587 29425
rect 27621 29391 27633 29425
rect 27575 29357 27633 29391
rect 27575 29323 27587 29357
rect 27621 29323 27633 29357
rect 27575 29289 27633 29323
rect 27575 29255 27587 29289
rect 27621 29255 27633 29289
rect 27575 29221 27633 29255
rect 27575 29187 27587 29221
rect 27621 29187 27633 29221
rect 27575 29153 27633 29187
rect 27575 29119 27587 29153
rect 27621 29119 27633 29153
rect 27575 29085 27633 29119
rect 27575 29051 27587 29085
rect 27621 29051 27633 29085
rect 27575 29017 27633 29051
rect 27575 28983 27587 29017
rect 27621 28983 27633 29017
rect 27575 28949 27633 28983
rect 27575 28915 27587 28949
rect 27621 28915 27633 28949
rect 27575 28881 27633 28915
rect 27575 28847 27587 28881
rect 27621 28847 27633 28881
rect 27575 28813 27633 28847
rect 27575 28779 27587 28813
rect 27621 28779 27633 28813
rect 27575 28745 27633 28779
rect 27575 28711 27587 28745
rect 27621 28711 27633 28745
rect 27575 28677 27633 28711
rect 27575 28643 27587 28677
rect 27621 28643 27633 28677
rect 27575 28627 27633 28643
rect 28033 29901 28091 29917
rect 28033 29867 28045 29901
rect 28079 29867 28091 29901
rect 28033 29833 28091 29867
rect 28033 29799 28045 29833
rect 28079 29799 28091 29833
rect 28033 29765 28091 29799
rect 28033 29731 28045 29765
rect 28079 29731 28091 29765
rect 28033 29697 28091 29731
rect 28033 29663 28045 29697
rect 28079 29663 28091 29697
rect 28033 29629 28091 29663
rect 28033 29595 28045 29629
rect 28079 29595 28091 29629
rect 28033 29561 28091 29595
rect 28033 29527 28045 29561
rect 28079 29527 28091 29561
rect 28033 29493 28091 29527
rect 28033 29459 28045 29493
rect 28079 29459 28091 29493
rect 28033 29425 28091 29459
rect 28033 29391 28045 29425
rect 28079 29391 28091 29425
rect 28033 29357 28091 29391
rect 28033 29323 28045 29357
rect 28079 29323 28091 29357
rect 28033 29289 28091 29323
rect 28033 29255 28045 29289
rect 28079 29255 28091 29289
rect 28033 29221 28091 29255
rect 28033 29187 28045 29221
rect 28079 29187 28091 29221
rect 28033 29153 28091 29187
rect 28033 29119 28045 29153
rect 28079 29119 28091 29153
rect 28033 29085 28091 29119
rect 28033 29051 28045 29085
rect 28079 29051 28091 29085
rect 28033 29017 28091 29051
rect 28033 28983 28045 29017
rect 28079 28983 28091 29017
rect 28033 28949 28091 28983
rect 28033 28915 28045 28949
rect 28079 28915 28091 28949
rect 28033 28881 28091 28915
rect 28033 28847 28045 28881
rect 28079 28847 28091 28881
rect 28033 28813 28091 28847
rect 28033 28779 28045 28813
rect 28079 28779 28091 28813
rect 28033 28745 28091 28779
rect 28033 28711 28045 28745
rect 28079 28711 28091 28745
rect 28033 28677 28091 28711
rect 28033 28643 28045 28677
rect 28079 28643 28091 28677
rect 28033 28627 28091 28643
rect 28491 29901 28549 29917
rect 28491 29867 28503 29901
rect 28537 29867 28549 29901
rect 28491 29833 28549 29867
rect 28491 29799 28503 29833
rect 28537 29799 28549 29833
rect 28491 29765 28549 29799
rect 28491 29731 28503 29765
rect 28537 29731 28549 29765
rect 28491 29697 28549 29731
rect 28491 29663 28503 29697
rect 28537 29663 28549 29697
rect 28491 29629 28549 29663
rect 28491 29595 28503 29629
rect 28537 29595 28549 29629
rect 28491 29561 28549 29595
rect 28491 29527 28503 29561
rect 28537 29527 28549 29561
rect 28491 29493 28549 29527
rect 28491 29459 28503 29493
rect 28537 29459 28549 29493
rect 28491 29425 28549 29459
rect 28491 29391 28503 29425
rect 28537 29391 28549 29425
rect 28491 29357 28549 29391
rect 28491 29323 28503 29357
rect 28537 29323 28549 29357
rect 28491 29289 28549 29323
rect 28491 29255 28503 29289
rect 28537 29255 28549 29289
rect 28491 29221 28549 29255
rect 28491 29187 28503 29221
rect 28537 29187 28549 29221
rect 28491 29153 28549 29187
rect 28491 29119 28503 29153
rect 28537 29119 28549 29153
rect 28491 29085 28549 29119
rect 28491 29051 28503 29085
rect 28537 29051 28549 29085
rect 28491 29017 28549 29051
rect 28491 28983 28503 29017
rect 28537 28983 28549 29017
rect 28491 28949 28549 28983
rect 28491 28915 28503 28949
rect 28537 28915 28549 28949
rect 28491 28881 28549 28915
rect 28491 28847 28503 28881
rect 28537 28847 28549 28881
rect 28491 28813 28549 28847
rect 28491 28779 28503 28813
rect 28537 28779 28549 28813
rect 28491 28745 28549 28779
rect 28491 28711 28503 28745
rect 28537 28711 28549 28745
rect 28491 28677 28549 28711
rect 28491 28643 28503 28677
rect 28537 28643 28549 28677
rect 28491 28627 28549 28643
rect 28949 29901 29007 29917
rect 28949 29867 28961 29901
rect 28995 29867 29007 29901
rect 28949 29833 29007 29867
rect 28949 29799 28961 29833
rect 28995 29799 29007 29833
rect 28949 29765 29007 29799
rect 28949 29731 28961 29765
rect 28995 29731 29007 29765
rect 28949 29697 29007 29731
rect 28949 29663 28961 29697
rect 28995 29663 29007 29697
rect 28949 29629 29007 29663
rect 28949 29595 28961 29629
rect 28995 29595 29007 29629
rect 28949 29561 29007 29595
rect 28949 29527 28961 29561
rect 28995 29527 29007 29561
rect 28949 29493 29007 29527
rect 28949 29459 28961 29493
rect 28995 29459 29007 29493
rect 28949 29425 29007 29459
rect 28949 29391 28961 29425
rect 28995 29391 29007 29425
rect 28949 29357 29007 29391
rect 28949 29323 28961 29357
rect 28995 29323 29007 29357
rect 28949 29289 29007 29323
rect 28949 29255 28961 29289
rect 28995 29255 29007 29289
rect 28949 29221 29007 29255
rect 28949 29187 28961 29221
rect 28995 29187 29007 29221
rect 28949 29153 29007 29187
rect 28949 29119 28961 29153
rect 28995 29119 29007 29153
rect 28949 29085 29007 29119
rect 28949 29051 28961 29085
rect 28995 29051 29007 29085
rect 28949 29017 29007 29051
rect 28949 28983 28961 29017
rect 28995 28983 29007 29017
rect 28949 28949 29007 28983
rect 28949 28915 28961 28949
rect 28995 28915 29007 28949
rect 28949 28881 29007 28915
rect 28949 28847 28961 28881
rect 28995 28847 29007 28881
rect 28949 28813 29007 28847
rect 28949 28779 28961 28813
rect 28995 28779 29007 28813
rect 28949 28745 29007 28779
rect 28949 28711 28961 28745
rect 28995 28711 29007 28745
rect 28949 28677 29007 28711
rect 28949 28643 28961 28677
rect 28995 28643 29007 28677
rect 28949 28627 29007 28643
rect 29407 29901 29465 29917
rect 29407 29867 29419 29901
rect 29453 29867 29465 29901
rect 29407 29833 29465 29867
rect 29407 29799 29419 29833
rect 29453 29799 29465 29833
rect 29407 29765 29465 29799
rect 29407 29731 29419 29765
rect 29453 29731 29465 29765
rect 29407 29697 29465 29731
rect 29407 29663 29419 29697
rect 29453 29663 29465 29697
rect 29407 29629 29465 29663
rect 29407 29595 29419 29629
rect 29453 29595 29465 29629
rect 29407 29561 29465 29595
rect 29407 29527 29419 29561
rect 29453 29527 29465 29561
rect 29407 29493 29465 29527
rect 29407 29459 29419 29493
rect 29453 29459 29465 29493
rect 29407 29425 29465 29459
rect 29407 29391 29419 29425
rect 29453 29391 29465 29425
rect 29407 29357 29465 29391
rect 29407 29323 29419 29357
rect 29453 29323 29465 29357
rect 29407 29289 29465 29323
rect 29407 29255 29419 29289
rect 29453 29255 29465 29289
rect 29407 29221 29465 29255
rect 29407 29187 29419 29221
rect 29453 29187 29465 29221
rect 29407 29153 29465 29187
rect 29407 29119 29419 29153
rect 29453 29119 29465 29153
rect 29407 29085 29465 29119
rect 29407 29051 29419 29085
rect 29453 29051 29465 29085
rect 29407 29017 29465 29051
rect 29407 28983 29419 29017
rect 29453 28983 29465 29017
rect 29407 28949 29465 28983
rect 29407 28915 29419 28949
rect 29453 28915 29465 28949
rect 29407 28881 29465 28915
rect 29407 28847 29419 28881
rect 29453 28847 29465 28881
rect 29407 28813 29465 28847
rect 29407 28779 29419 28813
rect 29453 28779 29465 28813
rect 29407 28745 29465 28779
rect 29407 28711 29419 28745
rect 29453 28711 29465 28745
rect 29407 28677 29465 28711
rect 29407 28643 29419 28677
rect 29453 28643 29465 28677
rect 29407 28627 29465 28643
rect 29865 29901 29923 29917
rect 29865 29867 29877 29901
rect 29911 29867 29923 29901
rect 29865 29833 29923 29867
rect 29865 29799 29877 29833
rect 29911 29799 29923 29833
rect 29865 29765 29923 29799
rect 29865 29731 29877 29765
rect 29911 29731 29923 29765
rect 29865 29697 29923 29731
rect 29865 29663 29877 29697
rect 29911 29663 29923 29697
rect 29865 29629 29923 29663
rect 29865 29595 29877 29629
rect 29911 29595 29923 29629
rect 29865 29561 29923 29595
rect 29865 29527 29877 29561
rect 29911 29527 29923 29561
rect 29865 29493 29923 29527
rect 29865 29459 29877 29493
rect 29911 29459 29923 29493
rect 29865 29425 29923 29459
rect 29865 29391 29877 29425
rect 29911 29391 29923 29425
rect 29865 29357 29923 29391
rect 29865 29323 29877 29357
rect 29911 29323 29923 29357
rect 29865 29289 29923 29323
rect 29865 29255 29877 29289
rect 29911 29255 29923 29289
rect 29865 29221 29923 29255
rect 29865 29187 29877 29221
rect 29911 29187 29923 29221
rect 29865 29153 29923 29187
rect 29865 29119 29877 29153
rect 29911 29119 29923 29153
rect 29865 29085 29923 29119
rect 29865 29051 29877 29085
rect 29911 29051 29923 29085
rect 29865 29017 29923 29051
rect 29865 28983 29877 29017
rect 29911 28983 29923 29017
rect 29865 28949 29923 28983
rect 29865 28915 29877 28949
rect 29911 28915 29923 28949
rect 29865 28881 29923 28915
rect 29865 28847 29877 28881
rect 29911 28847 29923 28881
rect 29865 28813 29923 28847
rect 29865 28779 29877 28813
rect 29911 28779 29923 28813
rect 29865 28745 29923 28779
rect 29865 28711 29877 28745
rect 29911 28711 29923 28745
rect 29865 28677 29923 28711
rect 29865 28643 29877 28677
rect 29911 28643 29923 28677
rect 29865 28627 29923 28643
rect 30323 29901 30381 29917
rect 30323 29867 30335 29901
rect 30369 29867 30381 29901
rect 30323 29833 30381 29867
rect 30323 29799 30335 29833
rect 30369 29799 30381 29833
rect 30323 29765 30381 29799
rect 30323 29731 30335 29765
rect 30369 29731 30381 29765
rect 30323 29697 30381 29731
rect 30323 29663 30335 29697
rect 30369 29663 30381 29697
rect 30323 29629 30381 29663
rect 30323 29595 30335 29629
rect 30369 29595 30381 29629
rect 30323 29561 30381 29595
rect 30323 29527 30335 29561
rect 30369 29527 30381 29561
rect 30323 29493 30381 29527
rect 30323 29459 30335 29493
rect 30369 29459 30381 29493
rect 30323 29425 30381 29459
rect 30323 29391 30335 29425
rect 30369 29391 30381 29425
rect 30323 29357 30381 29391
rect 30323 29323 30335 29357
rect 30369 29323 30381 29357
rect 30323 29289 30381 29323
rect 30323 29255 30335 29289
rect 30369 29255 30381 29289
rect 30323 29221 30381 29255
rect 30323 29187 30335 29221
rect 30369 29187 30381 29221
rect 30323 29153 30381 29187
rect 30323 29119 30335 29153
rect 30369 29119 30381 29153
rect 30323 29085 30381 29119
rect 30323 29051 30335 29085
rect 30369 29051 30381 29085
rect 30323 29017 30381 29051
rect 30323 28983 30335 29017
rect 30369 28983 30381 29017
rect 30323 28949 30381 28983
rect 30323 28915 30335 28949
rect 30369 28915 30381 28949
rect 30323 28881 30381 28915
rect 30323 28847 30335 28881
rect 30369 28847 30381 28881
rect 30323 28813 30381 28847
rect 30323 28779 30335 28813
rect 30369 28779 30381 28813
rect 30323 28745 30381 28779
rect 30323 28711 30335 28745
rect 30369 28711 30381 28745
rect 30323 28677 30381 28711
rect 30323 28643 30335 28677
rect 30369 28643 30381 28677
rect 30323 28627 30381 28643
rect 30781 29901 30839 29917
rect 30781 29867 30793 29901
rect 30827 29867 30839 29901
rect 30781 29833 30839 29867
rect 30781 29799 30793 29833
rect 30827 29799 30839 29833
rect 30781 29765 30839 29799
rect 30781 29731 30793 29765
rect 30827 29731 30839 29765
rect 30781 29697 30839 29731
rect 30781 29663 30793 29697
rect 30827 29663 30839 29697
rect 30781 29629 30839 29663
rect 30781 29595 30793 29629
rect 30827 29595 30839 29629
rect 30781 29561 30839 29595
rect 30781 29527 30793 29561
rect 30827 29527 30839 29561
rect 30781 29493 30839 29527
rect 30781 29459 30793 29493
rect 30827 29459 30839 29493
rect 30781 29425 30839 29459
rect 30781 29391 30793 29425
rect 30827 29391 30839 29425
rect 30781 29357 30839 29391
rect 30781 29323 30793 29357
rect 30827 29323 30839 29357
rect 30781 29289 30839 29323
rect 30781 29255 30793 29289
rect 30827 29255 30839 29289
rect 30781 29221 30839 29255
rect 30781 29187 30793 29221
rect 30827 29187 30839 29221
rect 30781 29153 30839 29187
rect 30781 29119 30793 29153
rect 30827 29119 30839 29153
rect 30781 29085 30839 29119
rect 30781 29051 30793 29085
rect 30827 29051 30839 29085
rect 30781 29017 30839 29051
rect 30781 28983 30793 29017
rect 30827 28983 30839 29017
rect 30781 28949 30839 28983
rect 30781 28915 30793 28949
rect 30827 28915 30839 28949
rect 30781 28881 30839 28915
rect 30781 28847 30793 28881
rect 30827 28847 30839 28881
rect 30781 28813 30839 28847
rect 30781 28779 30793 28813
rect 30827 28779 30839 28813
rect 30781 28745 30839 28779
rect 30781 28711 30793 28745
rect 30827 28711 30839 28745
rect 30781 28677 30839 28711
rect 30781 28643 30793 28677
rect 30827 28643 30839 28677
rect 30781 28627 30839 28643
rect 31239 29901 31297 29917
rect 31239 29867 31251 29901
rect 31285 29867 31297 29901
rect 31239 29833 31297 29867
rect 31239 29799 31251 29833
rect 31285 29799 31297 29833
rect 31239 29765 31297 29799
rect 31239 29731 31251 29765
rect 31285 29731 31297 29765
rect 31239 29697 31297 29731
rect 31239 29663 31251 29697
rect 31285 29663 31297 29697
rect 31239 29629 31297 29663
rect 31239 29595 31251 29629
rect 31285 29595 31297 29629
rect 31239 29561 31297 29595
rect 31239 29527 31251 29561
rect 31285 29527 31297 29561
rect 31239 29493 31297 29527
rect 31239 29459 31251 29493
rect 31285 29459 31297 29493
rect 31239 29425 31297 29459
rect 31239 29391 31251 29425
rect 31285 29391 31297 29425
rect 31239 29357 31297 29391
rect 31239 29323 31251 29357
rect 31285 29323 31297 29357
rect 31239 29289 31297 29323
rect 31239 29255 31251 29289
rect 31285 29255 31297 29289
rect 31239 29221 31297 29255
rect 31239 29187 31251 29221
rect 31285 29187 31297 29221
rect 31239 29153 31297 29187
rect 31239 29119 31251 29153
rect 31285 29119 31297 29153
rect 31239 29085 31297 29119
rect 31239 29051 31251 29085
rect 31285 29051 31297 29085
rect 31239 29017 31297 29051
rect 31239 28983 31251 29017
rect 31285 28983 31297 29017
rect 31239 28949 31297 28983
rect 31239 28915 31251 28949
rect 31285 28915 31297 28949
rect 31239 28881 31297 28915
rect 31239 28847 31251 28881
rect 31285 28847 31297 28881
rect 31239 28813 31297 28847
rect 31239 28779 31251 28813
rect 31285 28779 31297 28813
rect 31239 28745 31297 28779
rect 31239 28711 31251 28745
rect 31285 28711 31297 28745
rect 31239 28677 31297 28711
rect 31239 28643 31251 28677
rect 31285 28643 31297 28677
rect 31239 28627 31297 28643
rect 31697 29901 31755 29917
rect 31697 29867 31709 29901
rect 31743 29867 31755 29901
rect 31697 29833 31755 29867
rect 31697 29799 31709 29833
rect 31743 29799 31755 29833
rect 31697 29765 31755 29799
rect 31697 29731 31709 29765
rect 31743 29731 31755 29765
rect 31697 29697 31755 29731
rect 31697 29663 31709 29697
rect 31743 29663 31755 29697
rect 31697 29629 31755 29663
rect 31697 29595 31709 29629
rect 31743 29595 31755 29629
rect 31697 29561 31755 29595
rect 31697 29527 31709 29561
rect 31743 29527 31755 29561
rect 31697 29493 31755 29527
rect 31697 29459 31709 29493
rect 31743 29459 31755 29493
rect 31697 29425 31755 29459
rect 31697 29391 31709 29425
rect 31743 29391 31755 29425
rect 31697 29357 31755 29391
rect 31697 29323 31709 29357
rect 31743 29323 31755 29357
rect 31697 29289 31755 29323
rect 31697 29255 31709 29289
rect 31743 29255 31755 29289
rect 31697 29221 31755 29255
rect 31697 29187 31709 29221
rect 31743 29187 31755 29221
rect 31697 29153 31755 29187
rect 31697 29119 31709 29153
rect 31743 29119 31755 29153
rect 31697 29085 31755 29119
rect 31697 29051 31709 29085
rect 31743 29051 31755 29085
rect 31697 29017 31755 29051
rect 31697 28983 31709 29017
rect 31743 28983 31755 29017
rect 31697 28949 31755 28983
rect 31697 28915 31709 28949
rect 31743 28915 31755 28949
rect 31697 28881 31755 28915
rect 31697 28847 31709 28881
rect 31743 28847 31755 28881
rect 31697 28813 31755 28847
rect 31697 28779 31709 28813
rect 31743 28779 31755 28813
rect 31697 28745 31755 28779
rect 31697 28711 31709 28745
rect 31743 28711 31755 28745
rect 31697 28677 31755 28711
rect 31697 28643 31709 28677
rect 31743 28643 31755 28677
rect 31697 28627 31755 28643
rect 32155 29901 32213 29917
rect 32155 29867 32167 29901
rect 32201 29867 32213 29901
rect 32155 29833 32213 29867
rect 32155 29799 32167 29833
rect 32201 29799 32213 29833
rect 32155 29765 32213 29799
rect 32155 29731 32167 29765
rect 32201 29731 32213 29765
rect 32155 29697 32213 29731
rect 32155 29663 32167 29697
rect 32201 29663 32213 29697
rect 32155 29629 32213 29663
rect 32155 29595 32167 29629
rect 32201 29595 32213 29629
rect 32155 29561 32213 29595
rect 32155 29527 32167 29561
rect 32201 29527 32213 29561
rect 32155 29493 32213 29527
rect 32155 29459 32167 29493
rect 32201 29459 32213 29493
rect 32155 29425 32213 29459
rect 32155 29391 32167 29425
rect 32201 29391 32213 29425
rect 32155 29357 32213 29391
rect 32155 29323 32167 29357
rect 32201 29323 32213 29357
rect 32155 29289 32213 29323
rect 32155 29255 32167 29289
rect 32201 29255 32213 29289
rect 32155 29221 32213 29255
rect 32155 29187 32167 29221
rect 32201 29187 32213 29221
rect 32155 29153 32213 29187
rect 32155 29119 32167 29153
rect 32201 29119 32213 29153
rect 32155 29085 32213 29119
rect 32155 29051 32167 29085
rect 32201 29051 32213 29085
rect 32155 29017 32213 29051
rect 32155 28983 32167 29017
rect 32201 28983 32213 29017
rect 32155 28949 32213 28983
rect 32155 28915 32167 28949
rect 32201 28915 32213 28949
rect 32155 28881 32213 28915
rect 32155 28847 32167 28881
rect 32201 28847 32213 28881
rect 32155 28813 32213 28847
rect 32155 28779 32167 28813
rect 32201 28779 32213 28813
rect 32155 28745 32213 28779
rect 32155 28711 32167 28745
rect 32201 28711 32213 28745
rect 32155 28677 32213 28711
rect 32155 28643 32167 28677
rect 32201 28643 32213 28677
rect 32155 28627 32213 28643
rect 32613 29901 32671 29917
rect 32613 29867 32625 29901
rect 32659 29867 32671 29901
rect 32613 29833 32671 29867
rect 32613 29799 32625 29833
rect 32659 29799 32671 29833
rect 32613 29765 32671 29799
rect 32613 29731 32625 29765
rect 32659 29731 32671 29765
rect 32613 29697 32671 29731
rect 32613 29663 32625 29697
rect 32659 29663 32671 29697
rect 32613 29629 32671 29663
rect 32613 29595 32625 29629
rect 32659 29595 32671 29629
rect 32613 29561 32671 29595
rect 32613 29527 32625 29561
rect 32659 29527 32671 29561
rect 32613 29493 32671 29527
rect 32613 29459 32625 29493
rect 32659 29459 32671 29493
rect 32613 29425 32671 29459
rect 32613 29391 32625 29425
rect 32659 29391 32671 29425
rect 32613 29357 32671 29391
rect 32613 29323 32625 29357
rect 32659 29323 32671 29357
rect 32613 29289 32671 29323
rect 32613 29255 32625 29289
rect 32659 29255 32671 29289
rect 32613 29221 32671 29255
rect 32613 29187 32625 29221
rect 32659 29187 32671 29221
rect 32613 29153 32671 29187
rect 32613 29119 32625 29153
rect 32659 29119 32671 29153
rect 32613 29085 32671 29119
rect 32613 29051 32625 29085
rect 32659 29051 32671 29085
rect 32613 29017 32671 29051
rect 32613 28983 32625 29017
rect 32659 28983 32671 29017
rect 32613 28949 32671 28983
rect 32613 28915 32625 28949
rect 32659 28915 32671 28949
rect 32613 28881 32671 28915
rect 32613 28847 32625 28881
rect 32659 28847 32671 28881
rect 32613 28813 32671 28847
rect 32613 28779 32625 28813
rect 32659 28779 32671 28813
rect 32613 28745 32671 28779
rect 32613 28711 32625 28745
rect 32659 28711 32671 28745
rect 32613 28677 32671 28711
rect 32613 28643 32625 28677
rect 32659 28643 32671 28677
rect 32613 28627 32671 28643
rect 33071 29901 33129 29917
rect 33071 29867 33083 29901
rect 33117 29867 33129 29901
rect 33071 29833 33129 29867
rect 33071 29799 33083 29833
rect 33117 29799 33129 29833
rect 33071 29765 33129 29799
rect 33071 29731 33083 29765
rect 33117 29731 33129 29765
rect 33071 29697 33129 29731
rect 33071 29663 33083 29697
rect 33117 29663 33129 29697
rect 33071 29629 33129 29663
rect 33071 29595 33083 29629
rect 33117 29595 33129 29629
rect 33071 29561 33129 29595
rect 33071 29527 33083 29561
rect 33117 29527 33129 29561
rect 33071 29493 33129 29527
rect 33071 29459 33083 29493
rect 33117 29459 33129 29493
rect 33071 29425 33129 29459
rect 33071 29391 33083 29425
rect 33117 29391 33129 29425
rect 33071 29357 33129 29391
rect 33071 29323 33083 29357
rect 33117 29323 33129 29357
rect 33071 29289 33129 29323
rect 33071 29255 33083 29289
rect 33117 29255 33129 29289
rect 33071 29221 33129 29255
rect 33071 29187 33083 29221
rect 33117 29187 33129 29221
rect 33071 29153 33129 29187
rect 33071 29119 33083 29153
rect 33117 29119 33129 29153
rect 33071 29085 33129 29119
rect 33071 29051 33083 29085
rect 33117 29051 33129 29085
rect 33071 29017 33129 29051
rect 33071 28983 33083 29017
rect 33117 28983 33129 29017
rect 33071 28949 33129 28983
rect 33071 28915 33083 28949
rect 33117 28915 33129 28949
rect 33071 28881 33129 28915
rect 33071 28847 33083 28881
rect 33117 28847 33129 28881
rect 33071 28813 33129 28847
rect 33071 28779 33083 28813
rect 33117 28779 33129 28813
rect 33071 28745 33129 28779
rect 33071 28711 33083 28745
rect 33117 28711 33129 28745
rect 33071 28677 33129 28711
rect 33071 28643 33083 28677
rect 33117 28643 33129 28677
rect 33071 28627 33129 28643
rect 33529 29901 33587 29917
rect 33529 29867 33541 29901
rect 33575 29867 33587 29901
rect 33529 29833 33587 29867
rect 33529 29799 33541 29833
rect 33575 29799 33587 29833
rect 33529 29765 33587 29799
rect 33529 29731 33541 29765
rect 33575 29731 33587 29765
rect 33529 29697 33587 29731
rect 33529 29663 33541 29697
rect 33575 29663 33587 29697
rect 33529 29629 33587 29663
rect 33529 29595 33541 29629
rect 33575 29595 33587 29629
rect 33529 29561 33587 29595
rect 33529 29527 33541 29561
rect 33575 29527 33587 29561
rect 33529 29493 33587 29527
rect 33529 29459 33541 29493
rect 33575 29459 33587 29493
rect 33529 29425 33587 29459
rect 33529 29391 33541 29425
rect 33575 29391 33587 29425
rect 33529 29357 33587 29391
rect 33529 29323 33541 29357
rect 33575 29323 33587 29357
rect 33529 29289 33587 29323
rect 33529 29255 33541 29289
rect 33575 29255 33587 29289
rect 33529 29221 33587 29255
rect 33529 29187 33541 29221
rect 33575 29187 33587 29221
rect 33529 29153 33587 29187
rect 33529 29119 33541 29153
rect 33575 29119 33587 29153
rect 33529 29085 33587 29119
rect 33529 29051 33541 29085
rect 33575 29051 33587 29085
rect 33529 29017 33587 29051
rect 33529 28983 33541 29017
rect 33575 28983 33587 29017
rect 33529 28949 33587 28983
rect 33529 28915 33541 28949
rect 33575 28915 33587 28949
rect 33529 28881 33587 28915
rect 33529 28847 33541 28881
rect 33575 28847 33587 28881
rect 33529 28813 33587 28847
rect 33529 28779 33541 28813
rect 33575 28779 33587 28813
rect 33529 28745 33587 28779
rect 33529 28711 33541 28745
rect 33575 28711 33587 28745
rect 33529 28677 33587 28711
rect 33529 28643 33541 28677
rect 33575 28643 33587 28677
rect 33529 28627 33587 28643
rect 34077 29901 34135 29917
rect 34077 29867 34089 29901
rect 34123 29867 34135 29901
rect 34077 29833 34135 29867
rect 34077 29799 34089 29833
rect 34123 29799 34135 29833
rect 34077 29765 34135 29799
rect 34077 29731 34089 29765
rect 34123 29731 34135 29765
rect 34077 29697 34135 29731
rect 34077 29663 34089 29697
rect 34123 29663 34135 29697
rect 34077 29629 34135 29663
rect 34077 29595 34089 29629
rect 34123 29595 34135 29629
rect 34077 29561 34135 29595
rect 34077 29527 34089 29561
rect 34123 29527 34135 29561
rect 34077 29493 34135 29527
rect 34077 29459 34089 29493
rect 34123 29459 34135 29493
rect 34077 29425 34135 29459
rect 34077 29391 34089 29425
rect 34123 29391 34135 29425
rect 34077 29357 34135 29391
rect 34077 29323 34089 29357
rect 34123 29323 34135 29357
rect 34077 29289 34135 29323
rect 34077 29255 34089 29289
rect 34123 29255 34135 29289
rect 34077 29221 34135 29255
rect 34077 29187 34089 29221
rect 34123 29187 34135 29221
rect 34077 29153 34135 29187
rect 34077 29119 34089 29153
rect 34123 29119 34135 29153
rect 34077 29085 34135 29119
rect 34077 29051 34089 29085
rect 34123 29051 34135 29085
rect 34077 29017 34135 29051
rect 34077 28983 34089 29017
rect 34123 28983 34135 29017
rect 34077 28949 34135 28983
rect 34077 28915 34089 28949
rect 34123 28915 34135 28949
rect 34077 28881 34135 28915
rect 34077 28847 34089 28881
rect 34123 28847 34135 28881
rect 34077 28813 34135 28847
rect 34077 28779 34089 28813
rect 34123 28779 34135 28813
rect 34077 28745 34135 28779
rect 34077 28711 34089 28745
rect 34123 28711 34135 28745
rect 34077 28677 34135 28711
rect 34077 28643 34089 28677
rect 34123 28643 34135 28677
rect 34077 28627 34135 28643
rect 34535 29901 34593 29917
rect 34535 29867 34547 29901
rect 34581 29867 34593 29901
rect 34535 29833 34593 29867
rect 34535 29799 34547 29833
rect 34581 29799 34593 29833
rect 34535 29765 34593 29799
rect 34535 29731 34547 29765
rect 34581 29731 34593 29765
rect 34535 29697 34593 29731
rect 34535 29663 34547 29697
rect 34581 29663 34593 29697
rect 34535 29629 34593 29663
rect 34535 29595 34547 29629
rect 34581 29595 34593 29629
rect 34535 29561 34593 29595
rect 34535 29527 34547 29561
rect 34581 29527 34593 29561
rect 34535 29493 34593 29527
rect 34535 29459 34547 29493
rect 34581 29459 34593 29493
rect 34535 29425 34593 29459
rect 34535 29391 34547 29425
rect 34581 29391 34593 29425
rect 34535 29357 34593 29391
rect 34535 29323 34547 29357
rect 34581 29323 34593 29357
rect 34535 29289 34593 29323
rect 34535 29255 34547 29289
rect 34581 29255 34593 29289
rect 34535 29221 34593 29255
rect 34535 29187 34547 29221
rect 34581 29187 34593 29221
rect 34535 29153 34593 29187
rect 34535 29119 34547 29153
rect 34581 29119 34593 29153
rect 34535 29085 34593 29119
rect 34535 29051 34547 29085
rect 34581 29051 34593 29085
rect 34535 29017 34593 29051
rect 34535 28983 34547 29017
rect 34581 28983 34593 29017
rect 34535 28949 34593 28983
rect 34535 28915 34547 28949
rect 34581 28915 34593 28949
rect 34535 28881 34593 28915
rect 34535 28847 34547 28881
rect 34581 28847 34593 28881
rect 34535 28813 34593 28847
rect 34535 28779 34547 28813
rect 34581 28779 34593 28813
rect 34535 28745 34593 28779
rect 34535 28711 34547 28745
rect 34581 28711 34593 28745
rect 34535 28677 34593 28711
rect 34535 28643 34547 28677
rect 34581 28643 34593 28677
rect 34535 28627 34593 28643
rect 34993 29901 35051 29917
rect 34993 29867 35005 29901
rect 35039 29867 35051 29901
rect 34993 29833 35051 29867
rect 34993 29799 35005 29833
rect 35039 29799 35051 29833
rect 34993 29765 35051 29799
rect 34993 29731 35005 29765
rect 35039 29731 35051 29765
rect 34993 29697 35051 29731
rect 34993 29663 35005 29697
rect 35039 29663 35051 29697
rect 34993 29629 35051 29663
rect 34993 29595 35005 29629
rect 35039 29595 35051 29629
rect 34993 29561 35051 29595
rect 34993 29527 35005 29561
rect 35039 29527 35051 29561
rect 34993 29493 35051 29527
rect 34993 29459 35005 29493
rect 35039 29459 35051 29493
rect 34993 29425 35051 29459
rect 34993 29391 35005 29425
rect 35039 29391 35051 29425
rect 34993 29357 35051 29391
rect 34993 29323 35005 29357
rect 35039 29323 35051 29357
rect 34993 29289 35051 29323
rect 34993 29255 35005 29289
rect 35039 29255 35051 29289
rect 34993 29221 35051 29255
rect 34993 29187 35005 29221
rect 35039 29187 35051 29221
rect 34993 29153 35051 29187
rect 34993 29119 35005 29153
rect 35039 29119 35051 29153
rect 34993 29085 35051 29119
rect 34993 29051 35005 29085
rect 35039 29051 35051 29085
rect 34993 29017 35051 29051
rect 34993 28983 35005 29017
rect 35039 28983 35051 29017
rect 34993 28949 35051 28983
rect 34993 28915 35005 28949
rect 35039 28915 35051 28949
rect 34993 28881 35051 28915
rect 34993 28847 35005 28881
rect 35039 28847 35051 28881
rect 34993 28813 35051 28847
rect 34993 28779 35005 28813
rect 35039 28779 35051 28813
rect 34993 28745 35051 28779
rect 34993 28711 35005 28745
rect 35039 28711 35051 28745
rect 34993 28677 35051 28711
rect 34993 28643 35005 28677
rect 35039 28643 35051 28677
rect 34993 28627 35051 28643
rect 35451 29901 35509 29917
rect 35451 29867 35463 29901
rect 35497 29867 35509 29901
rect 35451 29833 35509 29867
rect 35451 29799 35463 29833
rect 35497 29799 35509 29833
rect 35451 29765 35509 29799
rect 35451 29731 35463 29765
rect 35497 29731 35509 29765
rect 35451 29697 35509 29731
rect 35451 29663 35463 29697
rect 35497 29663 35509 29697
rect 35451 29629 35509 29663
rect 35451 29595 35463 29629
rect 35497 29595 35509 29629
rect 35451 29561 35509 29595
rect 35451 29527 35463 29561
rect 35497 29527 35509 29561
rect 35451 29493 35509 29527
rect 35451 29459 35463 29493
rect 35497 29459 35509 29493
rect 35451 29425 35509 29459
rect 35451 29391 35463 29425
rect 35497 29391 35509 29425
rect 35451 29357 35509 29391
rect 35451 29323 35463 29357
rect 35497 29323 35509 29357
rect 35451 29289 35509 29323
rect 35451 29255 35463 29289
rect 35497 29255 35509 29289
rect 35451 29221 35509 29255
rect 35451 29187 35463 29221
rect 35497 29187 35509 29221
rect 35451 29153 35509 29187
rect 35451 29119 35463 29153
rect 35497 29119 35509 29153
rect 35451 29085 35509 29119
rect 35451 29051 35463 29085
rect 35497 29051 35509 29085
rect 35451 29017 35509 29051
rect 35451 28983 35463 29017
rect 35497 28983 35509 29017
rect 35451 28949 35509 28983
rect 35451 28915 35463 28949
rect 35497 28915 35509 28949
rect 35451 28881 35509 28915
rect 35451 28847 35463 28881
rect 35497 28847 35509 28881
rect 35451 28813 35509 28847
rect 35451 28779 35463 28813
rect 35497 28779 35509 28813
rect 35451 28745 35509 28779
rect 35451 28711 35463 28745
rect 35497 28711 35509 28745
rect 35451 28677 35509 28711
rect 35451 28643 35463 28677
rect 35497 28643 35509 28677
rect 35451 28627 35509 28643
rect 35909 29901 35967 29917
rect 35909 29867 35921 29901
rect 35955 29867 35967 29901
rect 35909 29833 35967 29867
rect 35909 29799 35921 29833
rect 35955 29799 35967 29833
rect 35909 29765 35967 29799
rect 35909 29731 35921 29765
rect 35955 29731 35967 29765
rect 35909 29697 35967 29731
rect 35909 29663 35921 29697
rect 35955 29663 35967 29697
rect 35909 29629 35967 29663
rect 35909 29595 35921 29629
rect 35955 29595 35967 29629
rect 35909 29561 35967 29595
rect 35909 29527 35921 29561
rect 35955 29527 35967 29561
rect 35909 29493 35967 29527
rect 35909 29459 35921 29493
rect 35955 29459 35967 29493
rect 35909 29425 35967 29459
rect 35909 29391 35921 29425
rect 35955 29391 35967 29425
rect 35909 29357 35967 29391
rect 35909 29323 35921 29357
rect 35955 29323 35967 29357
rect 35909 29289 35967 29323
rect 35909 29255 35921 29289
rect 35955 29255 35967 29289
rect 35909 29221 35967 29255
rect 35909 29187 35921 29221
rect 35955 29187 35967 29221
rect 35909 29153 35967 29187
rect 35909 29119 35921 29153
rect 35955 29119 35967 29153
rect 35909 29085 35967 29119
rect 35909 29051 35921 29085
rect 35955 29051 35967 29085
rect 35909 29017 35967 29051
rect 35909 28983 35921 29017
rect 35955 28983 35967 29017
rect 35909 28949 35967 28983
rect 35909 28915 35921 28949
rect 35955 28915 35967 28949
rect 35909 28881 35967 28915
rect 35909 28847 35921 28881
rect 35955 28847 35967 28881
rect 35909 28813 35967 28847
rect 35909 28779 35921 28813
rect 35955 28779 35967 28813
rect 35909 28745 35967 28779
rect 35909 28711 35921 28745
rect 35955 28711 35967 28745
rect 35909 28677 35967 28711
rect 35909 28643 35921 28677
rect 35955 28643 35967 28677
rect 35909 28627 35967 28643
rect 36367 29901 36425 29917
rect 36367 29867 36379 29901
rect 36413 29867 36425 29901
rect 36367 29833 36425 29867
rect 36367 29799 36379 29833
rect 36413 29799 36425 29833
rect 36367 29765 36425 29799
rect 36367 29731 36379 29765
rect 36413 29731 36425 29765
rect 36367 29697 36425 29731
rect 36367 29663 36379 29697
rect 36413 29663 36425 29697
rect 36367 29629 36425 29663
rect 36367 29595 36379 29629
rect 36413 29595 36425 29629
rect 36367 29561 36425 29595
rect 36367 29527 36379 29561
rect 36413 29527 36425 29561
rect 36367 29493 36425 29527
rect 36367 29459 36379 29493
rect 36413 29459 36425 29493
rect 36367 29425 36425 29459
rect 36367 29391 36379 29425
rect 36413 29391 36425 29425
rect 36367 29357 36425 29391
rect 36367 29323 36379 29357
rect 36413 29323 36425 29357
rect 36367 29289 36425 29323
rect 36367 29255 36379 29289
rect 36413 29255 36425 29289
rect 36367 29221 36425 29255
rect 36367 29187 36379 29221
rect 36413 29187 36425 29221
rect 36367 29153 36425 29187
rect 36367 29119 36379 29153
rect 36413 29119 36425 29153
rect 36367 29085 36425 29119
rect 36367 29051 36379 29085
rect 36413 29051 36425 29085
rect 36367 29017 36425 29051
rect 36367 28983 36379 29017
rect 36413 28983 36425 29017
rect 36367 28949 36425 28983
rect 36367 28915 36379 28949
rect 36413 28915 36425 28949
rect 36367 28881 36425 28915
rect 36367 28847 36379 28881
rect 36413 28847 36425 28881
rect 36367 28813 36425 28847
rect 36367 28779 36379 28813
rect 36413 28779 36425 28813
rect 36367 28745 36425 28779
rect 36367 28711 36379 28745
rect 36413 28711 36425 28745
rect 36367 28677 36425 28711
rect 36367 28643 36379 28677
rect 36413 28643 36425 28677
rect 36367 28627 36425 28643
rect 36825 29901 36883 29917
rect 36825 29867 36837 29901
rect 36871 29867 36883 29901
rect 36825 29833 36883 29867
rect 36825 29799 36837 29833
rect 36871 29799 36883 29833
rect 36825 29765 36883 29799
rect 36825 29731 36837 29765
rect 36871 29731 36883 29765
rect 36825 29697 36883 29731
rect 36825 29663 36837 29697
rect 36871 29663 36883 29697
rect 36825 29629 36883 29663
rect 36825 29595 36837 29629
rect 36871 29595 36883 29629
rect 36825 29561 36883 29595
rect 36825 29527 36837 29561
rect 36871 29527 36883 29561
rect 36825 29493 36883 29527
rect 36825 29459 36837 29493
rect 36871 29459 36883 29493
rect 36825 29425 36883 29459
rect 36825 29391 36837 29425
rect 36871 29391 36883 29425
rect 36825 29357 36883 29391
rect 36825 29323 36837 29357
rect 36871 29323 36883 29357
rect 36825 29289 36883 29323
rect 36825 29255 36837 29289
rect 36871 29255 36883 29289
rect 36825 29221 36883 29255
rect 36825 29187 36837 29221
rect 36871 29187 36883 29221
rect 36825 29153 36883 29187
rect 36825 29119 36837 29153
rect 36871 29119 36883 29153
rect 36825 29085 36883 29119
rect 36825 29051 36837 29085
rect 36871 29051 36883 29085
rect 36825 29017 36883 29051
rect 36825 28983 36837 29017
rect 36871 28983 36883 29017
rect 36825 28949 36883 28983
rect 36825 28915 36837 28949
rect 36871 28915 36883 28949
rect 36825 28881 36883 28915
rect 36825 28847 36837 28881
rect 36871 28847 36883 28881
rect 36825 28813 36883 28847
rect 36825 28779 36837 28813
rect 36871 28779 36883 28813
rect 36825 28745 36883 28779
rect 36825 28711 36837 28745
rect 36871 28711 36883 28745
rect 36825 28677 36883 28711
rect 36825 28643 36837 28677
rect 36871 28643 36883 28677
rect 36825 28627 36883 28643
rect 9577 26141 9635 26157
rect 9577 26107 9589 26141
rect 9623 26107 9635 26141
rect 9577 26073 9635 26107
rect 9577 26039 9589 26073
rect 9623 26039 9635 26073
rect 9577 26005 9635 26039
rect 9577 25971 9589 26005
rect 9623 25971 9635 26005
rect 9577 25937 9635 25971
rect 9577 25903 9589 25937
rect 9623 25903 9635 25937
rect 9577 25869 9635 25903
rect 9577 25835 9589 25869
rect 9623 25835 9635 25869
rect 9577 25801 9635 25835
rect 9577 25767 9589 25801
rect 9623 25767 9635 25801
rect 9577 25733 9635 25767
rect 9577 25699 9589 25733
rect 9623 25699 9635 25733
rect 9577 25665 9635 25699
rect 9577 25631 9589 25665
rect 9623 25631 9635 25665
rect 9577 25597 9635 25631
rect 9577 25563 9589 25597
rect 9623 25563 9635 25597
rect 9577 25529 9635 25563
rect 9577 25495 9589 25529
rect 9623 25495 9635 25529
rect 9577 25461 9635 25495
rect 9577 25427 9589 25461
rect 9623 25427 9635 25461
rect 9577 25393 9635 25427
rect 9577 25359 9589 25393
rect 9623 25359 9635 25393
rect 9577 25325 9635 25359
rect 9577 25291 9589 25325
rect 9623 25291 9635 25325
rect 9577 25257 9635 25291
rect 9577 25223 9589 25257
rect 9623 25223 9635 25257
rect 9577 25189 9635 25223
rect 9577 25155 9589 25189
rect 9623 25155 9635 25189
rect 9577 25121 9635 25155
rect 9577 25087 9589 25121
rect 9623 25087 9635 25121
rect 9577 25053 9635 25087
rect 9577 25019 9589 25053
rect 9623 25019 9635 25053
rect 9577 24985 9635 25019
rect 9577 24951 9589 24985
rect 9623 24951 9635 24985
rect 9577 24917 9635 24951
rect 9577 24883 9589 24917
rect 9623 24883 9635 24917
rect 9577 24867 9635 24883
rect 10035 26141 10093 26157
rect 10035 26107 10047 26141
rect 10081 26107 10093 26141
rect 10035 26073 10093 26107
rect 10035 26039 10047 26073
rect 10081 26039 10093 26073
rect 10035 26005 10093 26039
rect 10035 25971 10047 26005
rect 10081 25971 10093 26005
rect 10035 25937 10093 25971
rect 10035 25903 10047 25937
rect 10081 25903 10093 25937
rect 10035 25869 10093 25903
rect 10035 25835 10047 25869
rect 10081 25835 10093 25869
rect 10035 25801 10093 25835
rect 10035 25767 10047 25801
rect 10081 25767 10093 25801
rect 10035 25733 10093 25767
rect 10035 25699 10047 25733
rect 10081 25699 10093 25733
rect 10035 25665 10093 25699
rect 10035 25631 10047 25665
rect 10081 25631 10093 25665
rect 10035 25597 10093 25631
rect 10035 25563 10047 25597
rect 10081 25563 10093 25597
rect 10035 25529 10093 25563
rect 10035 25495 10047 25529
rect 10081 25495 10093 25529
rect 10035 25461 10093 25495
rect 10035 25427 10047 25461
rect 10081 25427 10093 25461
rect 10035 25393 10093 25427
rect 10035 25359 10047 25393
rect 10081 25359 10093 25393
rect 10035 25325 10093 25359
rect 10035 25291 10047 25325
rect 10081 25291 10093 25325
rect 10035 25257 10093 25291
rect 10035 25223 10047 25257
rect 10081 25223 10093 25257
rect 10035 25189 10093 25223
rect 10035 25155 10047 25189
rect 10081 25155 10093 25189
rect 10035 25121 10093 25155
rect 10035 25087 10047 25121
rect 10081 25087 10093 25121
rect 10035 25053 10093 25087
rect 10035 25019 10047 25053
rect 10081 25019 10093 25053
rect 10035 24985 10093 25019
rect 10035 24951 10047 24985
rect 10081 24951 10093 24985
rect 10035 24917 10093 24951
rect 10035 24883 10047 24917
rect 10081 24883 10093 24917
rect 10035 24867 10093 24883
rect 10493 26141 10551 26157
rect 10493 26107 10505 26141
rect 10539 26107 10551 26141
rect 10493 26073 10551 26107
rect 10493 26039 10505 26073
rect 10539 26039 10551 26073
rect 10493 26005 10551 26039
rect 10493 25971 10505 26005
rect 10539 25971 10551 26005
rect 10493 25937 10551 25971
rect 10493 25903 10505 25937
rect 10539 25903 10551 25937
rect 10493 25869 10551 25903
rect 10493 25835 10505 25869
rect 10539 25835 10551 25869
rect 10493 25801 10551 25835
rect 10493 25767 10505 25801
rect 10539 25767 10551 25801
rect 10493 25733 10551 25767
rect 10493 25699 10505 25733
rect 10539 25699 10551 25733
rect 10493 25665 10551 25699
rect 10493 25631 10505 25665
rect 10539 25631 10551 25665
rect 10493 25597 10551 25631
rect 10493 25563 10505 25597
rect 10539 25563 10551 25597
rect 10493 25529 10551 25563
rect 10493 25495 10505 25529
rect 10539 25495 10551 25529
rect 10493 25461 10551 25495
rect 10493 25427 10505 25461
rect 10539 25427 10551 25461
rect 10493 25393 10551 25427
rect 10493 25359 10505 25393
rect 10539 25359 10551 25393
rect 10493 25325 10551 25359
rect 10493 25291 10505 25325
rect 10539 25291 10551 25325
rect 10493 25257 10551 25291
rect 10493 25223 10505 25257
rect 10539 25223 10551 25257
rect 10493 25189 10551 25223
rect 10493 25155 10505 25189
rect 10539 25155 10551 25189
rect 10493 25121 10551 25155
rect 10493 25087 10505 25121
rect 10539 25087 10551 25121
rect 10493 25053 10551 25087
rect 10493 25019 10505 25053
rect 10539 25019 10551 25053
rect 10493 24985 10551 25019
rect 10493 24951 10505 24985
rect 10539 24951 10551 24985
rect 10493 24917 10551 24951
rect 10493 24883 10505 24917
rect 10539 24883 10551 24917
rect 10493 24867 10551 24883
rect 10951 26141 11009 26157
rect 10951 26107 10963 26141
rect 10997 26107 11009 26141
rect 10951 26073 11009 26107
rect 10951 26039 10963 26073
rect 10997 26039 11009 26073
rect 10951 26005 11009 26039
rect 10951 25971 10963 26005
rect 10997 25971 11009 26005
rect 10951 25937 11009 25971
rect 10951 25903 10963 25937
rect 10997 25903 11009 25937
rect 10951 25869 11009 25903
rect 10951 25835 10963 25869
rect 10997 25835 11009 25869
rect 10951 25801 11009 25835
rect 10951 25767 10963 25801
rect 10997 25767 11009 25801
rect 10951 25733 11009 25767
rect 10951 25699 10963 25733
rect 10997 25699 11009 25733
rect 10951 25665 11009 25699
rect 10951 25631 10963 25665
rect 10997 25631 11009 25665
rect 10951 25597 11009 25631
rect 10951 25563 10963 25597
rect 10997 25563 11009 25597
rect 10951 25529 11009 25563
rect 10951 25495 10963 25529
rect 10997 25495 11009 25529
rect 10951 25461 11009 25495
rect 10951 25427 10963 25461
rect 10997 25427 11009 25461
rect 10951 25393 11009 25427
rect 10951 25359 10963 25393
rect 10997 25359 11009 25393
rect 10951 25325 11009 25359
rect 10951 25291 10963 25325
rect 10997 25291 11009 25325
rect 10951 25257 11009 25291
rect 10951 25223 10963 25257
rect 10997 25223 11009 25257
rect 10951 25189 11009 25223
rect 10951 25155 10963 25189
rect 10997 25155 11009 25189
rect 10951 25121 11009 25155
rect 10951 25087 10963 25121
rect 10997 25087 11009 25121
rect 10951 25053 11009 25087
rect 10951 25019 10963 25053
rect 10997 25019 11009 25053
rect 10951 24985 11009 25019
rect 10951 24951 10963 24985
rect 10997 24951 11009 24985
rect 10951 24917 11009 24951
rect 10951 24883 10963 24917
rect 10997 24883 11009 24917
rect 10951 24867 11009 24883
rect 11409 26141 11467 26157
rect 11409 26107 11421 26141
rect 11455 26107 11467 26141
rect 11409 26073 11467 26107
rect 11409 26039 11421 26073
rect 11455 26039 11467 26073
rect 11409 26005 11467 26039
rect 11409 25971 11421 26005
rect 11455 25971 11467 26005
rect 11409 25937 11467 25971
rect 11409 25903 11421 25937
rect 11455 25903 11467 25937
rect 11409 25869 11467 25903
rect 11409 25835 11421 25869
rect 11455 25835 11467 25869
rect 11409 25801 11467 25835
rect 11409 25767 11421 25801
rect 11455 25767 11467 25801
rect 11409 25733 11467 25767
rect 11409 25699 11421 25733
rect 11455 25699 11467 25733
rect 11409 25665 11467 25699
rect 11409 25631 11421 25665
rect 11455 25631 11467 25665
rect 11409 25597 11467 25631
rect 11409 25563 11421 25597
rect 11455 25563 11467 25597
rect 11409 25529 11467 25563
rect 11409 25495 11421 25529
rect 11455 25495 11467 25529
rect 11409 25461 11467 25495
rect 11409 25427 11421 25461
rect 11455 25427 11467 25461
rect 11409 25393 11467 25427
rect 11409 25359 11421 25393
rect 11455 25359 11467 25393
rect 11409 25325 11467 25359
rect 11409 25291 11421 25325
rect 11455 25291 11467 25325
rect 11409 25257 11467 25291
rect 11409 25223 11421 25257
rect 11455 25223 11467 25257
rect 11409 25189 11467 25223
rect 11409 25155 11421 25189
rect 11455 25155 11467 25189
rect 11409 25121 11467 25155
rect 11409 25087 11421 25121
rect 11455 25087 11467 25121
rect 11409 25053 11467 25087
rect 11409 25019 11421 25053
rect 11455 25019 11467 25053
rect 11409 24985 11467 25019
rect 11409 24951 11421 24985
rect 11455 24951 11467 24985
rect 11409 24917 11467 24951
rect 11409 24883 11421 24917
rect 11455 24883 11467 24917
rect 11409 24867 11467 24883
rect 11867 26141 11925 26157
rect 11867 26107 11879 26141
rect 11913 26107 11925 26141
rect 11867 26073 11925 26107
rect 11867 26039 11879 26073
rect 11913 26039 11925 26073
rect 11867 26005 11925 26039
rect 11867 25971 11879 26005
rect 11913 25971 11925 26005
rect 11867 25937 11925 25971
rect 11867 25903 11879 25937
rect 11913 25903 11925 25937
rect 11867 25869 11925 25903
rect 11867 25835 11879 25869
rect 11913 25835 11925 25869
rect 11867 25801 11925 25835
rect 11867 25767 11879 25801
rect 11913 25767 11925 25801
rect 11867 25733 11925 25767
rect 11867 25699 11879 25733
rect 11913 25699 11925 25733
rect 11867 25665 11925 25699
rect 11867 25631 11879 25665
rect 11913 25631 11925 25665
rect 11867 25597 11925 25631
rect 11867 25563 11879 25597
rect 11913 25563 11925 25597
rect 11867 25529 11925 25563
rect 11867 25495 11879 25529
rect 11913 25495 11925 25529
rect 11867 25461 11925 25495
rect 11867 25427 11879 25461
rect 11913 25427 11925 25461
rect 11867 25393 11925 25427
rect 11867 25359 11879 25393
rect 11913 25359 11925 25393
rect 11867 25325 11925 25359
rect 11867 25291 11879 25325
rect 11913 25291 11925 25325
rect 11867 25257 11925 25291
rect 11867 25223 11879 25257
rect 11913 25223 11925 25257
rect 11867 25189 11925 25223
rect 11867 25155 11879 25189
rect 11913 25155 11925 25189
rect 11867 25121 11925 25155
rect 11867 25087 11879 25121
rect 11913 25087 11925 25121
rect 11867 25053 11925 25087
rect 11867 25019 11879 25053
rect 11913 25019 11925 25053
rect 11867 24985 11925 25019
rect 11867 24951 11879 24985
rect 11913 24951 11925 24985
rect 11867 24917 11925 24951
rect 11867 24883 11879 24917
rect 11913 24883 11925 24917
rect 11867 24867 11925 24883
rect 12325 26141 12383 26157
rect 12325 26107 12337 26141
rect 12371 26107 12383 26141
rect 12325 26073 12383 26107
rect 12325 26039 12337 26073
rect 12371 26039 12383 26073
rect 12325 26005 12383 26039
rect 12325 25971 12337 26005
rect 12371 25971 12383 26005
rect 12325 25937 12383 25971
rect 12325 25903 12337 25937
rect 12371 25903 12383 25937
rect 12325 25869 12383 25903
rect 12325 25835 12337 25869
rect 12371 25835 12383 25869
rect 12325 25801 12383 25835
rect 12325 25767 12337 25801
rect 12371 25767 12383 25801
rect 12325 25733 12383 25767
rect 12325 25699 12337 25733
rect 12371 25699 12383 25733
rect 12325 25665 12383 25699
rect 12325 25631 12337 25665
rect 12371 25631 12383 25665
rect 12325 25597 12383 25631
rect 12325 25563 12337 25597
rect 12371 25563 12383 25597
rect 12325 25529 12383 25563
rect 12325 25495 12337 25529
rect 12371 25495 12383 25529
rect 12325 25461 12383 25495
rect 12325 25427 12337 25461
rect 12371 25427 12383 25461
rect 12325 25393 12383 25427
rect 12325 25359 12337 25393
rect 12371 25359 12383 25393
rect 12325 25325 12383 25359
rect 12325 25291 12337 25325
rect 12371 25291 12383 25325
rect 12325 25257 12383 25291
rect 12325 25223 12337 25257
rect 12371 25223 12383 25257
rect 12325 25189 12383 25223
rect 12325 25155 12337 25189
rect 12371 25155 12383 25189
rect 12325 25121 12383 25155
rect 12325 25087 12337 25121
rect 12371 25087 12383 25121
rect 12325 25053 12383 25087
rect 12325 25019 12337 25053
rect 12371 25019 12383 25053
rect 12325 24985 12383 25019
rect 12325 24951 12337 24985
rect 12371 24951 12383 24985
rect 12325 24917 12383 24951
rect 12325 24883 12337 24917
rect 12371 24883 12383 24917
rect 12325 24867 12383 24883
rect 12783 26141 12841 26157
rect 12783 26107 12795 26141
rect 12829 26107 12841 26141
rect 12783 26073 12841 26107
rect 12783 26039 12795 26073
rect 12829 26039 12841 26073
rect 12783 26005 12841 26039
rect 12783 25971 12795 26005
rect 12829 25971 12841 26005
rect 12783 25937 12841 25971
rect 12783 25903 12795 25937
rect 12829 25903 12841 25937
rect 12783 25869 12841 25903
rect 12783 25835 12795 25869
rect 12829 25835 12841 25869
rect 12783 25801 12841 25835
rect 12783 25767 12795 25801
rect 12829 25767 12841 25801
rect 12783 25733 12841 25767
rect 12783 25699 12795 25733
rect 12829 25699 12841 25733
rect 12783 25665 12841 25699
rect 12783 25631 12795 25665
rect 12829 25631 12841 25665
rect 12783 25597 12841 25631
rect 12783 25563 12795 25597
rect 12829 25563 12841 25597
rect 12783 25529 12841 25563
rect 12783 25495 12795 25529
rect 12829 25495 12841 25529
rect 12783 25461 12841 25495
rect 12783 25427 12795 25461
rect 12829 25427 12841 25461
rect 12783 25393 12841 25427
rect 12783 25359 12795 25393
rect 12829 25359 12841 25393
rect 12783 25325 12841 25359
rect 12783 25291 12795 25325
rect 12829 25291 12841 25325
rect 12783 25257 12841 25291
rect 12783 25223 12795 25257
rect 12829 25223 12841 25257
rect 12783 25189 12841 25223
rect 12783 25155 12795 25189
rect 12829 25155 12841 25189
rect 12783 25121 12841 25155
rect 12783 25087 12795 25121
rect 12829 25087 12841 25121
rect 12783 25053 12841 25087
rect 12783 25019 12795 25053
rect 12829 25019 12841 25053
rect 12783 24985 12841 25019
rect 12783 24951 12795 24985
rect 12829 24951 12841 24985
rect 12783 24917 12841 24951
rect 12783 24883 12795 24917
rect 12829 24883 12841 24917
rect 12783 24867 12841 24883
rect 13241 26141 13299 26157
rect 13241 26107 13253 26141
rect 13287 26107 13299 26141
rect 13241 26073 13299 26107
rect 13241 26039 13253 26073
rect 13287 26039 13299 26073
rect 13241 26005 13299 26039
rect 13241 25971 13253 26005
rect 13287 25971 13299 26005
rect 13241 25937 13299 25971
rect 13241 25903 13253 25937
rect 13287 25903 13299 25937
rect 13241 25869 13299 25903
rect 13241 25835 13253 25869
rect 13287 25835 13299 25869
rect 13241 25801 13299 25835
rect 13241 25767 13253 25801
rect 13287 25767 13299 25801
rect 13241 25733 13299 25767
rect 13241 25699 13253 25733
rect 13287 25699 13299 25733
rect 13241 25665 13299 25699
rect 13241 25631 13253 25665
rect 13287 25631 13299 25665
rect 13241 25597 13299 25631
rect 13241 25563 13253 25597
rect 13287 25563 13299 25597
rect 13241 25529 13299 25563
rect 13241 25495 13253 25529
rect 13287 25495 13299 25529
rect 13241 25461 13299 25495
rect 13241 25427 13253 25461
rect 13287 25427 13299 25461
rect 13241 25393 13299 25427
rect 13241 25359 13253 25393
rect 13287 25359 13299 25393
rect 13241 25325 13299 25359
rect 13241 25291 13253 25325
rect 13287 25291 13299 25325
rect 13241 25257 13299 25291
rect 13241 25223 13253 25257
rect 13287 25223 13299 25257
rect 13241 25189 13299 25223
rect 13241 25155 13253 25189
rect 13287 25155 13299 25189
rect 13241 25121 13299 25155
rect 13241 25087 13253 25121
rect 13287 25087 13299 25121
rect 13241 25053 13299 25087
rect 13241 25019 13253 25053
rect 13287 25019 13299 25053
rect 13241 24985 13299 25019
rect 13241 24951 13253 24985
rect 13287 24951 13299 24985
rect 13241 24917 13299 24951
rect 13241 24883 13253 24917
rect 13287 24883 13299 24917
rect 13241 24867 13299 24883
rect 13699 26141 13757 26157
rect 13699 26107 13711 26141
rect 13745 26107 13757 26141
rect 13699 26073 13757 26107
rect 13699 26039 13711 26073
rect 13745 26039 13757 26073
rect 13699 26005 13757 26039
rect 13699 25971 13711 26005
rect 13745 25971 13757 26005
rect 13699 25937 13757 25971
rect 13699 25903 13711 25937
rect 13745 25903 13757 25937
rect 13699 25869 13757 25903
rect 13699 25835 13711 25869
rect 13745 25835 13757 25869
rect 13699 25801 13757 25835
rect 13699 25767 13711 25801
rect 13745 25767 13757 25801
rect 13699 25733 13757 25767
rect 13699 25699 13711 25733
rect 13745 25699 13757 25733
rect 13699 25665 13757 25699
rect 13699 25631 13711 25665
rect 13745 25631 13757 25665
rect 13699 25597 13757 25631
rect 13699 25563 13711 25597
rect 13745 25563 13757 25597
rect 13699 25529 13757 25563
rect 13699 25495 13711 25529
rect 13745 25495 13757 25529
rect 13699 25461 13757 25495
rect 13699 25427 13711 25461
rect 13745 25427 13757 25461
rect 13699 25393 13757 25427
rect 13699 25359 13711 25393
rect 13745 25359 13757 25393
rect 13699 25325 13757 25359
rect 13699 25291 13711 25325
rect 13745 25291 13757 25325
rect 13699 25257 13757 25291
rect 13699 25223 13711 25257
rect 13745 25223 13757 25257
rect 13699 25189 13757 25223
rect 13699 25155 13711 25189
rect 13745 25155 13757 25189
rect 13699 25121 13757 25155
rect 13699 25087 13711 25121
rect 13745 25087 13757 25121
rect 13699 25053 13757 25087
rect 13699 25019 13711 25053
rect 13745 25019 13757 25053
rect 13699 24985 13757 25019
rect 13699 24951 13711 24985
rect 13745 24951 13757 24985
rect 13699 24917 13757 24951
rect 13699 24883 13711 24917
rect 13745 24883 13757 24917
rect 13699 24867 13757 24883
rect 14157 26141 14215 26157
rect 14157 26107 14169 26141
rect 14203 26107 14215 26141
rect 14157 26073 14215 26107
rect 14157 26039 14169 26073
rect 14203 26039 14215 26073
rect 14157 26005 14215 26039
rect 14157 25971 14169 26005
rect 14203 25971 14215 26005
rect 14157 25937 14215 25971
rect 14157 25903 14169 25937
rect 14203 25903 14215 25937
rect 14157 25869 14215 25903
rect 14157 25835 14169 25869
rect 14203 25835 14215 25869
rect 14157 25801 14215 25835
rect 14157 25767 14169 25801
rect 14203 25767 14215 25801
rect 14157 25733 14215 25767
rect 14157 25699 14169 25733
rect 14203 25699 14215 25733
rect 14157 25665 14215 25699
rect 14157 25631 14169 25665
rect 14203 25631 14215 25665
rect 14157 25597 14215 25631
rect 14157 25563 14169 25597
rect 14203 25563 14215 25597
rect 14157 25529 14215 25563
rect 14157 25495 14169 25529
rect 14203 25495 14215 25529
rect 14157 25461 14215 25495
rect 14157 25427 14169 25461
rect 14203 25427 14215 25461
rect 14157 25393 14215 25427
rect 14157 25359 14169 25393
rect 14203 25359 14215 25393
rect 14157 25325 14215 25359
rect 14157 25291 14169 25325
rect 14203 25291 14215 25325
rect 14157 25257 14215 25291
rect 14157 25223 14169 25257
rect 14203 25223 14215 25257
rect 14157 25189 14215 25223
rect 14157 25155 14169 25189
rect 14203 25155 14215 25189
rect 14157 25121 14215 25155
rect 14157 25087 14169 25121
rect 14203 25087 14215 25121
rect 14157 25053 14215 25087
rect 14157 25019 14169 25053
rect 14203 25019 14215 25053
rect 14157 24985 14215 25019
rect 14157 24951 14169 24985
rect 14203 24951 14215 24985
rect 14157 24917 14215 24951
rect 14157 24883 14169 24917
rect 14203 24883 14215 24917
rect 14157 24867 14215 24883
rect 14615 26141 14673 26157
rect 14615 26107 14627 26141
rect 14661 26107 14673 26141
rect 14615 26073 14673 26107
rect 14615 26039 14627 26073
rect 14661 26039 14673 26073
rect 14615 26005 14673 26039
rect 14615 25971 14627 26005
rect 14661 25971 14673 26005
rect 14615 25937 14673 25971
rect 14615 25903 14627 25937
rect 14661 25903 14673 25937
rect 14615 25869 14673 25903
rect 14615 25835 14627 25869
rect 14661 25835 14673 25869
rect 14615 25801 14673 25835
rect 14615 25767 14627 25801
rect 14661 25767 14673 25801
rect 14615 25733 14673 25767
rect 14615 25699 14627 25733
rect 14661 25699 14673 25733
rect 14615 25665 14673 25699
rect 14615 25631 14627 25665
rect 14661 25631 14673 25665
rect 14615 25597 14673 25631
rect 14615 25563 14627 25597
rect 14661 25563 14673 25597
rect 14615 25529 14673 25563
rect 14615 25495 14627 25529
rect 14661 25495 14673 25529
rect 14615 25461 14673 25495
rect 14615 25427 14627 25461
rect 14661 25427 14673 25461
rect 14615 25393 14673 25427
rect 14615 25359 14627 25393
rect 14661 25359 14673 25393
rect 14615 25325 14673 25359
rect 14615 25291 14627 25325
rect 14661 25291 14673 25325
rect 14615 25257 14673 25291
rect 14615 25223 14627 25257
rect 14661 25223 14673 25257
rect 14615 25189 14673 25223
rect 14615 25155 14627 25189
rect 14661 25155 14673 25189
rect 14615 25121 14673 25155
rect 14615 25087 14627 25121
rect 14661 25087 14673 25121
rect 14615 25053 14673 25087
rect 14615 25019 14627 25053
rect 14661 25019 14673 25053
rect 14615 24985 14673 25019
rect 14615 24951 14627 24985
rect 14661 24951 14673 24985
rect 14615 24917 14673 24951
rect 14615 24883 14627 24917
rect 14661 24883 14673 24917
rect 14615 24867 14673 24883
rect 15073 26141 15131 26157
rect 15073 26107 15085 26141
rect 15119 26107 15131 26141
rect 15073 26073 15131 26107
rect 15073 26039 15085 26073
rect 15119 26039 15131 26073
rect 15073 26005 15131 26039
rect 15073 25971 15085 26005
rect 15119 25971 15131 26005
rect 15073 25937 15131 25971
rect 15073 25903 15085 25937
rect 15119 25903 15131 25937
rect 15073 25869 15131 25903
rect 15073 25835 15085 25869
rect 15119 25835 15131 25869
rect 15073 25801 15131 25835
rect 15073 25767 15085 25801
rect 15119 25767 15131 25801
rect 15073 25733 15131 25767
rect 15073 25699 15085 25733
rect 15119 25699 15131 25733
rect 15073 25665 15131 25699
rect 15073 25631 15085 25665
rect 15119 25631 15131 25665
rect 15073 25597 15131 25631
rect 15073 25563 15085 25597
rect 15119 25563 15131 25597
rect 15073 25529 15131 25563
rect 15073 25495 15085 25529
rect 15119 25495 15131 25529
rect 15073 25461 15131 25495
rect 15073 25427 15085 25461
rect 15119 25427 15131 25461
rect 15073 25393 15131 25427
rect 15073 25359 15085 25393
rect 15119 25359 15131 25393
rect 15073 25325 15131 25359
rect 15073 25291 15085 25325
rect 15119 25291 15131 25325
rect 15073 25257 15131 25291
rect 15073 25223 15085 25257
rect 15119 25223 15131 25257
rect 15073 25189 15131 25223
rect 15073 25155 15085 25189
rect 15119 25155 15131 25189
rect 15073 25121 15131 25155
rect 15073 25087 15085 25121
rect 15119 25087 15131 25121
rect 15073 25053 15131 25087
rect 15073 25019 15085 25053
rect 15119 25019 15131 25053
rect 15073 24985 15131 25019
rect 15073 24951 15085 24985
rect 15119 24951 15131 24985
rect 15073 24917 15131 24951
rect 15073 24883 15085 24917
rect 15119 24883 15131 24917
rect 28590 25740 29270 25792
rect 28590 25706 28644 25740
rect 28678 25706 28734 25740
rect 28768 25706 28824 25740
rect 28858 25706 28914 25740
rect 28948 25706 29004 25740
rect 29038 25706 29094 25740
rect 29128 25706 29184 25740
rect 29218 25706 29270 25740
rect 28590 25650 29270 25706
rect 28590 25616 28644 25650
rect 28678 25616 28734 25650
rect 28768 25616 28824 25650
rect 28858 25616 28914 25650
rect 28948 25616 29004 25650
rect 29038 25616 29094 25650
rect 29128 25616 29184 25650
rect 29218 25616 29270 25650
rect 28590 25560 29270 25616
rect 28590 25526 28644 25560
rect 28678 25526 28734 25560
rect 28768 25526 28824 25560
rect 28858 25526 28914 25560
rect 28948 25526 29004 25560
rect 29038 25526 29094 25560
rect 29128 25526 29184 25560
rect 29218 25526 29270 25560
rect 28590 25470 29270 25526
rect 28590 25436 28644 25470
rect 28678 25436 28734 25470
rect 28768 25436 28824 25470
rect 28858 25436 28914 25470
rect 28948 25436 29004 25470
rect 29038 25436 29094 25470
rect 29128 25436 29184 25470
rect 29218 25436 29270 25470
rect 28590 25380 29270 25436
rect 28590 25346 28644 25380
rect 28678 25346 28734 25380
rect 28768 25346 28824 25380
rect 28858 25346 28914 25380
rect 28948 25346 29004 25380
rect 29038 25346 29094 25380
rect 29128 25346 29184 25380
rect 29218 25346 29270 25380
rect 28590 25290 29270 25346
rect 28590 25256 28644 25290
rect 28678 25256 28734 25290
rect 28768 25256 28824 25290
rect 28858 25256 28914 25290
rect 28948 25256 29004 25290
rect 29038 25256 29094 25290
rect 29128 25256 29184 25290
rect 29218 25256 29270 25290
rect 28590 25200 29270 25256
rect 28590 25166 28644 25200
rect 28678 25166 28734 25200
rect 28768 25166 28824 25200
rect 28858 25166 28914 25200
rect 28948 25166 29004 25200
rect 29038 25166 29094 25200
rect 29128 25166 29184 25200
rect 29218 25166 29270 25200
rect 28590 25112 29270 25166
rect 29930 25740 30610 25792
rect 29930 25706 29984 25740
rect 30018 25706 30074 25740
rect 30108 25706 30164 25740
rect 30198 25706 30254 25740
rect 30288 25706 30344 25740
rect 30378 25706 30434 25740
rect 30468 25706 30524 25740
rect 30558 25706 30610 25740
rect 29930 25650 30610 25706
rect 29930 25616 29984 25650
rect 30018 25616 30074 25650
rect 30108 25616 30164 25650
rect 30198 25616 30254 25650
rect 30288 25616 30344 25650
rect 30378 25616 30434 25650
rect 30468 25616 30524 25650
rect 30558 25616 30610 25650
rect 29930 25560 30610 25616
rect 29930 25526 29984 25560
rect 30018 25526 30074 25560
rect 30108 25526 30164 25560
rect 30198 25526 30254 25560
rect 30288 25526 30344 25560
rect 30378 25526 30434 25560
rect 30468 25526 30524 25560
rect 30558 25526 30610 25560
rect 29930 25470 30610 25526
rect 29930 25436 29984 25470
rect 30018 25436 30074 25470
rect 30108 25436 30164 25470
rect 30198 25436 30254 25470
rect 30288 25436 30344 25470
rect 30378 25436 30434 25470
rect 30468 25436 30524 25470
rect 30558 25436 30610 25470
rect 29930 25380 30610 25436
rect 29930 25346 29984 25380
rect 30018 25346 30074 25380
rect 30108 25346 30164 25380
rect 30198 25346 30254 25380
rect 30288 25346 30344 25380
rect 30378 25346 30434 25380
rect 30468 25346 30524 25380
rect 30558 25346 30610 25380
rect 29930 25290 30610 25346
rect 29930 25256 29984 25290
rect 30018 25256 30074 25290
rect 30108 25256 30164 25290
rect 30198 25256 30254 25290
rect 30288 25256 30344 25290
rect 30378 25256 30434 25290
rect 30468 25256 30524 25290
rect 30558 25256 30610 25290
rect 29930 25200 30610 25256
rect 29930 25166 29984 25200
rect 30018 25166 30074 25200
rect 30108 25166 30164 25200
rect 30198 25166 30254 25200
rect 30288 25166 30344 25200
rect 30378 25166 30434 25200
rect 30468 25166 30524 25200
rect 30558 25166 30610 25200
rect 29930 25112 30610 25166
rect 31270 25740 31950 25792
rect 31270 25706 31324 25740
rect 31358 25706 31414 25740
rect 31448 25706 31504 25740
rect 31538 25706 31594 25740
rect 31628 25706 31684 25740
rect 31718 25706 31774 25740
rect 31808 25706 31864 25740
rect 31898 25706 31950 25740
rect 31270 25650 31950 25706
rect 31270 25616 31324 25650
rect 31358 25616 31414 25650
rect 31448 25616 31504 25650
rect 31538 25616 31594 25650
rect 31628 25616 31684 25650
rect 31718 25616 31774 25650
rect 31808 25616 31864 25650
rect 31898 25616 31950 25650
rect 31270 25560 31950 25616
rect 31270 25526 31324 25560
rect 31358 25526 31414 25560
rect 31448 25526 31504 25560
rect 31538 25526 31594 25560
rect 31628 25526 31684 25560
rect 31718 25526 31774 25560
rect 31808 25526 31864 25560
rect 31898 25526 31950 25560
rect 31270 25470 31950 25526
rect 31270 25436 31324 25470
rect 31358 25436 31414 25470
rect 31448 25436 31504 25470
rect 31538 25436 31594 25470
rect 31628 25436 31684 25470
rect 31718 25436 31774 25470
rect 31808 25436 31864 25470
rect 31898 25436 31950 25470
rect 31270 25380 31950 25436
rect 31270 25346 31324 25380
rect 31358 25346 31414 25380
rect 31448 25346 31504 25380
rect 31538 25346 31594 25380
rect 31628 25346 31684 25380
rect 31718 25346 31774 25380
rect 31808 25346 31864 25380
rect 31898 25346 31950 25380
rect 31270 25290 31950 25346
rect 31270 25256 31324 25290
rect 31358 25256 31414 25290
rect 31448 25256 31504 25290
rect 31538 25256 31594 25290
rect 31628 25256 31684 25290
rect 31718 25256 31774 25290
rect 31808 25256 31864 25290
rect 31898 25256 31950 25290
rect 31270 25200 31950 25256
rect 31270 25166 31324 25200
rect 31358 25166 31414 25200
rect 31448 25166 31504 25200
rect 31538 25166 31594 25200
rect 31628 25166 31684 25200
rect 31718 25166 31774 25200
rect 31808 25166 31864 25200
rect 31898 25166 31950 25200
rect 31270 25112 31950 25166
rect 32610 25740 33290 25792
rect 32610 25706 32664 25740
rect 32698 25706 32754 25740
rect 32788 25706 32844 25740
rect 32878 25706 32934 25740
rect 32968 25706 33024 25740
rect 33058 25706 33114 25740
rect 33148 25706 33204 25740
rect 33238 25706 33290 25740
rect 32610 25650 33290 25706
rect 32610 25616 32664 25650
rect 32698 25616 32754 25650
rect 32788 25616 32844 25650
rect 32878 25616 32934 25650
rect 32968 25616 33024 25650
rect 33058 25616 33114 25650
rect 33148 25616 33204 25650
rect 33238 25616 33290 25650
rect 32610 25560 33290 25616
rect 32610 25526 32664 25560
rect 32698 25526 32754 25560
rect 32788 25526 32844 25560
rect 32878 25526 32934 25560
rect 32968 25526 33024 25560
rect 33058 25526 33114 25560
rect 33148 25526 33204 25560
rect 33238 25526 33290 25560
rect 32610 25470 33290 25526
rect 32610 25436 32664 25470
rect 32698 25436 32754 25470
rect 32788 25436 32844 25470
rect 32878 25436 32934 25470
rect 32968 25436 33024 25470
rect 33058 25436 33114 25470
rect 33148 25436 33204 25470
rect 33238 25436 33290 25470
rect 32610 25380 33290 25436
rect 32610 25346 32664 25380
rect 32698 25346 32754 25380
rect 32788 25346 32844 25380
rect 32878 25346 32934 25380
rect 32968 25346 33024 25380
rect 33058 25346 33114 25380
rect 33148 25346 33204 25380
rect 33238 25346 33290 25380
rect 32610 25290 33290 25346
rect 32610 25256 32664 25290
rect 32698 25256 32754 25290
rect 32788 25256 32844 25290
rect 32878 25256 32934 25290
rect 32968 25256 33024 25290
rect 33058 25256 33114 25290
rect 33148 25256 33204 25290
rect 33238 25256 33290 25290
rect 32610 25200 33290 25256
rect 32610 25166 32664 25200
rect 32698 25166 32754 25200
rect 32788 25166 32844 25200
rect 32878 25166 32934 25200
rect 32968 25166 33024 25200
rect 33058 25166 33114 25200
rect 33148 25166 33204 25200
rect 33238 25166 33290 25200
rect 32610 25112 33290 25166
rect 33950 25740 34630 25792
rect 33950 25706 34004 25740
rect 34038 25706 34094 25740
rect 34128 25706 34184 25740
rect 34218 25706 34274 25740
rect 34308 25706 34364 25740
rect 34398 25706 34454 25740
rect 34488 25706 34544 25740
rect 34578 25706 34630 25740
rect 33950 25650 34630 25706
rect 33950 25616 34004 25650
rect 34038 25616 34094 25650
rect 34128 25616 34184 25650
rect 34218 25616 34274 25650
rect 34308 25616 34364 25650
rect 34398 25616 34454 25650
rect 34488 25616 34544 25650
rect 34578 25616 34630 25650
rect 33950 25560 34630 25616
rect 33950 25526 34004 25560
rect 34038 25526 34094 25560
rect 34128 25526 34184 25560
rect 34218 25526 34274 25560
rect 34308 25526 34364 25560
rect 34398 25526 34454 25560
rect 34488 25526 34544 25560
rect 34578 25526 34630 25560
rect 33950 25470 34630 25526
rect 33950 25436 34004 25470
rect 34038 25436 34094 25470
rect 34128 25436 34184 25470
rect 34218 25436 34274 25470
rect 34308 25436 34364 25470
rect 34398 25436 34454 25470
rect 34488 25436 34544 25470
rect 34578 25436 34630 25470
rect 33950 25380 34630 25436
rect 33950 25346 34004 25380
rect 34038 25346 34094 25380
rect 34128 25346 34184 25380
rect 34218 25346 34274 25380
rect 34308 25346 34364 25380
rect 34398 25346 34454 25380
rect 34488 25346 34544 25380
rect 34578 25346 34630 25380
rect 33950 25290 34630 25346
rect 33950 25256 34004 25290
rect 34038 25256 34094 25290
rect 34128 25256 34184 25290
rect 34218 25256 34274 25290
rect 34308 25256 34364 25290
rect 34398 25256 34454 25290
rect 34488 25256 34544 25290
rect 34578 25256 34630 25290
rect 33950 25200 34630 25256
rect 33950 25166 34004 25200
rect 34038 25166 34094 25200
rect 34128 25166 34184 25200
rect 34218 25166 34274 25200
rect 34308 25166 34364 25200
rect 34398 25166 34454 25200
rect 34488 25166 34544 25200
rect 34578 25166 34630 25200
rect 33950 25112 34630 25166
rect 35290 25740 35970 25792
rect 35290 25706 35344 25740
rect 35378 25706 35434 25740
rect 35468 25706 35524 25740
rect 35558 25706 35614 25740
rect 35648 25706 35704 25740
rect 35738 25706 35794 25740
rect 35828 25706 35884 25740
rect 35918 25706 35970 25740
rect 35290 25650 35970 25706
rect 35290 25616 35344 25650
rect 35378 25616 35434 25650
rect 35468 25616 35524 25650
rect 35558 25616 35614 25650
rect 35648 25616 35704 25650
rect 35738 25616 35794 25650
rect 35828 25616 35884 25650
rect 35918 25616 35970 25650
rect 35290 25560 35970 25616
rect 35290 25526 35344 25560
rect 35378 25526 35434 25560
rect 35468 25526 35524 25560
rect 35558 25526 35614 25560
rect 35648 25526 35704 25560
rect 35738 25526 35794 25560
rect 35828 25526 35884 25560
rect 35918 25526 35970 25560
rect 35290 25470 35970 25526
rect 35290 25436 35344 25470
rect 35378 25436 35434 25470
rect 35468 25436 35524 25470
rect 35558 25436 35614 25470
rect 35648 25436 35704 25470
rect 35738 25436 35794 25470
rect 35828 25436 35884 25470
rect 35918 25436 35970 25470
rect 35290 25380 35970 25436
rect 35290 25346 35344 25380
rect 35378 25346 35434 25380
rect 35468 25346 35524 25380
rect 35558 25346 35614 25380
rect 35648 25346 35704 25380
rect 35738 25346 35794 25380
rect 35828 25346 35884 25380
rect 35918 25346 35970 25380
rect 35290 25290 35970 25346
rect 35290 25256 35344 25290
rect 35378 25256 35434 25290
rect 35468 25256 35524 25290
rect 35558 25256 35614 25290
rect 35648 25256 35704 25290
rect 35738 25256 35794 25290
rect 35828 25256 35884 25290
rect 35918 25256 35970 25290
rect 35290 25200 35970 25256
rect 35290 25166 35344 25200
rect 35378 25166 35434 25200
rect 35468 25166 35524 25200
rect 35558 25166 35614 25200
rect 35648 25166 35704 25200
rect 35738 25166 35794 25200
rect 35828 25166 35884 25200
rect 35918 25166 35970 25200
rect 35290 25112 35970 25166
rect 36630 25740 37310 25792
rect 36630 25706 36684 25740
rect 36718 25706 36774 25740
rect 36808 25706 36864 25740
rect 36898 25706 36954 25740
rect 36988 25706 37044 25740
rect 37078 25706 37134 25740
rect 37168 25706 37224 25740
rect 37258 25706 37310 25740
rect 36630 25650 37310 25706
rect 36630 25616 36684 25650
rect 36718 25616 36774 25650
rect 36808 25616 36864 25650
rect 36898 25616 36954 25650
rect 36988 25616 37044 25650
rect 37078 25616 37134 25650
rect 37168 25616 37224 25650
rect 37258 25616 37310 25650
rect 36630 25560 37310 25616
rect 36630 25526 36684 25560
rect 36718 25526 36774 25560
rect 36808 25526 36864 25560
rect 36898 25526 36954 25560
rect 36988 25526 37044 25560
rect 37078 25526 37134 25560
rect 37168 25526 37224 25560
rect 37258 25526 37310 25560
rect 36630 25470 37310 25526
rect 36630 25436 36684 25470
rect 36718 25436 36774 25470
rect 36808 25436 36864 25470
rect 36898 25436 36954 25470
rect 36988 25436 37044 25470
rect 37078 25436 37134 25470
rect 37168 25436 37224 25470
rect 37258 25436 37310 25470
rect 36630 25380 37310 25436
rect 36630 25346 36684 25380
rect 36718 25346 36774 25380
rect 36808 25346 36864 25380
rect 36898 25346 36954 25380
rect 36988 25346 37044 25380
rect 37078 25346 37134 25380
rect 37168 25346 37224 25380
rect 37258 25346 37310 25380
rect 36630 25290 37310 25346
rect 36630 25256 36684 25290
rect 36718 25256 36774 25290
rect 36808 25256 36864 25290
rect 36898 25256 36954 25290
rect 36988 25256 37044 25290
rect 37078 25256 37134 25290
rect 37168 25256 37224 25290
rect 37258 25256 37310 25290
rect 36630 25200 37310 25256
rect 36630 25166 36684 25200
rect 36718 25166 36774 25200
rect 36808 25166 36864 25200
rect 36898 25166 36954 25200
rect 36988 25166 37044 25200
rect 37078 25166 37134 25200
rect 37168 25166 37224 25200
rect 37258 25166 37310 25200
rect 36630 25112 37310 25166
rect 37970 25740 38650 25792
rect 37970 25706 38024 25740
rect 38058 25706 38114 25740
rect 38148 25706 38204 25740
rect 38238 25706 38294 25740
rect 38328 25706 38384 25740
rect 38418 25706 38474 25740
rect 38508 25706 38564 25740
rect 38598 25706 38650 25740
rect 37970 25650 38650 25706
rect 37970 25616 38024 25650
rect 38058 25616 38114 25650
rect 38148 25616 38204 25650
rect 38238 25616 38294 25650
rect 38328 25616 38384 25650
rect 38418 25616 38474 25650
rect 38508 25616 38564 25650
rect 38598 25616 38650 25650
rect 37970 25560 38650 25616
rect 37970 25526 38024 25560
rect 38058 25526 38114 25560
rect 38148 25526 38204 25560
rect 38238 25526 38294 25560
rect 38328 25526 38384 25560
rect 38418 25526 38474 25560
rect 38508 25526 38564 25560
rect 38598 25526 38650 25560
rect 37970 25470 38650 25526
rect 37970 25436 38024 25470
rect 38058 25436 38114 25470
rect 38148 25436 38204 25470
rect 38238 25436 38294 25470
rect 38328 25436 38384 25470
rect 38418 25436 38474 25470
rect 38508 25436 38564 25470
rect 38598 25436 38650 25470
rect 37970 25380 38650 25436
rect 37970 25346 38024 25380
rect 38058 25346 38114 25380
rect 38148 25346 38204 25380
rect 38238 25346 38294 25380
rect 38328 25346 38384 25380
rect 38418 25346 38474 25380
rect 38508 25346 38564 25380
rect 38598 25346 38650 25380
rect 37970 25290 38650 25346
rect 37970 25256 38024 25290
rect 38058 25256 38114 25290
rect 38148 25256 38204 25290
rect 38238 25256 38294 25290
rect 38328 25256 38384 25290
rect 38418 25256 38474 25290
rect 38508 25256 38564 25290
rect 38598 25256 38650 25290
rect 37970 25200 38650 25256
rect 37970 25166 38024 25200
rect 38058 25166 38114 25200
rect 38148 25166 38204 25200
rect 38238 25166 38294 25200
rect 38328 25166 38384 25200
rect 38418 25166 38474 25200
rect 38508 25166 38564 25200
rect 38598 25166 38650 25200
rect 37970 25112 38650 25166
rect 15073 24867 15131 24883
rect 7715 22381 7773 22397
rect 7715 22347 7727 22381
rect 7761 22347 7773 22381
rect 7715 22313 7773 22347
rect 7715 22279 7727 22313
rect 7761 22279 7773 22313
rect 7715 22245 7773 22279
rect 7715 22211 7727 22245
rect 7761 22211 7773 22245
rect 7715 22177 7773 22211
rect 7715 22143 7727 22177
rect 7761 22143 7773 22177
rect 7715 22109 7773 22143
rect 7715 22075 7727 22109
rect 7761 22075 7773 22109
rect 7715 22041 7773 22075
rect 7715 22007 7727 22041
rect 7761 22007 7773 22041
rect 7715 21973 7773 22007
rect 7715 21939 7727 21973
rect 7761 21939 7773 21973
rect 7715 21905 7773 21939
rect 7715 21871 7727 21905
rect 7761 21871 7773 21905
rect 7715 21837 7773 21871
rect 7715 21803 7727 21837
rect 7761 21803 7773 21837
rect 7715 21769 7773 21803
rect 7715 21735 7727 21769
rect 7761 21735 7773 21769
rect 7715 21701 7773 21735
rect 7715 21667 7727 21701
rect 7761 21667 7773 21701
rect 7715 21633 7773 21667
rect 7715 21599 7727 21633
rect 7761 21599 7773 21633
rect 7715 21565 7773 21599
rect 7715 21531 7727 21565
rect 7761 21531 7773 21565
rect 7715 21497 7773 21531
rect 7715 21463 7727 21497
rect 7761 21463 7773 21497
rect 7715 21429 7773 21463
rect 7715 21395 7727 21429
rect 7761 21395 7773 21429
rect 7715 21361 7773 21395
rect 7715 21327 7727 21361
rect 7761 21327 7773 21361
rect 7715 21293 7773 21327
rect 7715 21259 7727 21293
rect 7761 21259 7773 21293
rect 7715 21225 7773 21259
rect 7715 21191 7727 21225
rect 7761 21191 7773 21225
rect 7715 21157 7773 21191
rect 7715 21123 7727 21157
rect 7761 21123 7773 21157
rect 7715 21107 7773 21123
rect 8173 22381 8231 22397
rect 8173 22347 8185 22381
rect 8219 22347 8231 22381
rect 8173 22313 8231 22347
rect 8173 22279 8185 22313
rect 8219 22279 8231 22313
rect 8173 22245 8231 22279
rect 8173 22211 8185 22245
rect 8219 22211 8231 22245
rect 8173 22177 8231 22211
rect 8173 22143 8185 22177
rect 8219 22143 8231 22177
rect 8173 22109 8231 22143
rect 8173 22075 8185 22109
rect 8219 22075 8231 22109
rect 8173 22041 8231 22075
rect 8173 22007 8185 22041
rect 8219 22007 8231 22041
rect 8173 21973 8231 22007
rect 8173 21939 8185 21973
rect 8219 21939 8231 21973
rect 8173 21905 8231 21939
rect 8173 21871 8185 21905
rect 8219 21871 8231 21905
rect 8173 21837 8231 21871
rect 8173 21803 8185 21837
rect 8219 21803 8231 21837
rect 8173 21769 8231 21803
rect 8173 21735 8185 21769
rect 8219 21735 8231 21769
rect 8173 21701 8231 21735
rect 8173 21667 8185 21701
rect 8219 21667 8231 21701
rect 8173 21633 8231 21667
rect 8173 21599 8185 21633
rect 8219 21599 8231 21633
rect 8173 21565 8231 21599
rect 8173 21531 8185 21565
rect 8219 21531 8231 21565
rect 8173 21497 8231 21531
rect 8173 21463 8185 21497
rect 8219 21463 8231 21497
rect 8173 21429 8231 21463
rect 8173 21395 8185 21429
rect 8219 21395 8231 21429
rect 8173 21361 8231 21395
rect 8173 21327 8185 21361
rect 8219 21327 8231 21361
rect 8173 21293 8231 21327
rect 8173 21259 8185 21293
rect 8219 21259 8231 21293
rect 8173 21225 8231 21259
rect 8173 21191 8185 21225
rect 8219 21191 8231 21225
rect 8173 21157 8231 21191
rect 8173 21123 8185 21157
rect 8219 21123 8231 21157
rect 8173 21107 8231 21123
rect 8631 22381 8689 22397
rect 8631 22347 8643 22381
rect 8677 22347 8689 22381
rect 8631 22313 8689 22347
rect 8631 22279 8643 22313
rect 8677 22279 8689 22313
rect 8631 22245 8689 22279
rect 8631 22211 8643 22245
rect 8677 22211 8689 22245
rect 8631 22177 8689 22211
rect 8631 22143 8643 22177
rect 8677 22143 8689 22177
rect 8631 22109 8689 22143
rect 8631 22075 8643 22109
rect 8677 22075 8689 22109
rect 8631 22041 8689 22075
rect 8631 22007 8643 22041
rect 8677 22007 8689 22041
rect 8631 21973 8689 22007
rect 8631 21939 8643 21973
rect 8677 21939 8689 21973
rect 8631 21905 8689 21939
rect 8631 21871 8643 21905
rect 8677 21871 8689 21905
rect 8631 21837 8689 21871
rect 8631 21803 8643 21837
rect 8677 21803 8689 21837
rect 8631 21769 8689 21803
rect 8631 21735 8643 21769
rect 8677 21735 8689 21769
rect 8631 21701 8689 21735
rect 8631 21667 8643 21701
rect 8677 21667 8689 21701
rect 8631 21633 8689 21667
rect 8631 21599 8643 21633
rect 8677 21599 8689 21633
rect 8631 21565 8689 21599
rect 8631 21531 8643 21565
rect 8677 21531 8689 21565
rect 8631 21497 8689 21531
rect 8631 21463 8643 21497
rect 8677 21463 8689 21497
rect 8631 21429 8689 21463
rect 8631 21395 8643 21429
rect 8677 21395 8689 21429
rect 8631 21361 8689 21395
rect 8631 21327 8643 21361
rect 8677 21327 8689 21361
rect 8631 21293 8689 21327
rect 8631 21259 8643 21293
rect 8677 21259 8689 21293
rect 8631 21225 8689 21259
rect 8631 21191 8643 21225
rect 8677 21191 8689 21225
rect 8631 21157 8689 21191
rect 8631 21123 8643 21157
rect 8677 21123 8689 21157
rect 8631 21107 8689 21123
rect 9089 22381 9147 22397
rect 9089 22347 9101 22381
rect 9135 22347 9147 22381
rect 9089 22313 9147 22347
rect 9089 22279 9101 22313
rect 9135 22279 9147 22313
rect 9089 22245 9147 22279
rect 9089 22211 9101 22245
rect 9135 22211 9147 22245
rect 9089 22177 9147 22211
rect 9089 22143 9101 22177
rect 9135 22143 9147 22177
rect 9089 22109 9147 22143
rect 9089 22075 9101 22109
rect 9135 22075 9147 22109
rect 9089 22041 9147 22075
rect 9089 22007 9101 22041
rect 9135 22007 9147 22041
rect 9089 21973 9147 22007
rect 9089 21939 9101 21973
rect 9135 21939 9147 21973
rect 9089 21905 9147 21939
rect 9089 21871 9101 21905
rect 9135 21871 9147 21905
rect 9089 21837 9147 21871
rect 9089 21803 9101 21837
rect 9135 21803 9147 21837
rect 9089 21769 9147 21803
rect 9089 21735 9101 21769
rect 9135 21735 9147 21769
rect 9089 21701 9147 21735
rect 9089 21667 9101 21701
rect 9135 21667 9147 21701
rect 9089 21633 9147 21667
rect 9089 21599 9101 21633
rect 9135 21599 9147 21633
rect 9089 21565 9147 21599
rect 9089 21531 9101 21565
rect 9135 21531 9147 21565
rect 9089 21497 9147 21531
rect 9089 21463 9101 21497
rect 9135 21463 9147 21497
rect 9089 21429 9147 21463
rect 9089 21395 9101 21429
rect 9135 21395 9147 21429
rect 9089 21361 9147 21395
rect 9089 21327 9101 21361
rect 9135 21327 9147 21361
rect 9089 21293 9147 21327
rect 9089 21259 9101 21293
rect 9135 21259 9147 21293
rect 9089 21225 9147 21259
rect 9089 21191 9101 21225
rect 9135 21191 9147 21225
rect 9089 21157 9147 21191
rect 9089 21123 9101 21157
rect 9135 21123 9147 21157
rect 9089 21107 9147 21123
rect 9547 22381 9605 22397
rect 9547 22347 9559 22381
rect 9593 22347 9605 22381
rect 9547 22313 9605 22347
rect 9547 22279 9559 22313
rect 9593 22279 9605 22313
rect 9547 22245 9605 22279
rect 9547 22211 9559 22245
rect 9593 22211 9605 22245
rect 9547 22177 9605 22211
rect 9547 22143 9559 22177
rect 9593 22143 9605 22177
rect 9547 22109 9605 22143
rect 9547 22075 9559 22109
rect 9593 22075 9605 22109
rect 9547 22041 9605 22075
rect 9547 22007 9559 22041
rect 9593 22007 9605 22041
rect 9547 21973 9605 22007
rect 9547 21939 9559 21973
rect 9593 21939 9605 21973
rect 9547 21905 9605 21939
rect 9547 21871 9559 21905
rect 9593 21871 9605 21905
rect 9547 21837 9605 21871
rect 9547 21803 9559 21837
rect 9593 21803 9605 21837
rect 9547 21769 9605 21803
rect 9547 21735 9559 21769
rect 9593 21735 9605 21769
rect 9547 21701 9605 21735
rect 9547 21667 9559 21701
rect 9593 21667 9605 21701
rect 9547 21633 9605 21667
rect 9547 21599 9559 21633
rect 9593 21599 9605 21633
rect 9547 21565 9605 21599
rect 9547 21531 9559 21565
rect 9593 21531 9605 21565
rect 9547 21497 9605 21531
rect 9547 21463 9559 21497
rect 9593 21463 9605 21497
rect 9547 21429 9605 21463
rect 9547 21395 9559 21429
rect 9593 21395 9605 21429
rect 9547 21361 9605 21395
rect 9547 21327 9559 21361
rect 9593 21327 9605 21361
rect 9547 21293 9605 21327
rect 9547 21259 9559 21293
rect 9593 21259 9605 21293
rect 9547 21225 9605 21259
rect 9547 21191 9559 21225
rect 9593 21191 9605 21225
rect 9547 21157 9605 21191
rect 9547 21123 9559 21157
rect 9593 21123 9605 21157
rect 9547 21107 9605 21123
rect 10005 22381 10063 22397
rect 10005 22347 10017 22381
rect 10051 22347 10063 22381
rect 10005 22313 10063 22347
rect 10005 22279 10017 22313
rect 10051 22279 10063 22313
rect 10005 22245 10063 22279
rect 10005 22211 10017 22245
rect 10051 22211 10063 22245
rect 10005 22177 10063 22211
rect 10005 22143 10017 22177
rect 10051 22143 10063 22177
rect 10005 22109 10063 22143
rect 10005 22075 10017 22109
rect 10051 22075 10063 22109
rect 10005 22041 10063 22075
rect 10005 22007 10017 22041
rect 10051 22007 10063 22041
rect 10005 21973 10063 22007
rect 10005 21939 10017 21973
rect 10051 21939 10063 21973
rect 10005 21905 10063 21939
rect 10005 21871 10017 21905
rect 10051 21871 10063 21905
rect 10005 21837 10063 21871
rect 10005 21803 10017 21837
rect 10051 21803 10063 21837
rect 10005 21769 10063 21803
rect 10005 21735 10017 21769
rect 10051 21735 10063 21769
rect 10005 21701 10063 21735
rect 10005 21667 10017 21701
rect 10051 21667 10063 21701
rect 10005 21633 10063 21667
rect 10005 21599 10017 21633
rect 10051 21599 10063 21633
rect 10005 21565 10063 21599
rect 10005 21531 10017 21565
rect 10051 21531 10063 21565
rect 10005 21497 10063 21531
rect 10005 21463 10017 21497
rect 10051 21463 10063 21497
rect 10005 21429 10063 21463
rect 10005 21395 10017 21429
rect 10051 21395 10063 21429
rect 10005 21361 10063 21395
rect 10005 21327 10017 21361
rect 10051 21327 10063 21361
rect 10005 21293 10063 21327
rect 10005 21259 10017 21293
rect 10051 21259 10063 21293
rect 10005 21225 10063 21259
rect 10005 21191 10017 21225
rect 10051 21191 10063 21225
rect 10005 21157 10063 21191
rect 10005 21123 10017 21157
rect 10051 21123 10063 21157
rect 10005 21107 10063 21123
rect 10463 22381 10521 22397
rect 10463 22347 10475 22381
rect 10509 22347 10521 22381
rect 10463 22313 10521 22347
rect 10463 22279 10475 22313
rect 10509 22279 10521 22313
rect 10463 22245 10521 22279
rect 10463 22211 10475 22245
rect 10509 22211 10521 22245
rect 10463 22177 10521 22211
rect 10463 22143 10475 22177
rect 10509 22143 10521 22177
rect 10463 22109 10521 22143
rect 10463 22075 10475 22109
rect 10509 22075 10521 22109
rect 10463 22041 10521 22075
rect 10463 22007 10475 22041
rect 10509 22007 10521 22041
rect 10463 21973 10521 22007
rect 10463 21939 10475 21973
rect 10509 21939 10521 21973
rect 10463 21905 10521 21939
rect 10463 21871 10475 21905
rect 10509 21871 10521 21905
rect 10463 21837 10521 21871
rect 10463 21803 10475 21837
rect 10509 21803 10521 21837
rect 10463 21769 10521 21803
rect 10463 21735 10475 21769
rect 10509 21735 10521 21769
rect 10463 21701 10521 21735
rect 10463 21667 10475 21701
rect 10509 21667 10521 21701
rect 10463 21633 10521 21667
rect 10463 21599 10475 21633
rect 10509 21599 10521 21633
rect 10463 21565 10521 21599
rect 10463 21531 10475 21565
rect 10509 21531 10521 21565
rect 10463 21497 10521 21531
rect 10463 21463 10475 21497
rect 10509 21463 10521 21497
rect 10463 21429 10521 21463
rect 10463 21395 10475 21429
rect 10509 21395 10521 21429
rect 10463 21361 10521 21395
rect 10463 21327 10475 21361
rect 10509 21327 10521 21361
rect 10463 21293 10521 21327
rect 10463 21259 10475 21293
rect 10509 21259 10521 21293
rect 10463 21225 10521 21259
rect 10463 21191 10475 21225
rect 10509 21191 10521 21225
rect 10463 21157 10521 21191
rect 10463 21123 10475 21157
rect 10509 21123 10521 21157
rect 10463 21107 10521 21123
rect 10921 22381 10979 22397
rect 10921 22347 10933 22381
rect 10967 22347 10979 22381
rect 10921 22313 10979 22347
rect 10921 22279 10933 22313
rect 10967 22279 10979 22313
rect 10921 22245 10979 22279
rect 10921 22211 10933 22245
rect 10967 22211 10979 22245
rect 10921 22177 10979 22211
rect 10921 22143 10933 22177
rect 10967 22143 10979 22177
rect 10921 22109 10979 22143
rect 10921 22075 10933 22109
rect 10967 22075 10979 22109
rect 10921 22041 10979 22075
rect 10921 22007 10933 22041
rect 10967 22007 10979 22041
rect 10921 21973 10979 22007
rect 10921 21939 10933 21973
rect 10967 21939 10979 21973
rect 10921 21905 10979 21939
rect 10921 21871 10933 21905
rect 10967 21871 10979 21905
rect 10921 21837 10979 21871
rect 10921 21803 10933 21837
rect 10967 21803 10979 21837
rect 10921 21769 10979 21803
rect 10921 21735 10933 21769
rect 10967 21735 10979 21769
rect 10921 21701 10979 21735
rect 10921 21667 10933 21701
rect 10967 21667 10979 21701
rect 10921 21633 10979 21667
rect 10921 21599 10933 21633
rect 10967 21599 10979 21633
rect 10921 21565 10979 21599
rect 10921 21531 10933 21565
rect 10967 21531 10979 21565
rect 10921 21497 10979 21531
rect 10921 21463 10933 21497
rect 10967 21463 10979 21497
rect 10921 21429 10979 21463
rect 10921 21395 10933 21429
rect 10967 21395 10979 21429
rect 10921 21361 10979 21395
rect 10921 21327 10933 21361
rect 10967 21327 10979 21361
rect 10921 21293 10979 21327
rect 10921 21259 10933 21293
rect 10967 21259 10979 21293
rect 10921 21225 10979 21259
rect 10921 21191 10933 21225
rect 10967 21191 10979 21225
rect 10921 21157 10979 21191
rect 10921 21123 10933 21157
rect 10967 21123 10979 21157
rect 10921 21107 10979 21123
rect 11379 22381 11437 22397
rect 11379 22347 11391 22381
rect 11425 22347 11437 22381
rect 11379 22313 11437 22347
rect 11379 22279 11391 22313
rect 11425 22279 11437 22313
rect 11379 22245 11437 22279
rect 11379 22211 11391 22245
rect 11425 22211 11437 22245
rect 11379 22177 11437 22211
rect 11379 22143 11391 22177
rect 11425 22143 11437 22177
rect 11379 22109 11437 22143
rect 11379 22075 11391 22109
rect 11425 22075 11437 22109
rect 11379 22041 11437 22075
rect 11379 22007 11391 22041
rect 11425 22007 11437 22041
rect 11379 21973 11437 22007
rect 11379 21939 11391 21973
rect 11425 21939 11437 21973
rect 11379 21905 11437 21939
rect 11379 21871 11391 21905
rect 11425 21871 11437 21905
rect 11379 21837 11437 21871
rect 11379 21803 11391 21837
rect 11425 21803 11437 21837
rect 11379 21769 11437 21803
rect 11379 21735 11391 21769
rect 11425 21735 11437 21769
rect 11379 21701 11437 21735
rect 11379 21667 11391 21701
rect 11425 21667 11437 21701
rect 11379 21633 11437 21667
rect 11379 21599 11391 21633
rect 11425 21599 11437 21633
rect 11379 21565 11437 21599
rect 11379 21531 11391 21565
rect 11425 21531 11437 21565
rect 11379 21497 11437 21531
rect 11379 21463 11391 21497
rect 11425 21463 11437 21497
rect 11379 21429 11437 21463
rect 11379 21395 11391 21429
rect 11425 21395 11437 21429
rect 11379 21361 11437 21395
rect 11379 21327 11391 21361
rect 11425 21327 11437 21361
rect 11379 21293 11437 21327
rect 11379 21259 11391 21293
rect 11425 21259 11437 21293
rect 11379 21225 11437 21259
rect 11379 21191 11391 21225
rect 11425 21191 11437 21225
rect 11379 21157 11437 21191
rect 11379 21123 11391 21157
rect 11425 21123 11437 21157
rect 11379 21107 11437 21123
rect 11837 22381 11895 22397
rect 11837 22347 11849 22381
rect 11883 22347 11895 22381
rect 11837 22313 11895 22347
rect 11837 22279 11849 22313
rect 11883 22279 11895 22313
rect 11837 22245 11895 22279
rect 11837 22211 11849 22245
rect 11883 22211 11895 22245
rect 11837 22177 11895 22211
rect 11837 22143 11849 22177
rect 11883 22143 11895 22177
rect 11837 22109 11895 22143
rect 11837 22075 11849 22109
rect 11883 22075 11895 22109
rect 11837 22041 11895 22075
rect 11837 22007 11849 22041
rect 11883 22007 11895 22041
rect 11837 21973 11895 22007
rect 11837 21939 11849 21973
rect 11883 21939 11895 21973
rect 11837 21905 11895 21939
rect 11837 21871 11849 21905
rect 11883 21871 11895 21905
rect 11837 21837 11895 21871
rect 11837 21803 11849 21837
rect 11883 21803 11895 21837
rect 11837 21769 11895 21803
rect 11837 21735 11849 21769
rect 11883 21735 11895 21769
rect 11837 21701 11895 21735
rect 11837 21667 11849 21701
rect 11883 21667 11895 21701
rect 11837 21633 11895 21667
rect 11837 21599 11849 21633
rect 11883 21599 11895 21633
rect 11837 21565 11895 21599
rect 11837 21531 11849 21565
rect 11883 21531 11895 21565
rect 11837 21497 11895 21531
rect 11837 21463 11849 21497
rect 11883 21463 11895 21497
rect 11837 21429 11895 21463
rect 11837 21395 11849 21429
rect 11883 21395 11895 21429
rect 11837 21361 11895 21395
rect 11837 21327 11849 21361
rect 11883 21327 11895 21361
rect 11837 21293 11895 21327
rect 11837 21259 11849 21293
rect 11883 21259 11895 21293
rect 11837 21225 11895 21259
rect 11837 21191 11849 21225
rect 11883 21191 11895 21225
rect 11837 21157 11895 21191
rect 11837 21123 11849 21157
rect 11883 21123 11895 21157
rect 11837 21107 11895 21123
rect 12295 22381 12353 22397
rect 12295 22347 12307 22381
rect 12341 22347 12353 22381
rect 12295 22313 12353 22347
rect 12295 22279 12307 22313
rect 12341 22279 12353 22313
rect 12295 22245 12353 22279
rect 12295 22211 12307 22245
rect 12341 22211 12353 22245
rect 12295 22177 12353 22211
rect 12295 22143 12307 22177
rect 12341 22143 12353 22177
rect 12295 22109 12353 22143
rect 12295 22075 12307 22109
rect 12341 22075 12353 22109
rect 12295 22041 12353 22075
rect 12295 22007 12307 22041
rect 12341 22007 12353 22041
rect 12295 21973 12353 22007
rect 12295 21939 12307 21973
rect 12341 21939 12353 21973
rect 12295 21905 12353 21939
rect 12295 21871 12307 21905
rect 12341 21871 12353 21905
rect 12295 21837 12353 21871
rect 12295 21803 12307 21837
rect 12341 21803 12353 21837
rect 12295 21769 12353 21803
rect 12295 21735 12307 21769
rect 12341 21735 12353 21769
rect 12295 21701 12353 21735
rect 12295 21667 12307 21701
rect 12341 21667 12353 21701
rect 12295 21633 12353 21667
rect 12295 21599 12307 21633
rect 12341 21599 12353 21633
rect 12295 21565 12353 21599
rect 12295 21531 12307 21565
rect 12341 21531 12353 21565
rect 12295 21497 12353 21531
rect 12295 21463 12307 21497
rect 12341 21463 12353 21497
rect 12295 21429 12353 21463
rect 12295 21395 12307 21429
rect 12341 21395 12353 21429
rect 12295 21361 12353 21395
rect 12295 21327 12307 21361
rect 12341 21327 12353 21361
rect 12295 21293 12353 21327
rect 12295 21259 12307 21293
rect 12341 21259 12353 21293
rect 12295 21225 12353 21259
rect 12295 21191 12307 21225
rect 12341 21191 12353 21225
rect 12295 21157 12353 21191
rect 12295 21123 12307 21157
rect 12341 21123 12353 21157
rect 12295 21107 12353 21123
rect 12753 22381 12811 22397
rect 12753 22347 12765 22381
rect 12799 22347 12811 22381
rect 12753 22313 12811 22347
rect 12753 22279 12765 22313
rect 12799 22279 12811 22313
rect 12753 22245 12811 22279
rect 12753 22211 12765 22245
rect 12799 22211 12811 22245
rect 12753 22177 12811 22211
rect 12753 22143 12765 22177
rect 12799 22143 12811 22177
rect 12753 22109 12811 22143
rect 12753 22075 12765 22109
rect 12799 22075 12811 22109
rect 12753 22041 12811 22075
rect 12753 22007 12765 22041
rect 12799 22007 12811 22041
rect 12753 21973 12811 22007
rect 12753 21939 12765 21973
rect 12799 21939 12811 21973
rect 12753 21905 12811 21939
rect 12753 21871 12765 21905
rect 12799 21871 12811 21905
rect 12753 21837 12811 21871
rect 12753 21803 12765 21837
rect 12799 21803 12811 21837
rect 12753 21769 12811 21803
rect 12753 21735 12765 21769
rect 12799 21735 12811 21769
rect 12753 21701 12811 21735
rect 12753 21667 12765 21701
rect 12799 21667 12811 21701
rect 12753 21633 12811 21667
rect 12753 21599 12765 21633
rect 12799 21599 12811 21633
rect 12753 21565 12811 21599
rect 12753 21531 12765 21565
rect 12799 21531 12811 21565
rect 12753 21497 12811 21531
rect 12753 21463 12765 21497
rect 12799 21463 12811 21497
rect 12753 21429 12811 21463
rect 12753 21395 12765 21429
rect 12799 21395 12811 21429
rect 12753 21361 12811 21395
rect 12753 21327 12765 21361
rect 12799 21327 12811 21361
rect 12753 21293 12811 21327
rect 12753 21259 12765 21293
rect 12799 21259 12811 21293
rect 12753 21225 12811 21259
rect 12753 21191 12765 21225
rect 12799 21191 12811 21225
rect 12753 21157 12811 21191
rect 12753 21123 12765 21157
rect 12799 21123 12811 21157
rect 12753 21107 12811 21123
rect 13211 22381 13269 22397
rect 13211 22347 13223 22381
rect 13257 22347 13269 22381
rect 13211 22313 13269 22347
rect 13211 22279 13223 22313
rect 13257 22279 13269 22313
rect 13211 22245 13269 22279
rect 13211 22211 13223 22245
rect 13257 22211 13269 22245
rect 13211 22177 13269 22211
rect 13211 22143 13223 22177
rect 13257 22143 13269 22177
rect 13211 22109 13269 22143
rect 13211 22075 13223 22109
rect 13257 22075 13269 22109
rect 13211 22041 13269 22075
rect 13211 22007 13223 22041
rect 13257 22007 13269 22041
rect 13211 21973 13269 22007
rect 13211 21939 13223 21973
rect 13257 21939 13269 21973
rect 13211 21905 13269 21939
rect 13211 21871 13223 21905
rect 13257 21871 13269 21905
rect 13211 21837 13269 21871
rect 13211 21803 13223 21837
rect 13257 21803 13269 21837
rect 13211 21769 13269 21803
rect 13211 21735 13223 21769
rect 13257 21735 13269 21769
rect 13211 21701 13269 21735
rect 13211 21667 13223 21701
rect 13257 21667 13269 21701
rect 13211 21633 13269 21667
rect 13211 21599 13223 21633
rect 13257 21599 13269 21633
rect 13211 21565 13269 21599
rect 13211 21531 13223 21565
rect 13257 21531 13269 21565
rect 13211 21497 13269 21531
rect 13211 21463 13223 21497
rect 13257 21463 13269 21497
rect 13211 21429 13269 21463
rect 13211 21395 13223 21429
rect 13257 21395 13269 21429
rect 13211 21361 13269 21395
rect 13211 21327 13223 21361
rect 13257 21327 13269 21361
rect 13211 21293 13269 21327
rect 13211 21259 13223 21293
rect 13257 21259 13269 21293
rect 13211 21225 13269 21259
rect 13211 21191 13223 21225
rect 13257 21191 13269 21225
rect 13211 21157 13269 21191
rect 13211 21123 13223 21157
rect 13257 21123 13269 21157
rect 13211 21107 13269 21123
rect 21338 21980 22018 22032
rect 21338 21946 21392 21980
rect 21426 21946 21482 21980
rect 21516 21946 21572 21980
rect 21606 21946 21662 21980
rect 21696 21946 21752 21980
rect 21786 21946 21842 21980
rect 21876 21946 21932 21980
rect 21966 21946 22018 21980
rect 21338 21890 22018 21946
rect 21338 21856 21392 21890
rect 21426 21856 21482 21890
rect 21516 21856 21572 21890
rect 21606 21856 21662 21890
rect 21696 21856 21752 21890
rect 21786 21856 21842 21890
rect 21876 21856 21932 21890
rect 21966 21856 22018 21890
rect 21338 21800 22018 21856
rect 21338 21766 21392 21800
rect 21426 21766 21482 21800
rect 21516 21766 21572 21800
rect 21606 21766 21662 21800
rect 21696 21766 21752 21800
rect 21786 21766 21842 21800
rect 21876 21766 21932 21800
rect 21966 21766 22018 21800
rect 21338 21710 22018 21766
rect 21338 21676 21392 21710
rect 21426 21676 21482 21710
rect 21516 21676 21572 21710
rect 21606 21676 21662 21710
rect 21696 21676 21752 21710
rect 21786 21676 21842 21710
rect 21876 21676 21932 21710
rect 21966 21676 22018 21710
rect 21338 21620 22018 21676
rect 21338 21586 21392 21620
rect 21426 21586 21482 21620
rect 21516 21586 21572 21620
rect 21606 21586 21662 21620
rect 21696 21586 21752 21620
rect 21786 21586 21842 21620
rect 21876 21586 21932 21620
rect 21966 21586 22018 21620
rect 21338 21530 22018 21586
rect 21338 21496 21392 21530
rect 21426 21496 21482 21530
rect 21516 21496 21572 21530
rect 21606 21496 21662 21530
rect 21696 21496 21752 21530
rect 21786 21496 21842 21530
rect 21876 21496 21932 21530
rect 21966 21496 22018 21530
rect 21338 21440 22018 21496
rect 21338 21406 21392 21440
rect 21426 21406 21482 21440
rect 21516 21406 21572 21440
rect 21606 21406 21662 21440
rect 21696 21406 21752 21440
rect 21786 21406 21842 21440
rect 21876 21406 21932 21440
rect 21966 21406 22018 21440
rect 21338 21352 22018 21406
rect 28590 21980 29270 22032
rect 28590 21946 28644 21980
rect 28678 21946 28734 21980
rect 28768 21946 28824 21980
rect 28858 21946 28914 21980
rect 28948 21946 29004 21980
rect 29038 21946 29094 21980
rect 29128 21946 29184 21980
rect 29218 21946 29270 21980
rect 28590 21890 29270 21946
rect 28590 21856 28644 21890
rect 28678 21856 28734 21890
rect 28768 21856 28824 21890
rect 28858 21856 28914 21890
rect 28948 21856 29004 21890
rect 29038 21856 29094 21890
rect 29128 21856 29184 21890
rect 29218 21856 29270 21890
rect 28590 21800 29270 21856
rect 28590 21766 28644 21800
rect 28678 21766 28734 21800
rect 28768 21766 28824 21800
rect 28858 21766 28914 21800
rect 28948 21766 29004 21800
rect 29038 21766 29094 21800
rect 29128 21766 29184 21800
rect 29218 21766 29270 21800
rect 28590 21710 29270 21766
rect 28590 21676 28644 21710
rect 28678 21676 28734 21710
rect 28768 21676 28824 21710
rect 28858 21676 28914 21710
rect 28948 21676 29004 21710
rect 29038 21676 29094 21710
rect 29128 21676 29184 21710
rect 29218 21676 29270 21710
rect 28590 21620 29270 21676
rect 28590 21586 28644 21620
rect 28678 21586 28734 21620
rect 28768 21586 28824 21620
rect 28858 21586 28914 21620
rect 28948 21586 29004 21620
rect 29038 21586 29094 21620
rect 29128 21586 29184 21620
rect 29218 21586 29270 21620
rect 28590 21530 29270 21586
rect 28590 21496 28644 21530
rect 28678 21496 28734 21530
rect 28768 21496 28824 21530
rect 28858 21496 28914 21530
rect 28948 21496 29004 21530
rect 29038 21496 29094 21530
rect 29128 21496 29184 21530
rect 29218 21496 29270 21530
rect 28590 21440 29270 21496
rect 28590 21406 28644 21440
rect 28678 21406 28734 21440
rect 28768 21406 28824 21440
rect 28858 21406 28914 21440
rect 28948 21406 29004 21440
rect 29038 21406 29094 21440
rect 29128 21406 29184 21440
rect 29218 21406 29270 21440
rect 28590 21352 29270 21406
rect 29930 21980 30610 22032
rect 29930 21946 29984 21980
rect 30018 21946 30074 21980
rect 30108 21946 30164 21980
rect 30198 21946 30254 21980
rect 30288 21946 30344 21980
rect 30378 21946 30434 21980
rect 30468 21946 30524 21980
rect 30558 21946 30610 21980
rect 29930 21890 30610 21946
rect 29930 21856 29984 21890
rect 30018 21856 30074 21890
rect 30108 21856 30164 21890
rect 30198 21856 30254 21890
rect 30288 21856 30344 21890
rect 30378 21856 30434 21890
rect 30468 21856 30524 21890
rect 30558 21856 30610 21890
rect 29930 21800 30610 21856
rect 29930 21766 29984 21800
rect 30018 21766 30074 21800
rect 30108 21766 30164 21800
rect 30198 21766 30254 21800
rect 30288 21766 30344 21800
rect 30378 21766 30434 21800
rect 30468 21766 30524 21800
rect 30558 21766 30610 21800
rect 29930 21710 30610 21766
rect 29930 21676 29984 21710
rect 30018 21676 30074 21710
rect 30108 21676 30164 21710
rect 30198 21676 30254 21710
rect 30288 21676 30344 21710
rect 30378 21676 30434 21710
rect 30468 21676 30524 21710
rect 30558 21676 30610 21710
rect 29930 21620 30610 21676
rect 29930 21586 29984 21620
rect 30018 21586 30074 21620
rect 30108 21586 30164 21620
rect 30198 21586 30254 21620
rect 30288 21586 30344 21620
rect 30378 21586 30434 21620
rect 30468 21586 30524 21620
rect 30558 21586 30610 21620
rect 29930 21530 30610 21586
rect 29930 21496 29984 21530
rect 30018 21496 30074 21530
rect 30108 21496 30164 21530
rect 30198 21496 30254 21530
rect 30288 21496 30344 21530
rect 30378 21496 30434 21530
rect 30468 21496 30524 21530
rect 30558 21496 30610 21530
rect 29930 21440 30610 21496
rect 29930 21406 29984 21440
rect 30018 21406 30074 21440
rect 30108 21406 30164 21440
rect 30198 21406 30254 21440
rect 30288 21406 30344 21440
rect 30378 21406 30434 21440
rect 30468 21406 30524 21440
rect 30558 21406 30610 21440
rect 29930 21352 30610 21406
rect 31270 21980 31950 22032
rect 31270 21946 31324 21980
rect 31358 21946 31414 21980
rect 31448 21946 31504 21980
rect 31538 21946 31594 21980
rect 31628 21946 31684 21980
rect 31718 21946 31774 21980
rect 31808 21946 31864 21980
rect 31898 21946 31950 21980
rect 31270 21890 31950 21946
rect 31270 21856 31324 21890
rect 31358 21856 31414 21890
rect 31448 21856 31504 21890
rect 31538 21856 31594 21890
rect 31628 21856 31684 21890
rect 31718 21856 31774 21890
rect 31808 21856 31864 21890
rect 31898 21856 31950 21890
rect 31270 21800 31950 21856
rect 31270 21766 31324 21800
rect 31358 21766 31414 21800
rect 31448 21766 31504 21800
rect 31538 21766 31594 21800
rect 31628 21766 31684 21800
rect 31718 21766 31774 21800
rect 31808 21766 31864 21800
rect 31898 21766 31950 21800
rect 31270 21710 31950 21766
rect 31270 21676 31324 21710
rect 31358 21676 31414 21710
rect 31448 21676 31504 21710
rect 31538 21676 31594 21710
rect 31628 21676 31684 21710
rect 31718 21676 31774 21710
rect 31808 21676 31864 21710
rect 31898 21676 31950 21710
rect 31270 21620 31950 21676
rect 31270 21586 31324 21620
rect 31358 21586 31414 21620
rect 31448 21586 31504 21620
rect 31538 21586 31594 21620
rect 31628 21586 31684 21620
rect 31718 21586 31774 21620
rect 31808 21586 31864 21620
rect 31898 21586 31950 21620
rect 31270 21530 31950 21586
rect 31270 21496 31324 21530
rect 31358 21496 31414 21530
rect 31448 21496 31504 21530
rect 31538 21496 31594 21530
rect 31628 21496 31684 21530
rect 31718 21496 31774 21530
rect 31808 21496 31864 21530
rect 31898 21496 31950 21530
rect 31270 21440 31950 21496
rect 31270 21406 31324 21440
rect 31358 21406 31414 21440
rect 31448 21406 31504 21440
rect 31538 21406 31594 21440
rect 31628 21406 31684 21440
rect 31718 21406 31774 21440
rect 31808 21406 31864 21440
rect 31898 21406 31950 21440
rect 31270 21352 31950 21406
rect 32610 21980 33290 22032
rect 32610 21946 32664 21980
rect 32698 21946 32754 21980
rect 32788 21946 32844 21980
rect 32878 21946 32934 21980
rect 32968 21946 33024 21980
rect 33058 21946 33114 21980
rect 33148 21946 33204 21980
rect 33238 21946 33290 21980
rect 32610 21890 33290 21946
rect 32610 21856 32664 21890
rect 32698 21856 32754 21890
rect 32788 21856 32844 21890
rect 32878 21856 32934 21890
rect 32968 21856 33024 21890
rect 33058 21856 33114 21890
rect 33148 21856 33204 21890
rect 33238 21856 33290 21890
rect 32610 21800 33290 21856
rect 32610 21766 32664 21800
rect 32698 21766 32754 21800
rect 32788 21766 32844 21800
rect 32878 21766 32934 21800
rect 32968 21766 33024 21800
rect 33058 21766 33114 21800
rect 33148 21766 33204 21800
rect 33238 21766 33290 21800
rect 32610 21710 33290 21766
rect 32610 21676 32664 21710
rect 32698 21676 32754 21710
rect 32788 21676 32844 21710
rect 32878 21676 32934 21710
rect 32968 21676 33024 21710
rect 33058 21676 33114 21710
rect 33148 21676 33204 21710
rect 33238 21676 33290 21710
rect 32610 21620 33290 21676
rect 32610 21586 32664 21620
rect 32698 21586 32754 21620
rect 32788 21586 32844 21620
rect 32878 21586 32934 21620
rect 32968 21586 33024 21620
rect 33058 21586 33114 21620
rect 33148 21586 33204 21620
rect 33238 21586 33290 21620
rect 32610 21530 33290 21586
rect 32610 21496 32664 21530
rect 32698 21496 32754 21530
rect 32788 21496 32844 21530
rect 32878 21496 32934 21530
rect 32968 21496 33024 21530
rect 33058 21496 33114 21530
rect 33148 21496 33204 21530
rect 33238 21496 33290 21530
rect 32610 21440 33290 21496
rect 32610 21406 32664 21440
rect 32698 21406 32754 21440
rect 32788 21406 32844 21440
rect 32878 21406 32934 21440
rect 32968 21406 33024 21440
rect 33058 21406 33114 21440
rect 33148 21406 33204 21440
rect 33238 21406 33290 21440
rect 32610 21352 33290 21406
rect 33950 21980 34630 22032
rect 33950 21946 34004 21980
rect 34038 21946 34094 21980
rect 34128 21946 34184 21980
rect 34218 21946 34274 21980
rect 34308 21946 34364 21980
rect 34398 21946 34454 21980
rect 34488 21946 34544 21980
rect 34578 21946 34630 21980
rect 33950 21890 34630 21946
rect 33950 21856 34004 21890
rect 34038 21856 34094 21890
rect 34128 21856 34184 21890
rect 34218 21856 34274 21890
rect 34308 21856 34364 21890
rect 34398 21856 34454 21890
rect 34488 21856 34544 21890
rect 34578 21856 34630 21890
rect 33950 21800 34630 21856
rect 33950 21766 34004 21800
rect 34038 21766 34094 21800
rect 34128 21766 34184 21800
rect 34218 21766 34274 21800
rect 34308 21766 34364 21800
rect 34398 21766 34454 21800
rect 34488 21766 34544 21800
rect 34578 21766 34630 21800
rect 33950 21710 34630 21766
rect 33950 21676 34004 21710
rect 34038 21676 34094 21710
rect 34128 21676 34184 21710
rect 34218 21676 34274 21710
rect 34308 21676 34364 21710
rect 34398 21676 34454 21710
rect 34488 21676 34544 21710
rect 34578 21676 34630 21710
rect 33950 21620 34630 21676
rect 33950 21586 34004 21620
rect 34038 21586 34094 21620
rect 34128 21586 34184 21620
rect 34218 21586 34274 21620
rect 34308 21586 34364 21620
rect 34398 21586 34454 21620
rect 34488 21586 34544 21620
rect 34578 21586 34630 21620
rect 33950 21530 34630 21586
rect 33950 21496 34004 21530
rect 34038 21496 34094 21530
rect 34128 21496 34184 21530
rect 34218 21496 34274 21530
rect 34308 21496 34364 21530
rect 34398 21496 34454 21530
rect 34488 21496 34544 21530
rect 34578 21496 34630 21530
rect 33950 21440 34630 21496
rect 33950 21406 34004 21440
rect 34038 21406 34094 21440
rect 34128 21406 34184 21440
rect 34218 21406 34274 21440
rect 34308 21406 34364 21440
rect 34398 21406 34454 21440
rect 34488 21406 34544 21440
rect 34578 21406 34630 21440
rect 33950 21352 34630 21406
rect 35290 21980 35970 22032
rect 35290 21946 35344 21980
rect 35378 21946 35434 21980
rect 35468 21946 35524 21980
rect 35558 21946 35614 21980
rect 35648 21946 35704 21980
rect 35738 21946 35794 21980
rect 35828 21946 35884 21980
rect 35918 21946 35970 21980
rect 35290 21890 35970 21946
rect 35290 21856 35344 21890
rect 35378 21856 35434 21890
rect 35468 21856 35524 21890
rect 35558 21856 35614 21890
rect 35648 21856 35704 21890
rect 35738 21856 35794 21890
rect 35828 21856 35884 21890
rect 35918 21856 35970 21890
rect 35290 21800 35970 21856
rect 35290 21766 35344 21800
rect 35378 21766 35434 21800
rect 35468 21766 35524 21800
rect 35558 21766 35614 21800
rect 35648 21766 35704 21800
rect 35738 21766 35794 21800
rect 35828 21766 35884 21800
rect 35918 21766 35970 21800
rect 35290 21710 35970 21766
rect 35290 21676 35344 21710
rect 35378 21676 35434 21710
rect 35468 21676 35524 21710
rect 35558 21676 35614 21710
rect 35648 21676 35704 21710
rect 35738 21676 35794 21710
rect 35828 21676 35884 21710
rect 35918 21676 35970 21710
rect 35290 21620 35970 21676
rect 35290 21586 35344 21620
rect 35378 21586 35434 21620
rect 35468 21586 35524 21620
rect 35558 21586 35614 21620
rect 35648 21586 35704 21620
rect 35738 21586 35794 21620
rect 35828 21586 35884 21620
rect 35918 21586 35970 21620
rect 35290 21530 35970 21586
rect 35290 21496 35344 21530
rect 35378 21496 35434 21530
rect 35468 21496 35524 21530
rect 35558 21496 35614 21530
rect 35648 21496 35704 21530
rect 35738 21496 35794 21530
rect 35828 21496 35884 21530
rect 35918 21496 35970 21530
rect 35290 21440 35970 21496
rect 35290 21406 35344 21440
rect 35378 21406 35434 21440
rect 35468 21406 35524 21440
rect 35558 21406 35614 21440
rect 35648 21406 35704 21440
rect 35738 21406 35794 21440
rect 35828 21406 35884 21440
rect 35918 21406 35970 21440
rect 35290 21352 35970 21406
rect 36630 21980 37310 22032
rect 36630 21946 36684 21980
rect 36718 21946 36774 21980
rect 36808 21946 36864 21980
rect 36898 21946 36954 21980
rect 36988 21946 37044 21980
rect 37078 21946 37134 21980
rect 37168 21946 37224 21980
rect 37258 21946 37310 21980
rect 36630 21890 37310 21946
rect 36630 21856 36684 21890
rect 36718 21856 36774 21890
rect 36808 21856 36864 21890
rect 36898 21856 36954 21890
rect 36988 21856 37044 21890
rect 37078 21856 37134 21890
rect 37168 21856 37224 21890
rect 37258 21856 37310 21890
rect 36630 21800 37310 21856
rect 36630 21766 36684 21800
rect 36718 21766 36774 21800
rect 36808 21766 36864 21800
rect 36898 21766 36954 21800
rect 36988 21766 37044 21800
rect 37078 21766 37134 21800
rect 37168 21766 37224 21800
rect 37258 21766 37310 21800
rect 36630 21710 37310 21766
rect 36630 21676 36684 21710
rect 36718 21676 36774 21710
rect 36808 21676 36864 21710
rect 36898 21676 36954 21710
rect 36988 21676 37044 21710
rect 37078 21676 37134 21710
rect 37168 21676 37224 21710
rect 37258 21676 37310 21710
rect 36630 21620 37310 21676
rect 36630 21586 36684 21620
rect 36718 21586 36774 21620
rect 36808 21586 36864 21620
rect 36898 21586 36954 21620
rect 36988 21586 37044 21620
rect 37078 21586 37134 21620
rect 37168 21586 37224 21620
rect 37258 21586 37310 21620
rect 36630 21530 37310 21586
rect 36630 21496 36684 21530
rect 36718 21496 36774 21530
rect 36808 21496 36864 21530
rect 36898 21496 36954 21530
rect 36988 21496 37044 21530
rect 37078 21496 37134 21530
rect 37168 21496 37224 21530
rect 37258 21496 37310 21530
rect 36630 21440 37310 21496
rect 36630 21406 36684 21440
rect 36718 21406 36774 21440
rect 36808 21406 36864 21440
rect 36898 21406 36954 21440
rect 36988 21406 37044 21440
rect 37078 21406 37134 21440
rect 37168 21406 37224 21440
rect 37258 21406 37310 21440
rect 36630 21352 37310 21406
rect 37970 21980 38650 22032
rect 37970 21946 38024 21980
rect 38058 21946 38114 21980
rect 38148 21946 38204 21980
rect 38238 21946 38294 21980
rect 38328 21946 38384 21980
rect 38418 21946 38474 21980
rect 38508 21946 38564 21980
rect 38598 21946 38650 21980
rect 37970 21890 38650 21946
rect 37970 21856 38024 21890
rect 38058 21856 38114 21890
rect 38148 21856 38204 21890
rect 38238 21856 38294 21890
rect 38328 21856 38384 21890
rect 38418 21856 38474 21890
rect 38508 21856 38564 21890
rect 38598 21856 38650 21890
rect 37970 21800 38650 21856
rect 37970 21766 38024 21800
rect 38058 21766 38114 21800
rect 38148 21766 38204 21800
rect 38238 21766 38294 21800
rect 38328 21766 38384 21800
rect 38418 21766 38474 21800
rect 38508 21766 38564 21800
rect 38598 21766 38650 21800
rect 37970 21710 38650 21766
rect 37970 21676 38024 21710
rect 38058 21676 38114 21710
rect 38148 21676 38204 21710
rect 38238 21676 38294 21710
rect 38328 21676 38384 21710
rect 38418 21676 38474 21710
rect 38508 21676 38564 21710
rect 38598 21676 38650 21710
rect 37970 21620 38650 21676
rect 37970 21586 38024 21620
rect 38058 21586 38114 21620
rect 38148 21586 38204 21620
rect 38238 21586 38294 21620
rect 38328 21586 38384 21620
rect 38418 21586 38474 21620
rect 38508 21586 38564 21620
rect 38598 21586 38650 21620
rect 37970 21530 38650 21586
rect 37970 21496 38024 21530
rect 38058 21496 38114 21530
rect 38148 21496 38204 21530
rect 38238 21496 38294 21530
rect 38328 21496 38384 21530
rect 38418 21496 38474 21530
rect 38508 21496 38564 21530
rect 38598 21496 38650 21530
rect 37970 21440 38650 21496
rect 37970 21406 38024 21440
rect 38058 21406 38114 21440
rect 38148 21406 38204 21440
rect 38238 21406 38294 21440
rect 38328 21406 38384 21440
rect 38418 21406 38474 21440
rect 38508 21406 38564 21440
rect 38598 21406 38650 21440
rect 37970 21352 38650 21406
rect 23983 18621 24041 18637
rect 23983 18587 23995 18621
rect 24029 18587 24041 18621
rect 23983 18553 24041 18587
rect 23983 18519 23995 18553
rect 24029 18519 24041 18553
rect 23983 18485 24041 18519
rect 23983 18451 23995 18485
rect 24029 18451 24041 18485
rect 23983 18417 24041 18451
rect 23983 18383 23995 18417
rect 24029 18383 24041 18417
rect 23983 18349 24041 18383
rect 23983 18315 23995 18349
rect 24029 18315 24041 18349
rect 23983 18281 24041 18315
rect 23983 18247 23995 18281
rect 24029 18247 24041 18281
rect 23983 18213 24041 18247
rect 23983 18179 23995 18213
rect 24029 18179 24041 18213
rect 23983 18145 24041 18179
rect 23983 18111 23995 18145
rect 24029 18111 24041 18145
rect 23983 18077 24041 18111
rect 23983 18043 23995 18077
rect 24029 18043 24041 18077
rect 23983 18009 24041 18043
rect 23983 17975 23995 18009
rect 24029 17975 24041 18009
rect 23983 17941 24041 17975
rect 23983 17907 23995 17941
rect 24029 17907 24041 17941
rect 23983 17873 24041 17907
rect 23983 17839 23995 17873
rect 24029 17839 24041 17873
rect 23983 17805 24041 17839
rect 23983 17771 23995 17805
rect 24029 17771 24041 17805
rect 23983 17737 24041 17771
rect 23983 17703 23995 17737
rect 24029 17703 24041 17737
rect 23983 17669 24041 17703
rect 23983 17635 23995 17669
rect 24029 17635 24041 17669
rect 23983 17601 24041 17635
rect 23983 17567 23995 17601
rect 24029 17567 24041 17601
rect 23983 17533 24041 17567
rect 23983 17499 23995 17533
rect 24029 17499 24041 17533
rect 23983 17465 24041 17499
rect 23983 17431 23995 17465
rect 24029 17431 24041 17465
rect 23983 17397 24041 17431
rect 23983 17363 23995 17397
rect 24029 17363 24041 17397
rect 23983 17347 24041 17363
rect 24441 18621 24499 18637
rect 24441 18587 24453 18621
rect 24487 18587 24499 18621
rect 24441 18553 24499 18587
rect 24441 18519 24453 18553
rect 24487 18519 24499 18553
rect 24441 18485 24499 18519
rect 24441 18451 24453 18485
rect 24487 18451 24499 18485
rect 24441 18417 24499 18451
rect 24441 18383 24453 18417
rect 24487 18383 24499 18417
rect 24441 18349 24499 18383
rect 24441 18315 24453 18349
rect 24487 18315 24499 18349
rect 24441 18281 24499 18315
rect 24441 18247 24453 18281
rect 24487 18247 24499 18281
rect 24441 18213 24499 18247
rect 24441 18179 24453 18213
rect 24487 18179 24499 18213
rect 24441 18145 24499 18179
rect 24441 18111 24453 18145
rect 24487 18111 24499 18145
rect 24441 18077 24499 18111
rect 24441 18043 24453 18077
rect 24487 18043 24499 18077
rect 24441 18009 24499 18043
rect 24441 17975 24453 18009
rect 24487 17975 24499 18009
rect 24441 17941 24499 17975
rect 24441 17907 24453 17941
rect 24487 17907 24499 17941
rect 24441 17873 24499 17907
rect 24441 17839 24453 17873
rect 24487 17839 24499 17873
rect 24441 17805 24499 17839
rect 24441 17771 24453 17805
rect 24487 17771 24499 17805
rect 24441 17737 24499 17771
rect 24441 17703 24453 17737
rect 24487 17703 24499 17737
rect 24441 17669 24499 17703
rect 24441 17635 24453 17669
rect 24487 17635 24499 17669
rect 24441 17601 24499 17635
rect 24441 17567 24453 17601
rect 24487 17567 24499 17601
rect 24441 17533 24499 17567
rect 24441 17499 24453 17533
rect 24487 17499 24499 17533
rect 24441 17465 24499 17499
rect 24441 17431 24453 17465
rect 24487 17431 24499 17465
rect 24441 17397 24499 17431
rect 24441 17363 24453 17397
rect 24487 17363 24499 17397
rect 24441 17347 24499 17363
rect 24899 18621 24957 18637
rect 24899 18587 24911 18621
rect 24945 18587 24957 18621
rect 24899 18553 24957 18587
rect 24899 18519 24911 18553
rect 24945 18519 24957 18553
rect 24899 18485 24957 18519
rect 24899 18451 24911 18485
rect 24945 18451 24957 18485
rect 24899 18417 24957 18451
rect 24899 18383 24911 18417
rect 24945 18383 24957 18417
rect 24899 18349 24957 18383
rect 24899 18315 24911 18349
rect 24945 18315 24957 18349
rect 24899 18281 24957 18315
rect 24899 18247 24911 18281
rect 24945 18247 24957 18281
rect 24899 18213 24957 18247
rect 24899 18179 24911 18213
rect 24945 18179 24957 18213
rect 24899 18145 24957 18179
rect 24899 18111 24911 18145
rect 24945 18111 24957 18145
rect 24899 18077 24957 18111
rect 24899 18043 24911 18077
rect 24945 18043 24957 18077
rect 24899 18009 24957 18043
rect 24899 17975 24911 18009
rect 24945 17975 24957 18009
rect 24899 17941 24957 17975
rect 24899 17907 24911 17941
rect 24945 17907 24957 17941
rect 24899 17873 24957 17907
rect 24899 17839 24911 17873
rect 24945 17839 24957 17873
rect 24899 17805 24957 17839
rect 24899 17771 24911 17805
rect 24945 17771 24957 17805
rect 24899 17737 24957 17771
rect 24899 17703 24911 17737
rect 24945 17703 24957 17737
rect 24899 17669 24957 17703
rect 24899 17635 24911 17669
rect 24945 17635 24957 17669
rect 24899 17601 24957 17635
rect 24899 17567 24911 17601
rect 24945 17567 24957 17601
rect 24899 17533 24957 17567
rect 24899 17499 24911 17533
rect 24945 17499 24957 17533
rect 24899 17465 24957 17499
rect 24899 17431 24911 17465
rect 24945 17431 24957 17465
rect 24899 17397 24957 17431
rect 24899 17363 24911 17397
rect 24945 17363 24957 17397
rect 24899 17347 24957 17363
rect 25357 18621 25415 18637
rect 25357 18587 25369 18621
rect 25403 18587 25415 18621
rect 25357 18553 25415 18587
rect 25357 18519 25369 18553
rect 25403 18519 25415 18553
rect 25357 18485 25415 18519
rect 25357 18451 25369 18485
rect 25403 18451 25415 18485
rect 25357 18417 25415 18451
rect 25357 18383 25369 18417
rect 25403 18383 25415 18417
rect 25357 18349 25415 18383
rect 25357 18315 25369 18349
rect 25403 18315 25415 18349
rect 25357 18281 25415 18315
rect 25357 18247 25369 18281
rect 25403 18247 25415 18281
rect 25357 18213 25415 18247
rect 25357 18179 25369 18213
rect 25403 18179 25415 18213
rect 25357 18145 25415 18179
rect 25357 18111 25369 18145
rect 25403 18111 25415 18145
rect 25357 18077 25415 18111
rect 25357 18043 25369 18077
rect 25403 18043 25415 18077
rect 25357 18009 25415 18043
rect 25357 17975 25369 18009
rect 25403 17975 25415 18009
rect 25357 17941 25415 17975
rect 25357 17907 25369 17941
rect 25403 17907 25415 17941
rect 25357 17873 25415 17907
rect 25357 17839 25369 17873
rect 25403 17839 25415 17873
rect 25357 17805 25415 17839
rect 25357 17771 25369 17805
rect 25403 17771 25415 17805
rect 25357 17737 25415 17771
rect 25357 17703 25369 17737
rect 25403 17703 25415 17737
rect 25357 17669 25415 17703
rect 25357 17635 25369 17669
rect 25403 17635 25415 17669
rect 25357 17601 25415 17635
rect 25357 17567 25369 17601
rect 25403 17567 25415 17601
rect 25357 17533 25415 17567
rect 25357 17499 25369 17533
rect 25403 17499 25415 17533
rect 25357 17465 25415 17499
rect 25357 17431 25369 17465
rect 25403 17431 25415 17465
rect 25357 17397 25415 17431
rect 25357 17363 25369 17397
rect 25403 17363 25415 17397
rect 25357 17347 25415 17363
rect 25815 18621 25873 18637
rect 25815 18587 25827 18621
rect 25861 18587 25873 18621
rect 25815 18553 25873 18587
rect 25815 18519 25827 18553
rect 25861 18519 25873 18553
rect 25815 18485 25873 18519
rect 25815 18451 25827 18485
rect 25861 18451 25873 18485
rect 25815 18417 25873 18451
rect 25815 18383 25827 18417
rect 25861 18383 25873 18417
rect 25815 18349 25873 18383
rect 25815 18315 25827 18349
rect 25861 18315 25873 18349
rect 25815 18281 25873 18315
rect 25815 18247 25827 18281
rect 25861 18247 25873 18281
rect 25815 18213 25873 18247
rect 25815 18179 25827 18213
rect 25861 18179 25873 18213
rect 25815 18145 25873 18179
rect 25815 18111 25827 18145
rect 25861 18111 25873 18145
rect 25815 18077 25873 18111
rect 25815 18043 25827 18077
rect 25861 18043 25873 18077
rect 25815 18009 25873 18043
rect 25815 17975 25827 18009
rect 25861 17975 25873 18009
rect 25815 17941 25873 17975
rect 25815 17907 25827 17941
rect 25861 17907 25873 17941
rect 25815 17873 25873 17907
rect 25815 17839 25827 17873
rect 25861 17839 25873 17873
rect 25815 17805 25873 17839
rect 25815 17771 25827 17805
rect 25861 17771 25873 17805
rect 25815 17737 25873 17771
rect 25815 17703 25827 17737
rect 25861 17703 25873 17737
rect 25815 17669 25873 17703
rect 25815 17635 25827 17669
rect 25861 17635 25873 17669
rect 25815 17601 25873 17635
rect 25815 17567 25827 17601
rect 25861 17567 25873 17601
rect 25815 17533 25873 17567
rect 25815 17499 25827 17533
rect 25861 17499 25873 17533
rect 25815 17465 25873 17499
rect 25815 17431 25827 17465
rect 25861 17431 25873 17465
rect 25815 17397 25873 17431
rect 25815 17363 25827 17397
rect 25861 17363 25873 17397
rect 25815 17347 25873 17363
rect 26273 18621 26331 18637
rect 26273 18587 26285 18621
rect 26319 18587 26331 18621
rect 26273 18553 26331 18587
rect 26273 18519 26285 18553
rect 26319 18519 26331 18553
rect 26273 18485 26331 18519
rect 26273 18451 26285 18485
rect 26319 18451 26331 18485
rect 26273 18417 26331 18451
rect 26273 18383 26285 18417
rect 26319 18383 26331 18417
rect 26273 18349 26331 18383
rect 26273 18315 26285 18349
rect 26319 18315 26331 18349
rect 26273 18281 26331 18315
rect 26273 18247 26285 18281
rect 26319 18247 26331 18281
rect 26273 18213 26331 18247
rect 26273 18179 26285 18213
rect 26319 18179 26331 18213
rect 26273 18145 26331 18179
rect 26273 18111 26285 18145
rect 26319 18111 26331 18145
rect 26273 18077 26331 18111
rect 26273 18043 26285 18077
rect 26319 18043 26331 18077
rect 26273 18009 26331 18043
rect 26273 17975 26285 18009
rect 26319 17975 26331 18009
rect 26273 17941 26331 17975
rect 26273 17907 26285 17941
rect 26319 17907 26331 17941
rect 26273 17873 26331 17907
rect 26273 17839 26285 17873
rect 26319 17839 26331 17873
rect 26273 17805 26331 17839
rect 26273 17771 26285 17805
rect 26319 17771 26331 17805
rect 26273 17737 26331 17771
rect 26273 17703 26285 17737
rect 26319 17703 26331 17737
rect 26273 17669 26331 17703
rect 26273 17635 26285 17669
rect 26319 17635 26331 17669
rect 26273 17601 26331 17635
rect 26273 17567 26285 17601
rect 26319 17567 26331 17601
rect 26273 17533 26331 17567
rect 26273 17499 26285 17533
rect 26319 17499 26331 17533
rect 26273 17465 26331 17499
rect 26273 17431 26285 17465
rect 26319 17431 26331 17465
rect 26273 17397 26331 17431
rect 26273 17363 26285 17397
rect 26319 17363 26331 17397
rect 26273 17347 26331 17363
rect 26731 18621 26789 18637
rect 26731 18587 26743 18621
rect 26777 18587 26789 18621
rect 26731 18553 26789 18587
rect 26731 18519 26743 18553
rect 26777 18519 26789 18553
rect 26731 18485 26789 18519
rect 26731 18451 26743 18485
rect 26777 18451 26789 18485
rect 26731 18417 26789 18451
rect 26731 18383 26743 18417
rect 26777 18383 26789 18417
rect 26731 18349 26789 18383
rect 26731 18315 26743 18349
rect 26777 18315 26789 18349
rect 26731 18281 26789 18315
rect 26731 18247 26743 18281
rect 26777 18247 26789 18281
rect 26731 18213 26789 18247
rect 26731 18179 26743 18213
rect 26777 18179 26789 18213
rect 26731 18145 26789 18179
rect 26731 18111 26743 18145
rect 26777 18111 26789 18145
rect 26731 18077 26789 18111
rect 26731 18043 26743 18077
rect 26777 18043 26789 18077
rect 26731 18009 26789 18043
rect 26731 17975 26743 18009
rect 26777 17975 26789 18009
rect 26731 17941 26789 17975
rect 26731 17907 26743 17941
rect 26777 17907 26789 17941
rect 26731 17873 26789 17907
rect 26731 17839 26743 17873
rect 26777 17839 26789 17873
rect 26731 17805 26789 17839
rect 26731 17771 26743 17805
rect 26777 17771 26789 17805
rect 26731 17737 26789 17771
rect 26731 17703 26743 17737
rect 26777 17703 26789 17737
rect 26731 17669 26789 17703
rect 26731 17635 26743 17669
rect 26777 17635 26789 17669
rect 26731 17601 26789 17635
rect 26731 17567 26743 17601
rect 26777 17567 26789 17601
rect 26731 17533 26789 17567
rect 26731 17499 26743 17533
rect 26777 17499 26789 17533
rect 26731 17465 26789 17499
rect 26731 17431 26743 17465
rect 26777 17431 26789 17465
rect 26731 17397 26789 17431
rect 26731 17363 26743 17397
rect 26777 17363 26789 17397
rect 26731 17347 26789 17363
rect 28590 18220 29270 18272
rect 28590 18186 28644 18220
rect 28678 18186 28734 18220
rect 28768 18186 28824 18220
rect 28858 18186 28914 18220
rect 28948 18186 29004 18220
rect 29038 18186 29094 18220
rect 29128 18186 29184 18220
rect 29218 18186 29270 18220
rect 28590 18130 29270 18186
rect 28590 18096 28644 18130
rect 28678 18096 28734 18130
rect 28768 18096 28824 18130
rect 28858 18096 28914 18130
rect 28948 18096 29004 18130
rect 29038 18096 29094 18130
rect 29128 18096 29184 18130
rect 29218 18096 29270 18130
rect 28590 18040 29270 18096
rect 28590 18006 28644 18040
rect 28678 18006 28734 18040
rect 28768 18006 28824 18040
rect 28858 18006 28914 18040
rect 28948 18006 29004 18040
rect 29038 18006 29094 18040
rect 29128 18006 29184 18040
rect 29218 18006 29270 18040
rect 28590 17950 29270 18006
rect 28590 17916 28644 17950
rect 28678 17916 28734 17950
rect 28768 17916 28824 17950
rect 28858 17916 28914 17950
rect 28948 17916 29004 17950
rect 29038 17916 29094 17950
rect 29128 17916 29184 17950
rect 29218 17916 29270 17950
rect 28590 17860 29270 17916
rect 28590 17826 28644 17860
rect 28678 17826 28734 17860
rect 28768 17826 28824 17860
rect 28858 17826 28914 17860
rect 28948 17826 29004 17860
rect 29038 17826 29094 17860
rect 29128 17826 29184 17860
rect 29218 17826 29270 17860
rect 28590 17770 29270 17826
rect 28590 17736 28644 17770
rect 28678 17736 28734 17770
rect 28768 17736 28824 17770
rect 28858 17736 28914 17770
rect 28948 17736 29004 17770
rect 29038 17736 29094 17770
rect 29128 17736 29184 17770
rect 29218 17736 29270 17770
rect 28590 17680 29270 17736
rect 28590 17646 28644 17680
rect 28678 17646 28734 17680
rect 28768 17646 28824 17680
rect 28858 17646 28914 17680
rect 28948 17646 29004 17680
rect 29038 17646 29094 17680
rect 29128 17646 29184 17680
rect 29218 17646 29270 17680
rect 28590 17592 29270 17646
rect 29930 18220 30610 18272
rect 29930 18186 29984 18220
rect 30018 18186 30074 18220
rect 30108 18186 30164 18220
rect 30198 18186 30254 18220
rect 30288 18186 30344 18220
rect 30378 18186 30434 18220
rect 30468 18186 30524 18220
rect 30558 18186 30610 18220
rect 29930 18130 30610 18186
rect 29930 18096 29984 18130
rect 30018 18096 30074 18130
rect 30108 18096 30164 18130
rect 30198 18096 30254 18130
rect 30288 18096 30344 18130
rect 30378 18096 30434 18130
rect 30468 18096 30524 18130
rect 30558 18096 30610 18130
rect 29930 18040 30610 18096
rect 29930 18006 29984 18040
rect 30018 18006 30074 18040
rect 30108 18006 30164 18040
rect 30198 18006 30254 18040
rect 30288 18006 30344 18040
rect 30378 18006 30434 18040
rect 30468 18006 30524 18040
rect 30558 18006 30610 18040
rect 29930 17950 30610 18006
rect 29930 17916 29984 17950
rect 30018 17916 30074 17950
rect 30108 17916 30164 17950
rect 30198 17916 30254 17950
rect 30288 17916 30344 17950
rect 30378 17916 30434 17950
rect 30468 17916 30524 17950
rect 30558 17916 30610 17950
rect 29930 17860 30610 17916
rect 29930 17826 29984 17860
rect 30018 17826 30074 17860
rect 30108 17826 30164 17860
rect 30198 17826 30254 17860
rect 30288 17826 30344 17860
rect 30378 17826 30434 17860
rect 30468 17826 30524 17860
rect 30558 17826 30610 17860
rect 29930 17770 30610 17826
rect 29930 17736 29984 17770
rect 30018 17736 30074 17770
rect 30108 17736 30164 17770
rect 30198 17736 30254 17770
rect 30288 17736 30344 17770
rect 30378 17736 30434 17770
rect 30468 17736 30524 17770
rect 30558 17736 30610 17770
rect 29930 17680 30610 17736
rect 29930 17646 29984 17680
rect 30018 17646 30074 17680
rect 30108 17646 30164 17680
rect 30198 17646 30254 17680
rect 30288 17646 30344 17680
rect 30378 17646 30434 17680
rect 30468 17646 30524 17680
rect 30558 17646 30610 17680
rect 29930 17592 30610 17646
rect 31270 18220 31950 18272
rect 31270 18186 31324 18220
rect 31358 18186 31414 18220
rect 31448 18186 31504 18220
rect 31538 18186 31594 18220
rect 31628 18186 31684 18220
rect 31718 18186 31774 18220
rect 31808 18186 31864 18220
rect 31898 18186 31950 18220
rect 31270 18130 31950 18186
rect 31270 18096 31324 18130
rect 31358 18096 31414 18130
rect 31448 18096 31504 18130
rect 31538 18096 31594 18130
rect 31628 18096 31684 18130
rect 31718 18096 31774 18130
rect 31808 18096 31864 18130
rect 31898 18096 31950 18130
rect 31270 18040 31950 18096
rect 31270 18006 31324 18040
rect 31358 18006 31414 18040
rect 31448 18006 31504 18040
rect 31538 18006 31594 18040
rect 31628 18006 31684 18040
rect 31718 18006 31774 18040
rect 31808 18006 31864 18040
rect 31898 18006 31950 18040
rect 31270 17950 31950 18006
rect 31270 17916 31324 17950
rect 31358 17916 31414 17950
rect 31448 17916 31504 17950
rect 31538 17916 31594 17950
rect 31628 17916 31684 17950
rect 31718 17916 31774 17950
rect 31808 17916 31864 17950
rect 31898 17916 31950 17950
rect 31270 17860 31950 17916
rect 31270 17826 31324 17860
rect 31358 17826 31414 17860
rect 31448 17826 31504 17860
rect 31538 17826 31594 17860
rect 31628 17826 31684 17860
rect 31718 17826 31774 17860
rect 31808 17826 31864 17860
rect 31898 17826 31950 17860
rect 31270 17770 31950 17826
rect 31270 17736 31324 17770
rect 31358 17736 31414 17770
rect 31448 17736 31504 17770
rect 31538 17736 31594 17770
rect 31628 17736 31684 17770
rect 31718 17736 31774 17770
rect 31808 17736 31864 17770
rect 31898 17736 31950 17770
rect 31270 17680 31950 17736
rect 31270 17646 31324 17680
rect 31358 17646 31414 17680
rect 31448 17646 31504 17680
rect 31538 17646 31594 17680
rect 31628 17646 31684 17680
rect 31718 17646 31774 17680
rect 31808 17646 31864 17680
rect 31898 17646 31950 17680
rect 31270 17592 31950 17646
rect 32610 18220 33290 18272
rect 32610 18186 32664 18220
rect 32698 18186 32754 18220
rect 32788 18186 32844 18220
rect 32878 18186 32934 18220
rect 32968 18186 33024 18220
rect 33058 18186 33114 18220
rect 33148 18186 33204 18220
rect 33238 18186 33290 18220
rect 32610 18130 33290 18186
rect 32610 18096 32664 18130
rect 32698 18096 32754 18130
rect 32788 18096 32844 18130
rect 32878 18096 32934 18130
rect 32968 18096 33024 18130
rect 33058 18096 33114 18130
rect 33148 18096 33204 18130
rect 33238 18096 33290 18130
rect 32610 18040 33290 18096
rect 32610 18006 32664 18040
rect 32698 18006 32754 18040
rect 32788 18006 32844 18040
rect 32878 18006 32934 18040
rect 32968 18006 33024 18040
rect 33058 18006 33114 18040
rect 33148 18006 33204 18040
rect 33238 18006 33290 18040
rect 32610 17950 33290 18006
rect 32610 17916 32664 17950
rect 32698 17916 32754 17950
rect 32788 17916 32844 17950
rect 32878 17916 32934 17950
rect 32968 17916 33024 17950
rect 33058 17916 33114 17950
rect 33148 17916 33204 17950
rect 33238 17916 33290 17950
rect 32610 17860 33290 17916
rect 32610 17826 32664 17860
rect 32698 17826 32754 17860
rect 32788 17826 32844 17860
rect 32878 17826 32934 17860
rect 32968 17826 33024 17860
rect 33058 17826 33114 17860
rect 33148 17826 33204 17860
rect 33238 17826 33290 17860
rect 32610 17770 33290 17826
rect 32610 17736 32664 17770
rect 32698 17736 32754 17770
rect 32788 17736 32844 17770
rect 32878 17736 32934 17770
rect 32968 17736 33024 17770
rect 33058 17736 33114 17770
rect 33148 17736 33204 17770
rect 33238 17736 33290 17770
rect 32610 17680 33290 17736
rect 32610 17646 32664 17680
rect 32698 17646 32754 17680
rect 32788 17646 32844 17680
rect 32878 17646 32934 17680
rect 32968 17646 33024 17680
rect 33058 17646 33114 17680
rect 33148 17646 33204 17680
rect 33238 17646 33290 17680
rect 32610 17592 33290 17646
rect 33950 18220 34630 18272
rect 33950 18186 34004 18220
rect 34038 18186 34094 18220
rect 34128 18186 34184 18220
rect 34218 18186 34274 18220
rect 34308 18186 34364 18220
rect 34398 18186 34454 18220
rect 34488 18186 34544 18220
rect 34578 18186 34630 18220
rect 33950 18130 34630 18186
rect 33950 18096 34004 18130
rect 34038 18096 34094 18130
rect 34128 18096 34184 18130
rect 34218 18096 34274 18130
rect 34308 18096 34364 18130
rect 34398 18096 34454 18130
rect 34488 18096 34544 18130
rect 34578 18096 34630 18130
rect 33950 18040 34630 18096
rect 33950 18006 34004 18040
rect 34038 18006 34094 18040
rect 34128 18006 34184 18040
rect 34218 18006 34274 18040
rect 34308 18006 34364 18040
rect 34398 18006 34454 18040
rect 34488 18006 34544 18040
rect 34578 18006 34630 18040
rect 33950 17950 34630 18006
rect 33950 17916 34004 17950
rect 34038 17916 34094 17950
rect 34128 17916 34184 17950
rect 34218 17916 34274 17950
rect 34308 17916 34364 17950
rect 34398 17916 34454 17950
rect 34488 17916 34544 17950
rect 34578 17916 34630 17950
rect 33950 17860 34630 17916
rect 33950 17826 34004 17860
rect 34038 17826 34094 17860
rect 34128 17826 34184 17860
rect 34218 17826 34274 17860
rect 34308 17826 34364 17860
rect 34398 17826 34454 17860
rect 34488 17826 34544 17860
rect 34578 17826 34630 17860
rect 33950 17770 34630 17826
rect 33950 17736 34004 17770
rect 34038 17736 34094 17770
rect 34128 17736 34184 17770
rect 34218 17736 34274 17770
rect 34308 17736 34364 17770
rect 34398 17736 34454 17770
rect 34488 17736 34544 17770
rect 34578 17736 34630 17770
rect 33950 17680 34630 17736
rect 33950 17646 34004 17680
rect 34038 17646 34094 17680
rect 34128 17646 34184 17680
rect 34218 17646 34274 17680
rect 34308 17646 34364 17680
rect 34398 17646 34454 17680
rect 34488 17646 34544 17680
rect 34578 17646 34630 17680
rect 33950 17592 34630 17646
rect 35290 18220 35970 18272
rect 35290 18186 35344 18220
rect 35378 18186 35434 18220
rect 35468 18186 35524 18220
rect 35558 18186 35614 18220
rect 35648 18186 35704 18220
rect 35738 18186 35794 18220
rect 35828 18186 35884 18220
rect 35918 18186 35970 18220
rect 35290 18130 35970 18186
rect 35290 18096 35344 18130
rect 35378 18096 35434 18130
rect 35468 18096 35524 18130
rect 35558 18096 35614 18130
rect 35648 18096 35704 18130
rect 35738 18096 35794 18130
rect 35828 18096 35884 18130
rect 35918 18096 35970 18130
rect 35290 18040 35970 18096
rect 35290 18006 35344 18040
rect 35378 18006 35434 18040
rect 35468 18006 35524 18040
rect 35558 18006 35614 18040
rect 35648 18006 35704 18040
rect 35738 18006 35794 18040
rect 35828 18006 35884 18040
rect 35918 18006 35970 18040
rect 35290 17950 35970 18006
rect 35290 17916 35344 17950
rect 35378 17916 35434 17950
rect 35468 17916 35524 17950
rect 35558 17916 35614 17950
rect 35648 17916 35704 17950
rect 35738 17916 35794 17950
rect 35828 17916 35884 17950
rect 35918 17916 35970 17950
rect 35290 17860 35970 17916
rect 35290 17826 35344 17860
rect 35378 17826 35434 17860
rect 35468 17826 35524 17860
rect 35558 17826 35614 17860
rect 35648 17826 35704 17860
rect 35738 17826 35794 17860
rect 35828 17826 35884 17860
rect 35918 17826 35970 17860
rect 35290 17770 35970 17826
rect 35290 17736 35344 17770
rect 35378 17736 35434 17770
rect 35468 17736 35524 17770
rect 35558 17736 35614 17770
rect 35648 17736 35704 17770
rect 35738 17736 35794 17770
rect 35828 17736 35884 17770
rect 35918 17736 35970 17770
rect 35290 17680 35970 17736
rect 35290 17646 35344 17680
rect 35378 17646 35434 17680
rect 35468 17646 35524 17680
rect 35558 17646 35614 17680
rect 35648 17646 35704 17680
rect 35738 17646 35794 17680
rect 35828 17646 35884 17680
rect 35918 17646 35970 17680
rect 35290 17592 35970 17646
rect 36630 18220 37310 18272
rect 36630 18186 36684 18220
rect 36718 18186 36774 18220
rect 36808 18186 36864 18220
rect 36898 18186 36954 18220
rect 36988 18186 37044 18220
rect 37078 18186 37134 18220
rect 37168 18186 37224 18220
rect 37258 18186 37310 18220
rect 36630 18130 37310 18186
rect 36630 18096 36684 18130
rect 36718 18096 36774 18130
rect 36808 18096 36864 18130
rect 36898 18096 36954 18130
rect 36988 18096 37044 18130
rect 37078 18096 37134 18130
rect 37168 18096 37224 18130
rect 37258 18096 37310 18130
rect 36630 18040 37310 18096
rect 36630 18006 36684 18040
rect 36718 18006 36774 18040
rect 36808 18006 36864 18040
rect 36898 18006 36954 18040
rect 36988 18006 37044 18040
rect 37078 18006 37134 18040
rect 37168 18006 37224 18040
rect 37258 18006 37310 18040
rect 36630 17950 37310 18006
rect 36630 17916 36684 17950
rect 36718 17916 36774 17950
rect 36808 17916 36864 17950
rect 36898 17916 36954 17950
rect 36988 17916 37044 17950
rect 37078 17916 37134 17950
rect 37168 17916 37224 17950
rect 37258 17916 37310 17950
rect 36630 17860 37310 17916
rect 36630 17826 36684 17860
rect 36718 17826 36774 17860
rect 36808 17826 36864 17860
rect 36898 17826 36954 17860
rect 36988 17826 37044 17860
rect 37078 17826 37134 17860
rect 37168 17826 37224 17860
rect 37258 17826 37310 17860
rect 36630 17770 37310 17826
rect 36630 17736 36684 17770
rect 36718 17736 36774 17770
rect 36808 17736 36864 17770
rect 36898 17736 36954 17770
rect 36988 17736 37044 17770
rect 37078 17736 37134 17770
rect 37168 17736 37224 17770
rect 37258 17736 37310 17770
rect 36630 17680 37310 17736
rect 36630 17646 36684 17680
rect 36718 17646 36774 17680
rect 36808 17646 36864 17680
rect 36898 17646 36954 17680
rect 36988 17646 37044 17680
rect 37078 17646 37134 17680
rect 37168 17646 37224 17680
rect 37258 17646 37310 17680
rect 36630 17592 37310 17646
rect 37970 18220 38650 18272
rect 37970 18186 38024 18220
rect 38058 18186 38114 18220
rect 38148 18186 38204 18220
rect 38238 18186 38294 18220
rect 38328 18186 38384 18220
rect 38418 18186 38474 18220
rect 38508 18186 38564 18220
rect 38598 18186 38650 18220
rect 37970 18130 38650 18186
rect 37970 18096 38024 18130
rect 38058 18096 38114 18130
rect 38148 18096 38204 18130
rect 38238 18096 38294 18130
rect 38328 18096 38384 18130
rect 38418 18096 38474 18130
rect 38508 18096 38564 18130
rect 38598 18096 38650 18130
rect 37970 18040 38650 18096
rect 37970 18006 38024 18040
rect 38058 18006 38114 18040
rect 38148 18006 38204 18040
rect 38238 18006 38294 18040
rect 38328 18006 38384 18040
rect 38418 18006 38474 18040
rect 38508 18006 38564 18040
rect 38598 18006 38650 18040
rect 37970 17950 38650 18006
rect 37970 17916 38024 17950
rect 38058 17916 38114 17950
rect 38148 17916 38204 17950
rect 38238 17916 38294 17950
rect 38328 17916 38384 17950
rect 38418 17916 38474 17950
rect 38508 17916 38564 17950
rect 38598 17916 38650 17950
rect 37970 17860 38650 17916
rect 37970 17826 38024 17860
rect 38058 17826 38114 17860
rect 38148 17826 38204 17860
rect 38238 17826 38294 17860
rect 38328 17826 38384 17860
rect 38418 17826 38474 17860
rect 38508 17826 38564 17860
rect 38598 17826 38650 17860
rect 37970 17770 38650 17826
rect 37970 17736 38024 17770
rect 38058 17736 38114 17770
rect 38148 17736 38204 17770
rect 38238 17736 38294 17770
rect 38328 17736 38384 17770
rect 38418 17736 38474 17770
rect 38508 17736 38564 17770
rect 38598 17736 38650 17770
rect 37970 17680 38650 17736
rect 37970 17646 38024 17680
rect 38058 17646 38114 17680
rect 38148 17646 38204 17680
rect 38238 17646 38294 17680
rect 38328 17646 38384 17680
rect 38418 17646 38474 17680
rect 38508 17646 38564 17680
rect 38598 17646 38650 17680
rect 37970 17592 38650 17646
rect 28590 14460 29270 14512
rect 28590 14426 28644 14460
rect 28678 14426 28734 14460
rect 28768 14426 28824 14460
rect 28858 14426 28914 14460
rect 28948 14426 29004 14460
rect 29038 14426 29094 14460
rect 29128 14426 29184 14460
rect 29218 14426 29270 14460
rect 28590 14370 29270 14426
rect 28590 14336 28644 14370
rect 28678 14336 28734 14370
rect 28768 14336 28824 14370
rect 28858 14336 28914 14370
rect 28948 14336 29004 14370
rect 29038 14336 29094 14370
rect 29128 14336 29184 14370
rect 29218 14336 29270 14370
rect 28590 14280 29270 14336
rect 28590 14246 28644 14280
rect 28678 14246 28734 14280
rect 28768 14246 28824 14280
rect 28858 14246 28914 14280
rect 28948 14246 29004 14280
rect 29038 14246 29094 14280
rect 29128 14246 29184 14280
rect 29218 14246 29270 14280
rect 28590 14190 29270 14246
rect 28590 14156 28644 14190
rect 28678 14156 28734 14190
rect 28768 14156 28824 14190
rect 28858 14156 28914 14190
rect 28948 14156 29004 14190
rect 29038 14156 29094 14190
rect 29128 14156 29184 14190
rect 29218 14156 29270 14190
rect 28590 14100 29270 14156
rect 28590 14066 28644 14100
rect 28678 14066 28734 14100
rect 28768 14066 28824 14100
rect 28858 14066 28914 14100
rect 28948 14066 29004 14100
rect 29038 14066 29094 14100
rect 29128 14066 29184 14100
rect 29218 14066 29270 14100
rect 28590 14010 29270 14066
rect 28590 13976 28644 14010
rect 28678 13976 28734 14010
rect 28768 13976 28824 14010
rect 28858 13976 28914 14010
rect 28948 13976 29004 14010
rect 29038 13976 29094 14010
rect 29128 13976 29184 14010
rect 29218 13976 29270 14010
rect 28590 13920 29270 13976
rect 28590 13886 28644 13920
rect 28678 13886 28734 13920
rect 28768 13886 28824 13920
rect 28858 13886 28914 13920
rect 28948 13886 29004 13920
rect 29038 13886 29094 13920
rect 29128 13886 29184 13920
rect 29218 13886 29270 13920
rect 28590 13832 29270 13886
rect 29930 14460 30610 14512
rect 29930 14426 29984 14460
rect 30018 14426 30074 14460
rect 30108 14426 30164 14460
rect 30198 14426 30254 14460
rect 30288 14426 30344 14460
rect 30378 14426 30434 14460
rect 30468 14426 30524 14460
rect 30558 14426 30610 14460
rect 29930 14370 30610 14426
rect 29930 14336 29984 14370
rect 30018 14336 30074 14370
rect 30108 14336 30164 14370
rect 30198 14336 30254 14370
rect 30288 14336 30344 14370
rect 30378 14336 30434 14370
rect 30468 14336 30524 14370
rect 30558 14336 30610 14370
rect 29930 14280 30610 14336
rect 29930 14246 29984 14280
rect 30018 14246 30074 14280
rect 30108 14246 30164 14280
rect 30198 14246 30254 14280
rect 30288 14246 30344 14280
rect 30378 14246 30434 14280
rect 30468 14246 30524 14280
rect 30558 14246 30610 14280
rect 29930 14190 30610 14246
rect 29930 14156 29984 14190
rect 30018 14156 30074 14190
rect 30108 14156 30164 14190
rect 30198 14156 30254 14190
rect 30288 14156 30344 14190
rect 30378 14156 30434 14190
rect 30468 14156 30524 14190
rect 30558 14156 30610 14190
rect 29930 14100 30610 14156
rect 29930 14066 29984 14100
rect 30018 14066 30074 14100
rect 30108 14066 30164 14100
rect 30198 14066 30254 14100
rect 30288 14066 30344 14100
rect 30378 14066 30434 14100
rect 30468 14066 30524 14100
rect 30558 14066 30610 14100
rect 29930 14010 30610 14066
rect 29930 13976 29984 14010
rect 30018 13976 30074 14010
rect 30108 13976 30164 14010
rect 30198 13976 30254 14010
rect 30288 13976 30344 14010
rect 30378 13976 30434 14010
rect 30468 13976 30524 14010
rect 30558 13976 30610 14010
rect 29930 13920 30610 13976
rect 29930 13886 29984 13920
rect 30018 13886 30074 13920
rect 30108 13886 30164 13920
rect 30198 13886 30254 13920
rect 30288 13886 30344 13920
rect 30378 13886 30434 13920
rect 30468 13886 30524 13920
rect 30558 13886 30610 13920
rect 29930 13832 30610 13886
rect 31270 14460 31950 14512
rect 31270 14426 31324 14460
rect 31358 14426 31414 14460
rect 31448 14426 31504 14460
rect 31538 14426 31594 14460
rect 31628 14426 31684 14460
rect 31718 14426 31774 14460
rect 31808 14426 31864 14460
rect 31898 14426 31950 14460
rect 31270 14370 31950 14426
rect 31270 14336 31324 14370
rect 31358 14336 31414 14370
rect 31448 14336 31504 14370
rect 31538 14336 31594 14370
rect 31628 14336 31684 14370
rect 31718 14336 31774 14370
rect 31808 14336 31864 14370
rect 31898 14336 31950 14370
rect 31270 14280 31950 14336
rect 31270 14246 31324 14280
rect 31358 14246 31414 14280
rect 31448 14246 31504 14280
rect 31538 14246 31594 14280
rect 31628 14246 31684 14280
rect 31718 14246 31774 14280
rect 31808 14246 31864 14280
rect 31898 14246 31950 14280
rect 31270 14190 31950 14246
rect 31270 14156 31324 14190
rect 31358 14156 31414 14190
rect 31448 14156 31504 14190
rect 31538 14156 31594 14190
rect 31628 14156 31684 14190
rect 31718 14156 31774 14190
rect 31808 14156 31864 14190
rect 31898 14156 31950 14190
rect 31270 14100 31950 14156
rect 31270 14066 31324 14100
rect 31358 14066 31414 14100
rect 31448 14066 31504 14100
rect 31538 14066 31594 14100
rect 31628 14066 31684 14100
rect 31718 14066 31774 14100
rect 31808 14066 31864 14100
rect 31898 14066 31950 14100
rect 31270 14010 31950 14066
rect 31270 13976 31324 14010
rect 31358 13976 31414 14010
rect 31448 13976 31504 14010
rect 31538 13976 31594 14010
rect 31628 13976 31684 14010
rect 31718 13976 31774 14010
rect 31808 13976 31864 14010
rect 31898 13976 31950 14010
rect 31270 13920 31950 13976
rect 31270 13886 31324 13920
rect 31358 13886 31414 13920
rect 31448 13886 31504 13920
rect 31538 13886 31594 13920
rect 31628 13886 31684 13920
rect 31718 13886 31774 13920
rect 31808 13886 31864 13920
rect 31898 13886 31950 13920
rect 31270 13832 31950 13886
rect 32610 14460 33290 14512
rect 32610 14426 32664 14460
rect 32698 14426 32754 14460
rect 32788 14426 32844 14460
rect 32878 14426 32934 14460
rect 32968 14426 33024 14460
rect 33058 14426 33114 14460
rect 33148 14426 33204 14460
rect 33238 14426 33290 14460
rect 32610 14370 33290 14426
rect 32610 14336 32664 14370
rect 32698 14336 32754 14370
rect 32788 14336 32844 14370
rect 32878 14336 32934 14370
rect 32968 14336 33024 14370
rect 33058 14336 33114 14370
rect 33148 14336 33204 14370
rect 33238 14336 33290 14370
rect 32610 14280 33290 14336
rect 32610 14246 32664 14280
rect 32698 14246 32754 14280
rect 32788 14246 32844 14280
rect 32878 14246 32934 14280
rect 32968 14246 33024 14280
rect 33058 14246 33114 14280
rect 33148 14246 33204 14280
rect 33238 14246 33290 14280
rect 32610 14190 33290 14246
rect 32610 14156 32664 14190
rect 32698 14156 32754 14190
rect 32788 14156 32844 14190
rect 32878 14156 32934 14190
rect 32968 14156 33024 14190
rect 33058 14156 33114 14190
rect 33148 14156 33204 14190
rect 33238 14156 33290 14190
rect 32610 14100 33290 14156
rect 32610 14066 32664 14100
rect 32698 14066 32754 14100
rect 32788 14066 32844 14100
rect 32878 14066 32934 14100
rect 32968 14066 33024 14100
rect 33058 14066 33114 14100
rect 33148 14066 33204 14100
rect 33238 14066 33290 14100
rect 32610 14010 33290 14066
rect 32610 13976 32664 14010
rect 32698 13976 32754 14010
rect 32788 13976 32844 14010
rect 32878 13976 32934 14010
rect 32968 13976 33024 14010
rect 33058 13976 33114 14010
rect 33148 13976 33204 14010
rect 33238 13976 33290 14010
rect 32610 13920 33290 13976
rect 32610 13886 32664 13920
rect 32698 13886 32754 13920
rect 32788 13886 32844 13920
rect 32878 13886 32934 13920
rect 32968 13886 33024 13920
rect 33058 13886 33114 13920
rect 33148 13886 33204 13920
rect 33238 13886 33290 13920
rect 32610 13832 33290 13886
rect 33950 14460 34630 14512
rect 33950 14426 34004 14460
rect 34038 14426 34094 14460
rect 34128 14426 34184 14460
rect 34218 14426 34274 14460
rect 34308 14426 34364 14460
rect 34398 14426 34454 14460
rect 34488 14426 34544 14460
rect 34578 14426 34630 14460
rect 33950 14370 34630 14426
rect 33950 14336 34004 14370
rect 34038 14336 34094 14370
rect 34128 14336 34184 14370
rect 34218 14336 34274 14370
rect 34308 14336 34364 14370
rect 34398 14336 34454 14370
rect 34488 14336 34544 14370
rect 34578 14336 34630 14370
rect 33950 14280 34630 14336
rect 33950 14246 34004 14280
rect 34038 14246 34094 14280
rect 34128 14246 34184 14280
rect 34218 14246 34274 14280
rect 34308 14246 34364 14280
rect 34398 14246 34454 14280
rect 34488 14246 34544 14280
rect 34578 14246 34630 14280
rect 33950 14190 34630 14246
rect 33950 14156 34004 14190
rect 34038 14156 34094 14190
rect 34128 14156 34184 14190
rect 34218 14156 34274 14190
rect 34308 14156 34364 14190
rect 34398 14156 34454 14190
rect 34488 14156 34544 14190
rect 34578 14156 34630 14190
rect 33950 14100 34630 14156
rect 33950 14066 34004 14100
rect 34038 14066 34094 14100
rect 34128 14066 34184 14100
rect 34218 14066 34274 14100
rect 34308 14066 34364 14100
rect 34398 14066 34454 14100
rect 34488 14066 34544 14100
rect 34578 14066 34630 14100
rect 33950 14010 34630 14066
rect 33950 13976 34004 14010
rect 34038 13976 34094 14010
rect 34128 13976 34184 14010
rect 34218 13976 34274 14010
rect 34308 13976 34364 14010
rect 34398 13976 34454 14010
rect 34488 13976 34544 14010
rect 34578 13976 34630 14010
rect 33950 13920 34630 13976
rect 33950 13886 34004 13920
rect 34038 13886 34094 13920
rect 34128 13886 34184 13920
rect 34218 13886 34274 13920
rect 34308 13886 34364 13920
rect 34398 13886 34454 13920
rect 34488 13886 34544 13920
rect 34578 13886 34630 13920
rect 33950 13832 34630 13886
rect 35290 14460 35970 14512
rect 35290 14426 35344 14460
rect 35378 14426 35434 14460
rect 35468 14426 35524 14460
rect 35558 14426 35614 14460
rect 35648 14426 35704 14460
rect 35738 14426 35794 14460
rect 35828 14426 35884 14460
rect 35918 14426 35970 14460
rect 35290 14370 35970 14426
rect 35290 14336 35344 14370
rect 35378 14336 35434 14370
rect 35468 14336 35524 14370
rect 35558 14336 35614 14370
rect 35648 14336 35704 14370
rect 35738 14336 35794 14370
rect 35828 14336 35884 14370
rect 35918 14336 35970 14370
rect 35290 14280 35970 14336
rect 35290 14246 35344 14280
rect 35378 14246 35434 14280
rect 35468 14246 35524 14280
rect 35558 14246 35614 14280
rect 35648 14246 35704 14280
rect 35738 14246 35794 14280
rect 35828 14246 35884 14280
rect 35918 14246 35970 14280
rect 35290 14190 35970 14246
rect 35290 14156 35344 14190
rect 35378 14156 35434 14190
rect 35468 14156 35524 14190
rect 35558 14156 35614 14190
rect 35648 14156 35704 14190
rect 35738 14156 35794 14190
rect 35828 14156 35884 14190
rect 35918 14156 35970 14190
rect 35290 14100 35970 14156
rect 35290 14066 35344 14100
rect 35378 14066 35434 14100
rect 35468 14066 35524 14100
rect 35558 14066 35614 14100
rect 35648 14066 35704 14100
rect 35738 14066 35794 14100
rect 35828 14066 35884 14100
rect 35918 14066 35970 14100
rect 35290 14010 35970 14066
rect 35290 13976 35344 14010
rect 35378 13976 35434 14010
rect 35468 13976 35524 14010
rect 35558 13976 35614 14010
rect 35648 13976 35704 14010
rect 35738 13976 35794 14010
rect 35828 13976 35884 14010
rect 35918 13976 35970 14010
rect 35290 13920 35970 13976
rect 35290 13886 35344 13920
rect 35378 13886 35434 13920
rect 35468 13886 35524 13920
rect 35558 13886 35614 13920
rect 35648 13886 35704 13920
rect 35738 13886 35794 13920
rect 35828 13886 35884 13920
rect 35918 13886 35970 13920
rect 35290 13832 35970 13886
rect 36630 14460 37310 14512
rect 36630 14426 36684 14460
rect 36718 14426 36774 14460
rect 36808 14426 36864 14460
rect 36898 14426 36954 14460
rect 36988 14426 37044 14460
rect 37078 14426 37134 14460
rect 37168 14426 37224 14460
rect 37258 14426 37310 14460
rect 36630 14370 37310 14426
rect 36630 14336 36684 14370
rect 36718 14336 36774 14370
rect 36808 14336 36864 14370
rect 36898 14336 36954 14370
rect 36988 14336 37044 14370
rect 37078 14336 37134 14370
rect 37168 14336 37224 14370
rect 37258 14336 37310 14370
rect 36630 14280 37310 14336
rect 36630 14246 36684 14280
rect 36718 14246 36774 14280
rect 36808 14246 36864 14280
rect 36898 14246 36954 14280
rect 36988 14246 37044 14280
rect 37078 14246 37134 14280
rect 37168 14246 37224 14280
rect 37258 14246 37310 14280
rect 36630 14190 37310 14246
rect 36630 14156 36684 14190
rect 36718 14156 36774 14190
rect 36808 14156 36864 14190
rect 36898 14156 36954 14190
rect 36988 14156 37044 14190
rect 37078 14156 37134 14190
rect 37168 14156 37224 14190
rect 37258 14156 37310 14190
rect 36630 14100 37310 14156
rect 36630 14066 36684 14100
rect 36718 14066 36774 14100
rect 36808 14066 36864 14100
rect 36898 14066 36954 14100
rect 36988 14066 37044 14100
rect 37078 14066 37134 14100
rect 37168 14066 37224 14100
rect 37258 14066 37310 14100
rect 36630 14010 37310 14066
rect 36630 13976 36684 14010
rect 36718 13976 36774 14010
rect 36808 13976 36864 14010
rect 36898 13976 36954 14010
rect 36988 13976 37044 14010
rect 37078 13976 37134 14010
rect 37168 13976 37224 14010
rect 37258 13976 37310 14010
rect 36630 13920 37310 13976
rect 36630 13886 36684 13920
rect 36718 13886 36774 13920
rect 36808 13886 36864 13920
rect 36898 13886 36954 13920
rect 36988 13886 37044 13920
rect 37078 13886 37134 13920
rect 37168 13886 37224 13920
rect 37258 13886 37310 13920
rect 36630 13832 37310 13886
rect 37970 14460 38650 14512
rect 37970 14426 38024 14460
rect 38058 14426 38114 14460
rect 38148 14426 38204 14460
rect 38238 14426 38294 14460
rect 38328 14426 38384 14460
rect 38418 14426 38474 14460
rect 38508 14426 38564 14460
rect 38598 14426 38650 14460
rect 37970 14370 38650 14426
rect 37970 14336 38024 14370
rect 38058 14336 38114 14370
rect 38148 14336 38204 14370
rect 38238 14336 38294 14370
rect 38328 14336 38384 14370
rect 38418 14336 38474 14370
rect 38508 14336 38564 14370
rect 38598 14336 38650 14370
rect 37970 14280 38650 14336
rect 37970 14246 38024 14280
rect 38058 14246 38114 14280
rect 38148 14246 38204 14280
rect 38238 14246 38294 14280
rect 38328 14246 38384 14280
rect 38418 14246 38474 14280
rect 38508 14246 38564 14280
rect 38598 14246 38650 14280
rect 37970 14190 38650 14246
rect 37970 14156 38024 14190
rect 38058 14156 38114 14190
rect 38148 14156 38204 14190
rect 38238 14156 38294 14190
rect 38328 14156 38384 14190
rect 38418 14156 38474 14190
rect 38508 14156 38564 14190
rect 38598 14156 38650 14190
rect 37970 14100 38650 14156
rect 37970 14066 38024 14100
rect 38058 14066 38114 14100
rect 38148 14066 38204 14100
rect 38238 14066 38294 14100
rect 38328 14066 38384 14100
rect 38418 14066 38474 14100
rect 38508 14066 38564 14100
rect 38598 14066 38650 14100
rect 37970 14010 38650 14066
rect 37970 13976 38024 14010
rect 38058 13976 38114 14010
rect 38148 13976 38204 14010
rect 38238 13976 38294 14010
rect 38328 13976 38384 14010
rect 38418 13976 38474 14010
rect 38508 13976 38564 14010
rect 38598 13976 38650 14010
rect 37970 13920 38650 13976
rect 37970 13886 38024 13920
rect 38058 13886 38114 13920
rect 38148 13886 38204 13920
rect 38238 13886 38294 13920
rect 38328 13886 38384 13920
rect 38418 13886 38474 13920
rect 38508 13886 38564 13920
rect 38598 13886 38650 13920
rect 37970 13832 38650 13886
<< ndiffc >>
rect 5996 40875 6030 40909
rect 5996 40807 6030 40841
rect 5996 40739 6030 40773
rect 5996 40671 6030 40705
rect 5996 40603 6030 40637
rect 5996 40535 6030 40569
rect 5996 40467 6030 40501
rect 5996 40399 6030 40433
rect 5996 40331 6030 40365
rect 5996 40263 6030 40297
rect 5996 40195 6030 40229
rect 6454 40875 6488 40909
rect 6454 40807 6488 40841
rect 6454 40739 6488 40773
rect 6454 40671 6488 40705
rect 6454 40603 6488 40637
rect 6454 40535 6488 40569
rect 6454 40467 6488 40501
rect 6454 40399 6488 40433
rect 6454 40331 6488 40365
rect 6454 40263 6488 40297
rect 6454 40195 6488 40229
rect 28340 37115 28374 37149
rect 28340 37047 28374 37081
rect 28340 36979 28374 37013
rect 28340 36911 28374 36945
rect 28340 36843 28374 36877
rect 28340 36775 28374 36809
rect 28340 36707 28374 36741
rect 28340 36639 28374 36673
rect 28340 36571 28374 36605
rect 28340 36503 28374 36537
rect 28340 36435 28374 36469
rect 28798 37115 28832 37149
rect 28798 37047 28832 37081
rect 28798 36979 28832 37013
rect 28798 36911 28832 36945
rect 28798 36843 28832 36877
rect 28798 36775 28832 36809
rect 28798 36707 28832 36741
rect 28798 36639 28832 36673
rect 28798 36571 28832 36605
rect 28798 36503 28832 36537
rect 28798 36435 28832 36469
rect 22980 25835 23014 25869
rect 22980 25767 23014 25801
rect 22980 25699 23014 25733
rect 22980 25631 23014 25665
rect 22980 25563 23014 25597
rect 22980 25495 23014 25529
rect 22980 25427 23014 25461
rect 22980 25359 23014 25393
rect 22980 25291 23014 25325
rect 22980 25223 23014 25257
rect 22980 25155 23014 25189
rect 23438 25835 23472 25869
rect 23438 25767 23472 25801
rect 23438 25699 23472 25733
rect 23438 25631 23472 25665
rect 23438 25563 23472 25597
rect 23438 25495 23472 25529
rect 23438 25427 23472 25461
rect 23438 25359 23472 25393
rect 23438 25291 23472 25325
rect 23438 25223 23472 25257
rect 23438 25155 23472 25189
rect 23896 25835 23930 25869
rect 23896 25767 23930 25801
rect 23896 25699 23930 25733
rect 23896 25631 23930 25665
rect 23896 25563 23930 25597
rect 23896 25495 23930 25529
rect 23896 25427 23930 25461
rect 23896 25359 23930 25393
rect 23896 25291 23930 25325
rect 23896 25223 23930 25257
rect 23896 25155 23930 25189
rect 24354 25835 24388 25869
rect 24354 25767 24388 25801
rect 24354 25699 24388 25733
rect 24354 25631 24388 25665
rect 24354 25563 24388 25597
rect 24354 25495 24388 25529
rect 24354 25427 24388 25461
rect 24354 25359 24388 25393
rect 24354 25291 24388 25325
rect 24354 25223 24388 25257
rect 24354 25155 24388 25189
rect 24812 25835 24846 25869
rect 24812 25767 24846 25801
rect 24812 25699 24846 25733
rect 24812 25631 24846 25665
rect 24812 25563 24846 25597
rect 24812 25495 24846 25529
rect 24812 25427 24846 25461
rect 24812 25359 24846 25393
rect 24812 25291 24846 25325
rect 24812 25223 24846 25257
rect 24812 25155 24846 25189
rect 25270 25835 25304 25869
rect 25270 25767 25304 25801
rect 25270 25699 25304 25733
rect 25270 25631 25304 25665
rect 25270 25563 25304 25597
rect 25270 25495 25304 25529
rect 25270 25427 25304 25461
rect 25270 25359 25304 25393
rect 25270 25291 25304 25325
rect 25270 25223 25304 25257
rect 25270 25155 25304 25189
rect 25728 25835 25762 25869
rect 25728 25767 25762 25801
rect 25728 25699 25762 25733
rect 25728 25631 25762 25665
rect 25728 25563 25762 25597
rect 25728 25495 25762 25529
rect 25728 25427 25762 25461
rect 25728 25359 25762 25393
rect 25728 25291 25762 25325
rect 25728 25223 25762 25257
rect 25728 25155 25762 25189
rect 26186 25835 26220 25869
rect 26186 25767 26220 25801
rect 26186 25699 26220 25733
rect 26186 25631 26220 25665
rect 26186 25563 26220 25597
rect 26186 25495 26220 25529
rect 26186 25427 26220 25461
rect 26186 25359 26220 25393
rect 26186 25291 26220 25325
rect 26186 25223 26220 25257
rect 26186 25155 26220 25189
rect 26644 25835 26678 25869
rect 26644 25767 26678 25801
rect 26644 25699 26678 25733
rect 26644 25631 26678 25665
rect 26644 25563 26678 25597
rect 26644 25495 26678 25529
rect 26644 25427 26678 25461
rect 26644 25359 26678 25393
rect 26644 25291 26678 25325
rect 26644 25223 26678 25257
rect 26644 25155 26678 25189
rect 27102 25835 27136 25869
rect 27102 25767 27136 25801
rect 27102 25699 27136 25733
rect 27102 25631 27136 25665
rect 27102 25563 27136 25597
rect 27102 25495 27136 25529
rect 27102 25427 27136 25461
rect 27102 25359 27136 25393
rect 27102 25291 27136 25325
rect 27102 25223 27136 25257
rect 27102 25155 27136 25189
rect 22980 22075 23014 22109
rect 22980 22007 23014 22041
rect 22980 21939 23014 21973
rect 22980 21871 23014 21905
rect 22980 21803 23014 21837
rect 22980 21735 23014 21769
rect 22980 21667 23014 21701
rect 22980 21599 23014 21633
rect 22980 21531 23014 21565
rect 22980 21463 23014 21497
rect 22980 21395 23014 21429
rect 23438 22075 23472 22109
rect 23438 22007 23472 22041
rect 23438 21939 23472 21973
rect 23438 21871 23472 21905
rect 23438 21803 23472 21837
rect 23438 21735 23472 21769
rect 23438 21667 23472 21701
rect 23438 21599 23472 21633
rect 23438 21531 23472 21565
rect 23438 21463 23472 21497
rect 23438 21395 23472 21429
rect 23896 22075 23930 22109
rect 23896 22007 23930 22041
rect 23896 21939 23930 21973
rect 23896 21871 23930 21905
rect 23896 21803 23930 21837
rect 23896 21735 23930 21769
rect 23896 21667 23930 21701
rect 23896 21599 23930 21633
rect 23896 21531 23930 21565
rect 23896 21463 23930 21497
rect 23896 21395 23930 21429
rect 24354 22075 24388 22109
rect 24354 22007 24388 22041
rect 24354 21939 24388 21973
rect 24354 21871 24388 21905
rect 24354 21803 24388 21837
rect 24354 21735 24388 21769
rect 24354 21667 24388 21701
rect 24354 21599 24388 21633
rect 24354 21531 24388 21565
rect 24354 21463 24388 21497
rect 24354 21395 24388 21429
rect 24812 22075 24846 22109
rect 24812 22007 24846 22041
rect 24812 21939 24846 21973
rect 24812 21871 24846 21905
rect 24812 21803 24846 21837
rect 24812 21735 24846 21769
rect 24812 21667 24846 21701
rect 24812 21599 24846 21633
rect 24812 21531 24846 21565
rect 24812 21463 24846 21497
rect 24812 21395 24846 21429
rect 25270 22075 25304 22109
rect 25270 22007 25304 22041
rect 25270 21939 25304 21973
rect 25270 21871 25304 21905
rect 25270 21803 25304 21837
rect 25270 21735 25304 21769
rect 25270 21667 25304 21701
rect 25270 21599 25304 21633
rect 25270 21531 25304 21565
rect 25270 21463 25304 21497
rect 25270 21395 25304 21429
rect 25728 22075 25762 22109
rect 25728 22007 25762 22041
rect 25728 21939 25762 21973
rect 25728 21871 25762 21905
rect 25728 21803 25762 21837
rect 25728 21735 25762 21769
rect 25728 21667 25762 21701
rect 25728 21599 25762 21633
rect 25728 21531 25762 21565
rect 25728 21463 25762 21497
rect 25728 21395 25762 21429
rect 26186 22075 26220 22109
rect 26186 22007 26220 22041
rect 26186 21939 26220 21973
rect 26186 21871 26220 21905
rect 26186 21803 26220 21837
rect 26186 21735 26220 21769
rect 26186 21667 26220 21701
rect 26186 21599 26220 21633
rect 26186 21531 26220 21565
rect 26186 21463 26220 21497
rect 26186 21395 26220 21429
rect 26644 22075 26678 22109
rect 26644 22007 26678 22041
rect 26644 21939 26678 21973
rect 26644 21871 26678 21905
rect 26644 21803 26678 21837
rect 26644 21735 26678 21769
rect 26644 21667 26678 21701
rect 26644 21599 26678 21633
rect 26644 21531 26678 21565
rect 26644 21463 26678 21497
rect 26644 21395 26678 21429
rect 27102 22075 27136 22109
rect 27102 22007 27136 22041
rect 27102 21939 27136 21973
rect 27102 21871 27136 21905
rect 27102 21803 27136 21837
rect 27102 21735 27136 21769
rect 27102 21667 27136 21701
rect 27102 21599 27136 21633
rect 27102 21531 27136 21565
rect 27102 21463 27136 21497
rect 27102 21395 27136 21429
rect 6026 18315 6060 18349
rect 6026 18247 6060 18281
rect 6026 18179 6060 18213
rect 6026 18111 6060 18145
rect 6026 18043 6060 18077
rect 6026 17975 6060 18009
rect 6026 17907 6060 17941
rect 6026 17839 6060 17873
rect 6026 17771 6060 17805
rect 6026 17703 6060 17737
rect 6026 17635 6060 17669
rect 6484 18315 6518 18349
rect 6484 18247 6518 18281
rect 6484 18179 6518 18213
rect 6484 18111 6518 18145
rect 6484 18043 6518 18077
rect 6484 17975 6518 18009
rect 6484 17907 6518 17941
rect 6484 17839 6518 17873
rect 6484 17771 6518 17805
rect 6484 17703 6518 17737
rect 6484 17635 6518 17669
rect 6942 18315 6976 18349
rect 6942 18247 6976 18281
rect 6942 18179 6976 18213
rect 6942 18111 6976 18145
rect 6942 18043 6976 18077
rect 6942 17975 6976 18009
rect 6942 17907 6976 17941
rect 6942 17839 6976 17873
rect 6942 17771 6976 17805
rect 6942 17703 6976 17737
rect 6942 17635 6976 17669
rect 7400 18315 7434 18349
rect 7400 18247 7434 18281
rect 7400 18179 7434 18213
rect 7400 18111 7434 18145
rect 7400 18043 7434 18077
rect 7400 17975 7434 18009
rect 7400 17907 7434 17941
rect 7400 17839 7434 17873
rect 7400 17771 7434 17805
rect 7400 17703 7434 17737
rect 7400 17635 7434 17669
rect 7858 18315 7892 18349
rect 7858 18247 7892 18281
rect 7858 18179 7892 18213
rect 7858 18111 7892 18145
rect 7858 18043 7892 18077
rect 7858 17975 7892 18009
rect 7858 17907 7892 17941
rect 7858 17839 7892 17873
rect 7858 17771 7892 17805
rect 7858 17703 7892 17737
rect 7858 17635 7892 17669
rect 8316 18315 8350 18349
rect 8316 18247 8350 18281
rect 8316 18179 8350 18213
rect 8316 18111 8350 18145
rect 8316 18043 8350 18077
rect 8316 17975 8350 18009
rect 8316 17907 8350 17941
rect 8316 17839 8350 17873
rect 8316 17771 8350 17805
rect 8316 17703 8350 17737
rect 8316 17635 8350 17669
rect 8774 18315 8808 18349
rect 8774 18247 8808 18281
rect 8774 18179 8808 18213
rect 8774 18111 8808 18145
rect 8774 18043 8808 18077
rect 8774 17975 8808 18009
rect 8774 17907 8808 17941
rect 8774 17839 8808 17873
rect 8774 17771 8808 17805
rect 8774 17703 8808 17737
rect 8774 17635 8808 17669
rect 9232 18315 9266 18349
rect 9232 18247 9266 18281
rect 9232 18179 9266 18213
rect 9232 18111 9266 18145
rect 9232 18043 9266 18077
rect 9232 17975 9266 18009
rect 9232 17907 9266 17941
rect 9232 17839 9266 17873
rect 9232 17771 9266 17805
rect 9232 17703 9266 17737
rect 9232 17635 9266 17669
rect 9690 18315 9724 18349
rect 9690 18247 9724 18281
rect 9690 18179 9724 18213
rect 9690 18111 9724 18145
rect 9690 18043 9724 18077
rect 9690 17975 9724 18009
rect 9690 17907 9724 17941
rect 9690 17839 9724 17873
rect 9690 17771 9724 17805
rect 9690 17703 9724 17737
rect 9690 17635 9724 17669
rect 10148 18315 10182 18349
rect 10148 18247 10182 18281
rect 10148 18179 10182 18213
rect 10148 18111 10182 18145
rect 10148 18043 10182 18077
rect 10148 17975 10182 18009
rect 10148 17907 10182 17941
rect 10148 17839 10182 17873
rect 10148 17771 10182 17805
rect 10148 17703 10182 17737
rect 10148 17635 10182 17669
<< pdiffc >>
rect 15077 41147 15111 41181
rect 15077 41079 15111 41113
rect 15077 41011 15111 41045
rect 15077 40943 15111 40977
rect 15077 40875 15111 40909
rect 15077 40807 15111 40841
rect 15077 40739 15111 40773
rect 15077 40671 15111 40705
rect 15077 40603 15111 40637
rect 15077 40535 15111 40569
rect 15077 40467 15111 40501
rect 15077 40399 15111 40433
rect 15077 40331 15111 40365
rect 15077 40263 15111 40297
rect 15077 40195 15111 40229
rect 15077 40127 15111 40161
rect 15077 40059 15111 40093
rect 15077 39991 15111 40025
rect 15077 39923 15111 39957
rect 15535 41147 15569 41181
rect 15535 41079 15569 41113
rect 15535 41011 15569 41045
rect 15535 40943 15569 40977
rect 15535 40875 15569 40909
rect 15535 40807 15569 40841
rect 15535 40739 15569 40773
rect 15535 40671 15569 40705
rect 15535 40603 15569 40637
rect 15535 40535 15569 40569
rect 15535 40467 15569 40501
rect 15535 40399 15569 40433
rect 15535 40331 15569 40365
rect 15535 40263 15569 40297
rect 15535 40195 15569 40229
rect 15535 40127 15569 40161
rect 15535 40059 15569 40093
rect 15535 39991 15569 40025
rect 15535 39923 15569 39957
rect 15993 41147 16027 41181
rect 15993 41079 16027 41113
rect 15993 41011 16027 41045
rect 15993 40943 16027 40977
rect 15993 40875 16027 40909
rect 15993 40807 16027 40841
rect 15993 40739 16027 40773
rect 15993 40671 16027 40705
rect 15993 40603 16027 40637
rect 15993 40535 16027 40569
rect 15993 40467 16027 40501
rect 15993 40399 16027 40433
rect 15993 40331 16027 40365
rect 15993 40263 16027 40297
rect 15993 40195 16027 40229
rect 15993 40127 16027 40161
rect 15993 40059 16027 40093
rect 15993 39991 16027 40025
rect 15993 39923 16027 39957
rect 16451 41147 16485 41181
rect 16451 41079 16485 41113
rect 16451 41011 16485 41045
rect 16451 40943 16485 40977
rect 16451 40875 16485 40909
rect 16451 40807 16485 40841
rect 16451 40739 16485 40773
rect 16451 40671 16485 40705
rect 16451 40603 16485 40637
rect 16451 40535 16485 40569
rect 16451 40467 16485 40501
rect 16451 40399 16485 40433
rect 16451 40331 16485 40365
rect 16451 40263 16485 40297
rect 16451 40195 16485 40229
rect 16451 40127 16485 40161
rect 16451 40059 16485 40093
rect 16451 39991 16485 40025
rect 16451 39923 16485 39957
rect 16909 41147 16943 41181
rect 16909 41079 16943 41113
rect 16909 41011 16943 41045
rect 16909 40943 16943 40977
rect 16909 40875 16943 40909
rect 16909 40807 16943 40841
rect 16909 40739 16943 40773
rect 16909 40671 16943 40705
rect 16909 40603 16943 40637
rect 16909 40535 16943 40569
rect 16909 40467 16943 40501
rect 16909 40399 16943 40433
rect 16909 40331 16943 40365
rect 16909 40263 16943 40297
rect 16909 40195 16943 40229
rect 16909 40127 16943 40161
rect 16909 40059 16943 40093
rect 16909 39991 16943 40025
rect 16909 39923 16943 39957
rect 17367 41147 17401 41181
rect 17367 41079 17401 41113
rect 17367 41011 17401 41045
rect 17367 40943 17401 40977
rect 17367 40875 17401 40909
rect 17367 40807 17401 40841
rect 17367 40739 17401 40773
rect 17367 40671 17401 40705
rect 17367 40603 17401 40637
rect 17367 40535 17401 40569
rect 17367 40467 17401 40501
rect 17367 40399 17401 40433
rect 17367 40331 17401 40365
rect 17367 40263 17401 40297
rect 17367 40195 17401 40229
rect 17367 40127 17401 40161
rect 17367 40059 17401 40093
rect 17367 39991 17401 40025
rect 17367 39923 17401 39957
rect 17825 41147 17859 41181
rect 17825 41079 17859 41113
rect 17825 41011 17859 41045
rect 17825 40943 17859 40977
rect 17825 40875 17859 40909
rect 17825 40807 17859 40841
rect 17825 40739 17859 40773
rect 17825 40671 17859 40705
rect 17825 40603 17859 40637
rect 17825 40535 17859 40569
rect 17825 40467 17859 40501
rect 17825 40399 17859 40433
rect 17825 40331 17859 40365
rect 17825 40263 17859 40297
rect 17825 40195 17859 40229
rect 17825 40127 17859 40161
rect 17825 40059 17859 40093
rect 17825 39991 17859 40025
rect 17825 39923 17859 39957
rect 18283 41147 18317 41181
rect 18283 41079 18317 41113
rect 18283 41011 18317 41045
rect 18283 40943 18317 40977
rect 18283 40875 18317 40909
rect 18283 40807 18317 40841
rect 18283 40739 18317 40773
rect 18283 40671 18317 40705
rect 18283 40603 18317 40637
rect 18283 40535 18317 40569
rect 18283 40467 18317 40501
rect 18283 40399 18317 40433
rect 18283 40331 18317 40365
rect 18283 40263 18317 40297
rect 18283 40195 18317 40229
rect 18283 40127 18317 40161
rect 18283 40059 18317 40093
rect 18283 39991 18317 40025
rect 18283 39923 18317 39957
rect 18741 41147 18775 41181
rect 18741 41079 18775 41113
rect 18741 41011 18775 41045
rect 18741 40943 18775 40977
rect 18741 40875 18775 40909
rect 18741 40807 18775 40841
rect 18741 40739 18775 40773
rect 18741 40671 18775 40705
rect 18741 40603 18775 40637
rect 18741 40535 18775 40569
rect 18741 40467 18775 40501
rect 18741 40399 18775 40433
rect 18741 40331 18775 40365
rect 18741 40263 18775 40297
rect 18741 40195 18775 40229
rect 18741 40127 18775 40161
rect 18741 40059 18775 40093
rect 18741 39991 18775 40025
rect 18741 39923 18775 39957
rect 19199 41147 19233 41181
rect 19199 41079 19233 41113
rect 19199 41011 19233 41045
rect 19199 40943 19233 40977
rect 19199 40875 19233 40909
rect 19199 40807 19233 40841
rect 19199 40739 19233 40773
rect 19199 40671 19233 40705
rect 19199 40603 19233 40637
rect 19199 40535 19233 40569
rect 19199 40467 19233 40501
rect 19199 40399 19233 40433
rect 19199 40331 19233 40365
rect 19199 40263 19233 40297
rect 19199 40195 19233 40229
rect 19199 40127 19233 40161
rect 19199 40059 19233 40093
rect 19199 39991 19233 40025
rect 19199 39923 19233 39957
rect 19657 41147 19691 41181
rect 19657 41079 19691 41113
rect 19657 41011 19691 41045
rect 19657 40943 19691 40977
rect 19657 40875 19691 40909
rect 19657 40807 19691 40841
rect 19657 40739 19691 40773
rect 19657 40671 19691 40705
rect 19657 40603 19691 40637
rect 19657 40535 19691 40569
rect 19657 40467 19691 40501
rect 19657 40399 19691 40433
rect 19657 40331 19691 40365
rect 19657 40263 19691 40297
rect 19657 40195 19691 40229
rect 19657 40127 19691 40161
rect 19657 40059 19691 40093
rect 19657 39991 19691 40025
rect 19657 39923 19691 39957
rect 20115 41147 20149 41181
rect 20115 41079 20149 41113
rect 20115 41011 20149 41045
rect 20115 40943 20149 40977
rect 20115 40875 20149 40909
rect 20115 40807 20149 40841
rect 20115 40739 20149 40773
rect 20115 40671 20149 40705
rect 20115 40603 20149 40637
rect 20115 40535 20149 40569
rect 20115 40467 20149 40501
rect 20115 40399 20149 40433
rect 20115 40331 20149 40365
rect 20115 40263 20149 40297
rect 20115 40195 20149 40229
rect 20115 40127 20149 40161
rect 20115 40059 20149 40093
rect 20115 39991 20149 40025
rect 20115 39923 20149 39957
rect 20573 41147 20607 41181
rect 20573 41079 20607 41113
rect 20573 41011 20607 41045
rect 20573 40943 20607 40977
rect 20573 40875 20607 40909
rect 20573 40807 20607 40841
rect 20573 40739 20607 40773
rect 20573 40671 20607 40705
rect 20573 40603 20607 40637
rect 20573 40535 20607 40569
rect 20573 40467 20607 40501
rect 20573 40399 20607 40433
rect 20573 40331 20607 40365
rect 20573 40263 20607 40297
rect 20573 40195 20607 40229
rect 20573 40127 20607 40161
rect 20573 40059 20607 40093
rect 20573 39991 20607 40025
rect 20573 39923 20607 39957
rect 21031 41147 21065 41181
rect 21031 41079 21065 41113
rect 21031 41011 21065 41045
rect 21031 40943 21065 40977
rect 21031 40875 21065 40909
rect 21031 40807 21065 40841
rect 21031 40739 21065 40773
rect 21031 40671 21065 40705
rect 21031 40603 21065 40637
rect 21031 40535 21065 40569
rect 21031 40467 21065 40501
rect 21031 40399 21065 40433
rect 21031 40331 21065 40365
rect 21031 40263 21065 40297
rect 21031 40195 21065 40229
rect 21031 40127 21065 40161
rect 21031 40059 21065 40093
rect 21031 39991 21065 40025
rect 21031 39923 21065 39957
rect 21489 41147 21523 41181
rect 21489 41079 21523 41113
rect 21489 41011 21523 41045
rect 21489 40943 21523 40977
rect 21489 40875 21523 40909
rect 21489 40807 21523 40841
rect 21489 40739 21523 40773
rect 21489 40671 21523 40705
rect 21489 40603 21523 40637
rect 21489 40535 21523 40569
rect 21489 40467 21523 40501
rect 21489 40399 21523 40433
rect 21489 40331 21523 40365
rect 21489 40263 21523 40297
rect 21489 40195 21523 40229
rect 21489 40127 21523 40161
rect 21489 40059 21523 40093
rect 21489 39991 21523 40025
rect 21489 39923 21523 39957
rect 21947 41147 21981 41181
rect 21947 41079 21981 41113
rect 21947 41011 21981 41045
rect 21947 40943 21981 40977
rect 21947 40875 21981 40909
rect 21947 40807 21981 40841
rect 21947 40739 21981 40773
rect 21947 40671 21981 40705
rect 21947 40603 21981 40637
rect 21947 40535 21981 40569
rect 21947 40467 21981 40501
rect 21947 40399 21981 40433
rect 21947 40331 21981 40365
rect 21947 40263 21981 40297
rect 21947 40195 21981 40229
rect 21947 40127 21981 40161
rect 21947 40059 21981 40093
rect 21947 39991 21981 40025
rect 21947 39923 21981 39957
rect 22405 41147 22439 41181
rect 22405 41079 22439 41113
rect 22405 41011 22439 41045
rect 22405 40943 22439 40977
rect 22405 40875 22439 40909
rect 22405 40807 22439 40841
rect 22405 40739 22439 40773
rect 22405 40671 22439 40705
rect 22405 40603 22439 40637
rect 22405 40535 22439 40569
rect 22405 40467 22439 40501
rect 22405 40399 22439 40433
rect 22405 40331 22439 40365
rect 22405 40263 22439 40297
rect 22405 40195 22439 40229
rect 22405 40127 22439 40161
rect 22405 40059 22439 40093
rect 22405 39991 22439 40025
rect 22405 39923 22439 39957
rect 22863 41147 22897 41181
rect 22863 41079 22897 41113
rect 22863 41011 22897 41045
rect 22863 40943 22897 40977
rect 22863 40875 22897 40909
rect 22863 40807 22897 40841
rect 22863 40739 22897 40773
rect 22863 40671 22897 40705
rect 22863 40603 22897 40637
rect 22863 40535 22897 40569
rect 22863 40467 22897 40501
rect 22863 40399 22897 40433
rect 22863 40331 22897 40365
rect 22863 40263 22897 40297
rect 22863 40195 22897 40229
rect 22863 40127 22897 40161
rect 22863 40059 22897 40093
rect 22863 39991 22897 40025
rect 22863 39923 22897 39957
rect 23321 41147 23355 41181
rect 23321 41079 23355 41113
rect 23321 41011 23355 41045
rect 23321 40943 23355 40977
rect 23321 40875 23355 40909
rect 23321 40807 23355 40841
rect 23321 40739 23355 40773
rect 23321 40671 23355 40705
rect 23321 40603 23355 40637
rect 23321 40535 23355 40569
rect 23321 40467 23355 40501
rect 23321 40399 23355 40433
rect 23321 40331 23355 40365
rect 23321 40263 23355 40297
rect 23321 40195 23355 40229
rect 23321 40127 23355 40161
rect 23321 40059 23355 40093
rect 23321 39991 23355 40025
rect 23321 39923 23355 39957
rect 23779 41147 23813 41181
rect 23779 41079 23813 41113
rect 23779 41011 23813 41045
rect 23779 40943 23813 40977
rect 23779 40875 23813 40909
rect 23779 40807 23813 40841
rect 23779 40739 23813 40773
rect 23779 40671 23813 40705
rect 23779 40603 23813 40637
rect 23779 40535 23813 40569
rect 23779 40467 23813 40501
rect 23779 40399 23813 40433
rect 23779 40331 23813 40365
rect 23779 40263 23813 40297
rect 23779 40195 23813 40229
rect 23779 40127 23813 40161
rect 23779 40059 23813 40093
rect 23779 39991 23813 40025
rect 23779 39923 23813 39957
rect 24237 41147 24271 41181
rect 24237 41079 24271 41113
rect 24237 41011 24271 41045
rect 24237 40943 24271 40977
rect 24237 40875 24271 40909
rect 24237 40807 24271 40841
rect 24237 40739 24271 40773
rect 24237 40671 24271 40705
rect 24237 40603 24271 40637
rect 24237 40535 24271 40569
rect 24237 40467 24271 40501
rect 24237 40399 24271 40433
rect 24237 40331 24271 40365
rect 24237 40263 24271 40297
rect 24237 40195 24271 40229
rect 24237 40127 24271 40161
rect 24237 40059 24271 40093
rect 24237 39991 24271 40025
rect 24237 39923 24271 39957
rect 24695 41147 24729 41181
rect 24695 41079 24729 41113
rect 24695 41011 24729 41045
rect 24695 40943 24729 40977
rect 24695 40875 24729 40909
rect 24695 40807 24729 40841
rect 24695 40739 24729 40773
rect 24695 40671 24729 40705
rect 24695 40603 24729 40637
rect 24695 40535 24729 40569
rect 24695 40467 24729 40501
rect 24695 40399 24729 40433
rect 24695 40331 24729 40365
rect 24695 40263 24729 40297
rect 24695 40195 24729 40229
rect 24695 40127 24729 40161
rect 24695 40059 24729 40093
rect 24695 39991 24729 40025
rect 24695 39923 24729 39957
rect 25153 41147 25187 41181
rect 25153 41079 25187 41113
rect 25153 41011 25187 41045
rect 25153 40943 25187 40977
rect 25153 40875 25187 40909
rect 25153 40807 25187 40841
rect 25153 40739 25187 40773
rect 25153 40671 25187 40705
rect 25153 40603 25187 40637
rect 25153 40535 25187 40569
rect 25153 40467 25187 40501
rect 25153 40399 25187 40433
rect 25153 40331 25187 40365
rect 25153 40263 25187 40297
rect 25153 40195 25187 40229
rect 25153 40127 25187 40161
rect 25153 40059 25187 40093
rect 25153 39991 25187 40025
rect 25153 39923 25187 39957
rect 25611 41147 25645 41181
rect 25611 41079 25645 41113
rect 25611 41011 25645 41045
rect 25611 40943 25645 40977
rect 25611 40875 25645 40909
rect 25611 40807 25645 40841
rect 25611 40739 25645 40773
rect 25611 40671 25645 40705
rect 25611 40603 25645 40637
rect 25611 40535 25645 40569
rect 25611 40467 25645 40501
rect 25611 40399 25645 40433
rect 25611 40331 25645 40365
rect 25611 40263 25645 40297
rect 25611 40195 25645 40229
rect 25611 40127 25645 40161
rect 25611 40059 25645 40093
rect 25611 39991 25645 40025
rect 25611 39923 25645 39957
rect 26069 41147 26103 41181
rect 26069 41079 26103 41113
rect 26069 41011 26103 41045
rect 26069 40943 26103 40977
rect 26069 40875 26103 40909
rect 26069 40807 26103 40841
rect 26069 40739 26103 40773
rect 26069 40671 26103 40705
rect 26069 40603 26103 40637
rect 26069 40535 26103 40569
rect 26069 40467 26103 40501
rect 26069 40399 26103 40433
rect 26069 40331 26103 40365
rect 26069 40263 26103 40297
rect 26069 40195 26103 40229
rect 26069 40127 26103 40161
rect 26069 40059 26103 40093
rect 26069 39991 26103 40025
rect 26069 39923 26103 39957
rect 26527 41147 26561 41181
rect 26527 41079 26561 41113
rect 26527 41011 26561 41045
rect 26527 40943 26561 40977
rect 26527 40875 26561 40909
rect 26527 40807 26561 40841
rect 26527 40739 26561 40773
rect 26527 40671 26561 40705
rect 26527 40603 26561 40637
rect 26527 40535 26561 40569
rect 26527 40467 26561 40501
rect 26527 40399 26561 40433
rect 26527 40331 26561 40365
rect 26527 40263 26561 40297
rect 26527 40195 26561 40229
rect 26527 40127 26561 40161
rect 26527 40059 26561 40093
rect 26527 39991 26561 40025
rect 26527 39923 26561 39957
rect 26985 41147 27019 41181
rect 26985 41079 27019 41113
rect 26985 41011 27019 41045
rect 26985 40943 27019 40977
rect 26985 40875 27019 40909
rect 26985 40807 27019 40841
rect 26985 40739 27019 40773
rect 26985 40671 27019 40705
rect 26985 40603 27019 40637
rect 26985 40535 27019 40569
rect 26985 40467 27019 40501
rect 26985 40399 27019 40433
rect 26985 40331 27019 40365
rect 26985 40263 27019 40297
rect 26985 40195 27019 40229
rect 26985 40127 27019 40161
rect 26985 40059 27019 40093
rect 26985 39991 27019 40025
rect 26985 39923 27019 39957
rect 27443 41147 27477 41181
rect 27443 41079 27477 41113
rect 27443 41011 27477 41045
rect 27443 40943 27477 40977
rect 27443 40875 27477 40909
rect 27443 40807 27477 40841
rect 27443 40739 27477 40773
rect 27443 40671 27477 40705
rect 27443 40603 27477 40637
rect 27443 40535 27477 40569
rect 27443 40467 27477 40501
rect 27443 40399 27477 40433
rect 27443 40331 27477 40365
rect 27443 40263 27477 40297
rect 27443 40195 27477 40229
rect 27443 40127 27477 40161
rect 27443 40059 27477 40093
rect 27443 39991 27477 40025
rect 27443 39923 27477 39957
rect 27901 41147 27935 41181
rect 27901 41079 27935 41113
rect 27901 41011 27935 41045
rect 27901 40943 27935 40977
rect 27901 40875 27935 40909
rect 27901 40807 27935 40841
rect 27901 40739 27935 40773
rect 27901 40671 27935 40705
rect 27901 40603 27935 40637
rect 27901 40535 27935 40569
rect 27901 40467 27935 40501
rect 27901 40399 27935 40433
rect 27901 40331 27935 40365
rect 27901 40263 27935 40297
rect 27901 40195 27935 40229
rect 27901 40127 27935 40161
rect 27901 40059 27935 40093
rect 27901 39991 27935 40025
rect 27901 39923 27935 39957
rect 28359 41147 28393 41181
rect 28359 41079 28393 41113
rect 28359 41011 28393 41045
rect 28359 40943 28393 40977
rect 28359 40875 28393 40909
rect 28359 40807 28393 40841
rect 28359 40739 28393 40773
rect 28359 40671 28393 40705
rect 28359 40603 28393 40637
rect 28359 40535 28393 40569
rect 28359 40467 28393 40501
rect 28359 40399 28393 40433
rect 28359 40331 28393 40365
rect 28359 40263 28393 40297
rect 28359 40195 28393 40229
rect 28359 40127 28393 40161
rect 28359 40059 28393 40093
rect 28359 39991 28393 40025
rect 28359 39923 28393 39957
rect 28817 41147 28851 41181
rect 28817 41079 28851 41113
rect 28817 41011 28851 41045
rect 28817 40943 28851 40977
rect 28817 40875 28851 40909
rect 28817 40807 28851 40841
rect 28817 40739 28851 40773
rect 28817 40671 28851 40705
rect 28817 40603 28851 40637
rect 28817 40535 28851 40569
rect 28817 40467 28851 40501
rect 28817 40399 28851 40433
rect 28817 40331 28851 40365
rect 28817 40263 28851 40297
rect 28817 40195 28851 40229
rect 28817 40127 28851 40161
rect 28817 40059 28851 40093
rect 28817 39991 28851 40025
rect 28817 39923 28851 39957
rect 29275 41147 29309 41181
rect 29275 41079 29309 41113
rect 29275 41011 29309 41045
rect 29275 40943 29309 40977
rect 29275 40875 29309 40909
rect 29275 40807 29309 40841
rect 29275 40739 29309 40773
rect 29275 40671 29309 40705
rect 29275 40603 29309 40637
rect 29275 40535 29309 40569
rect 29275 40467 29309 40501
rect 29275 40399 29309 40433
rect 29275 40331 29309 40365
rect 29275 40263 29309 40297
rect 29275 40195 29309 40229
rect 29275 40127 29309 40161
rect 29275 40059 29309 40093
rect 29275 39991 29309 40025
rect 29275 39923 29309 39957
rect 29733 41147 29767 41181
rect 29733 41079 29767 41113
rect 29733 41011 29767 41045
rect 29733 40943 29767 40977
rect 29733 40875 29767 40909
rect 29733 40807 29767 40841
rect 29733 40739 29767 40773
rect 29733 40671 29767 40705
rect 29733 40603 29767 40637
rect 29733 40535 29767 40569
rect 29733 40467 29767 40501
rect 29733 40399 29767 40433
rect 29733 40331 29767 40365
rect 29733 40263 29767 40297
rect 29733 40195 29767 40229
rect 29733 40127 29767 40161
rect 29733 40059 29767 40093
rect 29733 39991 29767 40025
rect 29733 39923 29767 39957
rect 30191 41147 30225 41181
rect 30191 41079 30225 41113
rect 30191 41011 30225 41045
rect 30191 40943 30225 40977
rect 30191 40875 30225 40909
rect 30191 40807 30225 40841
rect 30191 40739 30225 40773
rect 30191 40671 30225 40705
rect 30191 40603 30225 40637
rect 30191 40535 30225 40569
rect 30191 40467 30225 40501
rect 30191 40399 30225 40433
rect 30191 40331 30225 40365
rect 30191 40263 30225 40297
rect 30191 40195 30225 40229
rect 30191 40127 30225 40161
rect 30191 40059 30225 40093
rect 30191 39991 30225 40025
rect 30191 39923 30225 39957
rect 30649 41147 30683 41181
rect 30649 41079 30683 41113
rect 30649 41011 30683 41045
rect 30649 40943 30683 40977
rect 30649 40875 30683 40909
rect 30649 40807 30683 40841
rect 30649 40739 30683 40773
rect 30649 40671 30683 40705
rect 30649 40603 30683 40637
rect 30649 40535 30683 40569
rect 30649 40467 30683 40501
rect 30649 40399 30683 40433
rect 30649 40331 30683 40365
rect 30649 40263 30683 40297
rect 30649 40195 30683 40229
rect 30649 40127 30683 40161
rect 30649 40059 30683 40093
rect 30649 39991 30683 40025
rect 30649 39923 30683 39957
rect 31107 41147 31141 41181
rect 31107 41079 31141 41113
rect 31107 41011 31141 41045
rect 31107 40943 31141 40977
rect 31107 40875 31141 40909
rect 31107 40807 31141 40841
rect 31107 40739 31141 40773
rect 31107 40671 31141 40705
rect 31107 40603 31141 40637
rect 31107 40535 31141 40569
rect 31107 40467 31141 40501
rect 31107 40399 31141 40433
rect 31107 40331 31141 40365
rect 31107 40263 31141 40297
rect 31107 40195 31141 40229
rect 31107 40127 31141 40161
rect 31107 40059 31141 40093
rect 31107 39991 31141 40025
rect 31107 39923 31141 39957
rect 31565 41147 31599 41181
rect 31565 41079 31599 41113
rect 31565 41011 31599 41045
rect 31565 40943 31599 40977
rect 31565 40875 31599 40909
rect 31565 40807 31599 40841
rect 31565 40739 31599 40773
rect 31565 40671 31599 40705
rect 31565 40603 31599 40637
rect 31565 40535 31599 40569
rect 31565 40467 31599 40501
rect 31565 40399 31599 40433
rect 31565 40331 31599 40365
rect 31565 40263 31599 40297
rect 31565 40195 31599 40229
rect 31565 40127 31599 40161
rect 31565 40059 31599 40093
rect 31565 39991 31599 40025
rect 31565 39923 31599 39957
rect 32023 41147 32057 41181
rect 32023 41079 32057 41113
rect 32023 41011 32057 41045
rect 32023 40943 32057 40977
rect 32023 40875 32057 40909
rect 32023 40807 32057 40841
rect 32023 40739 32057 40773
rect 32023 40671 32057 40705
rect 32023 40603 32057 40637
rect 32023 40535 32057 40569
rect 32023 40467 32057 40501
rect 32023 40399 32057 40433
rect 32023 40331 32057 40365
rect 32023 40263 32057 40297
rect 32023 40195 32057 40229
rect 32023 40127 32057 40161
rect 32023 40059 32057 40093
rect 32023 39991 32057 40025
rect 32023 39923 32057 39957
rect 32481 41147 32515 41181
rect 32481 41079 32515 41113
rect 32481 41011 32515 41045
rect 32481 40943 32515 40977
rect 32481 40875 32515 40909
rect 32481 40807 32515 40841
rect 32481 40739 32515 40773
rect 32481 40671 32515 40705
rect 32481 40603 32515 40637
rect 32481 40535 32515 40569
rect 32481 40467 32515 40501
rect 32481 40399 32515 40433
rect 32481 40331 32515 40365
rect 32481 40263 32515 40297
rect 32481 40195 32515 40229
rect 32481 40127 32515 40161
rect 32481 40059 32515 40093
rect 32481 39991 32515 40025
rect 32481 39923 32515 39957
rect 32939 41147 32973 41181
rect 32939 41079 32973 41113
rect 32939 41011 32973 41045
rect 32939 40943 32973 40977
rect 32939 40875 32973 40909
rect 32939 40807 32973 40841
rect 32939 40739 32973 40773
rect 32939 40671 32973 40705
rect 32939 40603 32973 40637
rect 32939 40535 32973 40569
rect 32939 40467 32973 40501
rect 32939 40399 32973 40433
rect 32939 40331 32973 40365
rect 32939 40263 32973 40297
rect 32939 40195 32973 40229
rect 32939 40127 32973 40161
rect 32939 40059 32973 40093
rect 32939 39991 32973 40025
rect 32939 39923 32973 39957
rect 33397 41147 33431 41181
rect 33397 41079 33431 41113
rect 33397 41011 33431 41045
rect 33397 40943 33431 40977
rect 33397 40875 33431 40909
rect 33397 40807 33431 40841
rect 33397 40739 33431 40773
rect 33397 40671 33431 40705
rect 33397 40603 33431 40637
rect 33397 40535 33431 40569
rect 33397 40467 33431 40501
rect 33397 40399 33431 40433
rect 33397 40331 33431 40365
rect 33397 40263 33431 40297
rect 33397 40195 33431 40229
rect 33397 40127 33431 40161
rect 33397 40059 33431 40093
rect 33397 39991 33431 40025
rect 33397 39923 33431 39957
rect 33855 41147 33889 41181
rect 33855 41079 33889 41113
rect 33855 41011 33889 41045
rect 33855 40943 33889 40977
rect 33855 40875 33889 40909
rect 33855 40807 33889 40841
rect 33855 40739 33889 40773
rect 33855 40671 33889 40705
rect 33855 40603 33889 40637
rect 33855 40535 33889 40569
rect 33855 40467 33889 40501
rect 33855 40399 33889 40433
rect 33855 40331 33889 40365
rect 33855 40263 33889 40297
rect 33855 40195 33889 40229
rect 33855 40127 33889 40161
rect 33855 40059 33889 40093
rect 33855 39991 33889 40025
rect 33855 39923 33889 39957
rect 34313 41147 34347 41181
rect 34313 41079 34347 41113
rect 34313 41011 34347 41045
rect 34313 40943 34347 40977
rect 34313 40875 34347 40909
rect 34313 40807 34347 40841
rect 34313 40739 34347 40773
rect 34313 40671 34347 40705
rect 34313 40603 34347 40637
rect 34313 40535 34347 40569
rect 34313 40467 34347 40501
rect 34313 40399 34347 40433
rect 34313 40331 34347 40365
rect 34313 40263 34347 40297
rect 34313 40195 34347 40229
rect 34313 40127 34347 40161
rect 34313 40059 34347 40093
rect 34313 39991 34347 40025
rect 34313 39923 34347 39957
rect 34771 41147 34805 41181
rect 34771 41079 34805 41113
rect 34771 41011 34805 41045
rect 34771 40943 34805 40977
rect 34771 40875 34805 40909
rect 34771 40807 34805 40841
rect 34771 40739 34805 40773
rect 34771 40671 34805 40705
rect 34771 40603 34805 40637
rect 34771 40535 34805 40569
rect 34771 40467 34805 40501
rect 34771 40399 34805 40433
rect 34771 40331 34805 40365
rect 34771 40263 34805 40297
rect 34771 40195 34805 40229
rect 34771 40127 34805 40161
rect 34771 40059 34805 40093
rect 34771 39991 34805 40025
rect 34771 39923 34805 39957
rect 35229 41147 35263 41181
rect 35229 41079 35263 41113
rect 35229 41011 35263 41045
rect 35229 40943 35263 40977
rect 35229 40875 35263 40909
rect 35229 40807 35263 40841
rect 35229 40739 35263 40773
rect 35229 40671 35263 40705
rect 35229 40603 35263 40637
rect 35229 40535 35263 40569
rect 35229 40467 35263 40501
rect 35229 40399 35263 40433
rect 35229 40331 35263 40365
rect 35229 40263 35263 40297
rect 35229 40195 35263 40229
rect 35229 40127 35263 40161
rect 35229 40059 35263 40093
rect 35229 39991 35263 40025
rect 35229 39923 35263 39957
rect 35687 41147 35721 41181
rect 35687 41079 35721 41113
rect 35687 41011 35721 41045
rect 35687 40943 35721 40977
rect 35687 40875 35721 40909
rect 35687 40807 35721 40841
rect 35687 40739 35721 40773
rect 35687 40671 35721 40705
rect 35687 40603 35721 40637
rect 35687 40535 35721 40569
rect 35687 40467 35721 40501
rect 35687 40399 35721 40433
rect 35687 40331 35721 40365
rect 35687 40263 35721 40297
rect 35687 40195 35721 40229
rect 35687 40127 35721 40161
rect 35687 40059 35721 40093
rect 35687 39991 35721 40025
rect 35687 39923 35721 39957
rect 36145 41147 36179 41181
rect 36145 41079 36179 41113
rect 36145 41011 36179 41045
rect 36145 40943 36179 40977
rect 36145 40875 36179 40909
rect 36145 40807 36179 40841
rect 36145 40739 36179 40773
rect 36145 40671 36179 40705
rect 36145 40603 36179 40637
rect 36145 40535 36179 40569
rect 36145 40467 36179 40501
rect 36145 40399 36179 40433
rect 36145 40331 36179 40365
rect 36145 40263 36179 40297
rect 36145 40195 36179 40229
rect 36145 40127 36179 40161
rect 36145 40059 36179 40093
rect 36145 39991 36179 40025
rect 36145 39923 36179 39957
rect 36603 41147 36637 41181
rect 36603 41079 36637 41113
rect 36603 41011 36637 41045
rect 36603 40943 36637 40977
rect 36603 40875 36637 40909
rect 36603 40807 36637 40841
rect 36603 40739 36637 40773
rect 36603 40671 36637 40705
rect 36603 40603 36637 40637
rect 36603 40535 36637 40569
rect 36603 40467 36637 40501
rect 36603 40399 36637 40433
rect 36603 40331 36637 40365
rect 36603 40263 36637 40297
rect 36603 40195 36637 40229
rect 36603 40127 36637 40161
rect 36603 40059 36637 40093
rect 36603 39991 36637 40025
rect 36603 39923 36637 39957
rect 37061 41147 37095 41181
rect 37061 41079 37095 41113
rect 37061 41011 37095 41045
rect 37061 40943 37095 40977
rect 37061 40875 37095 40909
rect 37061 40807 37095 40841
rect 37061 40739 37095 40773
rect 37061 40671 37095 40705
rect 37061 40603 37095 40637
rect 37061 40535 37095 40569
rect 37061 40467 37095 40501
rect 37061 40399 37095 40433
rect 37061 40331 37095 40365
rect 37061 40263 37095 40297
rect 37061 40195 37095 40229
rect 37061 40127 37095 40161
rect 37061 40059 37095 40093
rect 37061 39991 37095 40025
rect 37061 39923 37095 39957
rect 37519 41147 37553 41181
rect 37519 41079 37553 41113
rect 37519 41011 37553 41045
rect 37519 40943 37553 40977
rect 37519 40875 37553 40909
rect 37519 40807 37553 40841
rect 37519 40739 37553 40773
rect 37519 40671 37553 40705
rect 37519 40603 37553 40637
rect 37519 40535 37553 40569
rect 37519 40467 37553 40501
rect 37519 40399 37553 40433
rect 37519 40331 37553 40365
rect 37519 40263 37553 40297
rect 37519 40195 37553 40229
rect 37519 40127 37553 40161
rect 37519 40059 37553 40093
rect 37519 39991 37553 40025
rect 37519 39923 37553 39957
rect 37977 41147 38011 41181
rect 37977 41079 38011 41113
rect 37977 41011 38011 41045
rect 37977 40943 38011 40977
rect 37977 40875 38011 40909
rect 37977 40807 38011 40841
rect 37977 40739 38011 40773
rect 37977 40671 38011 40705
rect 37977 40603 38011 40637
rect 37977 40535 38011 40569
rect 37977 40467 38011 40501
rect 37977 40399 38011 40433
rect 37977 40331 38011 40365
rect 37977 40263 38011 40297
rect 37977 40195 38011 40229
rect 37977 40127 38011 40161
rect 37977 40059 38011 40093
rect 37977 39991 38011 40025
rect 37977 39923 38011 39957
rect 38435 41147 38469 41181
rect 38435 41079 38469 41113
rect 38435 41011 38469 41045
rect 38435 40943 38469 40977
rect 38435 40875 38469 40909
rect 38435 40807 38469 40841
rect 38435 40739 38469 40773
rect 38435 40671 38469 40705
rect 38435 40603 38469 40637
rect 38435 40535 38469 40569
rect 38435 40467 38469 40501
rect 38435 40399 38469 40433
rect 38435 40331 38469 40365
rect 38435 40263 38469 40297
rect 38435 40195 38469 40229
rect 38435 40127 38469 40161
rect 38435 40059 38469 40093
rect 38435 39991 38469 40025
rect 38435 39923 38469 39957
rect 38893 41147 38927 41181
rect 38893 41079 38927 41113
rect 38893 41011 38927 41045
rect 38893 40943 38927 40977
rect 38893 40875 38927 40909
rect 38893 40807 38927 40841
rect 38893 40739 38927 40773
rect 38893 40671 38927 40705
rect 38893 40603 38927 40637
rect 38893 40535 38927 40569
rect 38893 40467 38927 40501
rect 38893 40399 38927 40433
rect 38893 40331 38927 40365
rect 38893 40263 38927 40297
rect 38893 40195 38927 40229
rect 38893 40127 38927 40161
rect 38893 40059 38927 40093
rect 38893 39991 38927 40025
rect 38893 39923 38927 39957
rect 39351 41147 39385 41181
rect 39351 41079 39385 41113
rect 39351 41011 39385 41045
rect 39351 40943 39385 40977
rect 39351 40875 39385 40909
rect 39351 40807 39385 40841
rect 39351 40739 39385 40773
rect 39351 40671 39385 40705
rect 39351 40603 39385 40637
rect 39351 40535 39385 40569
rect 39351 40467 39385 40501
rect 39351 40399 39385 40433
rect 39351 40331 39385 40365
rect 39351 40263 39385 40297
rect 39351 40195 39385 40229
rect 39351 40127 39385 40161
rect 39351 40059 39385 40093
rect 39351 39991 39385 40025
rect 39351 39923 39385 39957
rect 39809 41147 39843 41181
rect 39809 41079 39843 41113
rect 39809 41011 39843 41045
rect 39809 40943 39843 40977
rect 39809 40875 39843 40909
rect 39809 40807 39843 40841
rect 39809 40739 39843 40773
rect 39809 40671 39843 40705
rect 39809 40603 39843 40637
rect 39809 40535 39843 40569
rect 39809 40467 39843 40501
rect 39809 40399 39843 40433
rect 39809 40331 39843 40365
rect 39809 40263 39843 40297
rect 39809 40195 39843 40229
rect 39809 40127 39843 40161
rect 39809 40059 39843 40093
rect 39809 39991 39843 40025
rect 39809 39923 39843 39957
rect 40267 41147 40301 41181
rect 40267 41079 40301 41113
rect 40267 41011 40301 41045
rect 40267 40943 40301 40977
rect 40267 40875 40301 40909
rect 40267 40807 40301 40841
rect 40267 40739 40301 40773
rect 40267 40671 40301 40705
rect 40267 40603 40301 40637
rect 40267 40535 40301 40569
rect 40267 40467 40301 40501
rect 40267 40399 40301 40433
rect 40267 40331 40301 40365
rect 40267 40263 40301 40297
rect 40267 40195 40301 40229
rect 40267 40127 40301 40161
rect 40267 40059 40301 40093
rect 40267 39991 40301 40025
rect 40267 39923 40301 39957
rect 40725 41147 40759 41181
rect 40725 41079 40759 41113
rect 40725 41011 40759 41045
rect 40725 40943 40759 40977
rect 40725 40875 40759 40909
rect 40725 40807 40759 40841
rect 40725 40739 40759 40773
rect 40725 40671 40759 40705
rect 40725 40603 40759 40637
rect 40725 40535 40759 40569
rect 40725 40467 40759 40501
rect 40725 40399 40759 40433
rect 40725 40331 40759 40365
rect 40725 40263 40759 40297
rect 40725 40195 40759 40229
rect 40725 40127 40759 40161
rect 40725 40059 40759 40093
rect 40725 39991 40759 40025
rect 40725 39923 40759 39957
rect 41183 41147 41217 41181
rect 41183 41079 41217 41113
rect 41183 41011 41217 41045
rect 41183 40943 41217 40977
rect 41183 40875 41217 40909
rect 41183 40807 41217 40841
rect 41183 40739 41217 40773
rect 41183 40671 41217 40705
rect 41183 40603 41217 40637
rect 41183 40535 41217 40569
rect 41183 40467 41217 40501
rect 41183 40399 41217 40433
rect 41183 40331 41217 40365
rect 41183 40263 41217 40297
rect 41183 40195 41217 40229
rect 41183 40127 41217 40161
rect 41183 40059 41217 40093
rect 41183 39991 41217 40025
rect 41183 39923 41217 39957
rect 41641 41147 41675 41181
rect 41641 41079 41675 41113
rect 41641 41011 41675 41045
rect 41641 40943 41675 40977
rect 41641 40875 41675 40909
rect 41641 40807 41675 40841
rect 41641 40739 41675 40773
rect 41641 40671 41675 40705
rect 41641 40603 41675 40637
rect 41641 40535 41675 40569
rect 41641 40467 41675 40501
rect 41641 40399 41675 40433
rect 41641 40331 41675 40365
rect 41641 40263 41675 40297
rect 41641 40195 41675 40229
rect 41641 40127 41675 40161
rect 41641 40059 41675 40093
rect 41641 39991 41675 40025
rect 41641 39923 41675 39957
rect 42099 41147 42133 41181
rect 42099 41079 42133 41113
rect 42099 41011 42133 41045
rect 42099 40943 42133 40977
rect 42099 40875 42133 40909
rect 42099 40807 42133 40841
rect 42099 40739 42133 40773
rect 42099 40671 42133 40705
rect 42099 40603 42133 40637
rect 42099 40535 42133 40569
rect 42099 40467 42133 40501
rect 42099 40399 42133 40433
rect 42099 40331 42133 40365
rect 42099 40263 42133 40297
rect 42099 40195 42133 40229
rect 42099 40127 42133 40161
rect 42099 40059 42133 40093
rect 42099 39991 42133 40025
rect 42099 39923 42133 39957
rect 42557 41147 42591 41181
rect 42557 41079 42591 41113
rect 42557 41011 42591 41045
rect 42557 40943 42591 40977
rect 42557 40875 42591 40909
rect 42557 40807 42591 40841
rect 42557 40739 42591 40773
rect 42557 40671 42591 40705
rect 42557 40603 42591 40637
rect 42557 40535 42591 40569
rect 42557 40467 42591 40501
rect 42557 40399 42591 40433
rect 42557 40331 42591 40365
rect 42557 40263 42591 40297
rect 42557 40195 42591 40229
rect 42557 40127 42591 40161
rect 42557 40059 42591 40093
rect 42557 39991 42591 40025
rect 42557 39923 42591 39957
rect 30408 36986 30442 37020
rect 30498 36986 30532 37020
rect 30588 36986 30622 37020
rect 30678 36986 30712 37020
rect 30768 36986 30802 37020
rect 30858 36986 30892 37020
rect 30948 36986 30982 37020
rect 30408 36896 30442 36930
rect 30498 36896 30532 36930
rect 30588 36896 30622 36930
rect 30678 36896 30712 36930
rect 30768 36896 30802 36930
rect 30858 36896 30892 36930
rect 30948 36896 30982 36930
rect 30408 36806 30442 36840
rect 30498 36806 30532 36840
rect 30588 36806 30622 36840
rect 30678 36806 30712 36840
rect 30768 36806 30802 36840
rect 30858 36806 30892 36840
rect 30948 36806 30982 36840
rect 30408 36716 30442 36750
rect 30498 36716 30532 36750
rect 30588 36716 30622 36750
rect 30678 36716 30712 36750
rect 30768 36716 30802 36750
rect 30858 36716 30892 36750
rect 30948 36716 30982 36750
rect 30408 36626 30442 36660
rect 30498 36626 30532 36660
rect 30588 36626 30622 36660
rect 30678 36626 30712 36660
rect 30768 36626 30802 36660
rect 30858 36626 30892 36660
rect 30948 36626 30982 36660
rect 30408 36536 30442 36570
rect 30498 36536 30532 36570
rect 30588 36536 30622 36570
rect 30678 36536 30712 36570
rect 30768 36536 30802 36570
rect 30858 36536 30892 36570
rect 30948 36536 30982 36570
rect 30408 36446 30442 36480
rect 30498 36446 30532 36480
rect 30588 36446 30622 36480
rect 30678 36446 30712 36480
rect 30768 36446 30802 36480
rect 30858 36446 30892 36480
rect 30948 36446 30982 36480
rect 31748 36986 31782 37020
rect 31838 36986 31872 37020
rect 31928 36986 31962 37020
rect 32018 36986 32052 37020
rect 32108 36986 32142 37020
rect 32198 36986 32232 37020
rect 32288 36986 32322 37020
rect 31748 36896 31782 36930
rect 31838 36896 31872 36930
rect 31928 36896 31962 36930
rect 32018 36896 32052 36930
rect 32108 36896 32142 36930
rect 32198 36896 32232 36930
rect 32288 36896 32322 36930
rect 31748 36806 31782 36840
rect 31838 36806 31872 36840
rect 31928 36806 31962 36840
rect 32018 36806 32052 36840
rect 32108 36806 32142 36840
rect 32198 36806 32232 36840
rect 32288 36806 32322 36840
rect 31748 36716 31782 36750
rect 31838 36716 31872 36750
rect 31928 36716 31962 36750
rect 32018 36716 32052 36750
rect 32108 36716 32142 36750
rect 32198 36716 32232 36750
rect 32288 36716 32322 36750
rect 31748 36626 31782 36660
rect 31838 36626 31872 36660
rect 31928 36626 31962 36660
rect 32018 36626 32052 36660
rect 32108 36626 32142 36660
rect 32198 36626 32232 36660
rect 32288 36626 32322 36660
rect 31748 36536 31782 36570
rect 31838 36536 31872 36570
rect 31928 36536 31962 36570
rect 32018 36536 32052 36570
rect 32108 36536 32142 36570
rect 32198 36536 32232 36570
rect 32288 36536 32322 36570
rect 31748 36446 31782 36480
rect 31838 36446 31872 36480
rect 31928 36446 31962 36480
rect 32018 36446 32052 36480
rect 32108 36446 32142 36480
rect 32198 36446 32232 36480
rect 32288 36446 32322 36480
rect 33088 36986 33122 37020
rect 33178 36986 33212 37020
rect 33268 36986 33302 37020
rect 33358 36986 33392 37020
rect 33448 36986 33482 37020
rect 33538 36986 33572 37020
rect 33628 36986 33662 37020
rect 33088 36896 33122 36930
rect 33178 36896 33212 36930
rect 33268 36896 33302 36930
rect 33358 36896 33392 36930
rect 33448 36896 33482 36930
rect 33538 36896 33572 36930
rect 33628 36896 33662 36930
rect 33088 36806 33122 36840
rect 33178 36806 33212 36840
rect 33268 36806 33302 36840
rect 33358 36806 33392 36840
rect 33448 36806 33482 36840
rect 33538 36806 33572 36840
rect 33628 36806 33662 36840
rect 33088 36716 33122 36750
rect 33178 36716 33212 36750
rect 33268 36716 33302 36750
rect 33358 36716 33392 36750
rect 33448 36716 33482 36750
rect 33538 36716 33572 36750
rect 33628 36716 33662 36750
rect 33088 36626 33122 36660
rect 33178 36626 33212 36660
rect 33268 36626 33302 36660
rect 33358 36626 33392 36660
rect 33448 36626 33482 36660
rect 33538 36626 33572 36660
rect 33628 36626 33662 36660
rect 33088 36536 33122 36570
rect 33178 36536 33212 36570
rect 33268 36536 33302 36570
rect 33358 36536 33392 36570
rect 33448 36536 33482 36570
rect 33538 36536 33572 36570
rect 33628 36536 33662 36570
rect 33088 36446 33122 36480
rect 33178 36446 33212 36480
rect 33268 36446 33302 36480
rect 33358 36446 33392 36480
rect 33448 36446 33482 36480
rect 33538 36446 33572 36480
rect 33628 36446 33662 36480
rect 34428 36986 34462 37020
rect 34518 36986 34552 37020
rect 34608 36986 34642 37020
rect 34698 36986 34732 37020
rect 34788 36986 34822 37020
rect 34878 36986 34912 37020
rect 34968 36986 35002 37020
rect 34428 36896 34462 36930
rect 34518 36896 34552 36930
rect 34608 36896 34642 36930
rect 34698 36896 34732 36930
rect 34788 36896 34822 36930
rect 34878 36896 34912 36930
rect 34968 36896 35002 36930
rect 34428 36806 34462 36840
rect 34518 36806 34552 36840
rect 34608 36806 34642 36840
rect 34698 36806 34732 36840
rect 34788 36806 34822 36840
rect 34878 36806 34912 36840
rect 34968 36806 35002 36840
rect 34428 36716 34462 36750
rect 34518 36716 34552 36750
rect 34608 36716 34642 36750
rect 34698 36716 34732 36750
rect 34788 36716 34822 36750
rect 34878 36716 34912 36750
rect 34968 36716 35002 36750
rect 34428 36626 34462 36660
rect 34518 36626 34552 36660
rect 34608 36626 34642 36660
rect 34698 36626 34732 36660
rect 34788 36626 34822 36660
rect 34878 36626 34912 36660
rect 34968 36626 35002 36660
rect 34428 36536 34462 36570
rect 34518 36536 34552 36570
rect 34608 36536 34642 36570
rect 34698 36536 34732 36570
rect 34788 36536 34822 36570
rect 34878 36536 34912 36570
rect 34968 36536 35002 36570
rect 34428 36446 34462 36480
rect 34518 36446 34552 36480
rect 34608 36446 34642 36480
rect 34698 36446 34732 36480
rect 34788 36446 34822 36480
rect 34878 36446 34912 36480
rect 34968 36446 35002 36480
rect 35768 36986 35802 37020
rect 35858 36986 35892 37020
rect 35948 36986 35982 37020
rect 36038 36986 36072 37020
rect 36128 36986 36162 37020
rect 36218 36986 36252 37020
rect 36308 36986 36342 37020
rect 35768 36896 35802 36930
rect 35858 36896 35892 36930
rect 35948 36896 35982 36930
rect 36038 36896 36072 36930
rect 36128 36896 36162 36930
rect 36218 36896 36252 36930
rect 36308 36896 36342 36930
rect 35768 36806 35802 36840
rect 35858 36806 35892 36840
rect 35948 36806 35982 36840
rect 36038 36806 36072 36840
rect 36128 36806 36162 36840
rect 36218 36806 36252 36840
rect 36308 36806 36342 36840
rect 35768 36716 35802 36750
rect 35858 36716 35892 36750
rect 35948 36716 35982 36750
rect 36038 36716 36072 36750
rect 36128 36716 36162 36750
rect 36218 36716 36252 36750
rect 36308 36716 36342 36750
rect 35768 36626 35802 36660
rect 35858 36626 35892 36660
rect 35948 36626 35982 36660
rect 36038 36626 36072 36660
rect 36128 36626 36162 36660
rect 36218 36626 36252 36660
rect 36308 36626 36342 36660
rect 35768 36536 35802 36570
rect 35858 36536 35892 36570
rect 35948 36536 35982 36570
rect 36038 36536 36072 36570
rect 36128 36536 36162 36570
rect 36218 36536 36252 36570
rect 36308 36536 36342 36570
rect 35768 36446 35802 36480
rect 35858 36446 35892 36480
rect 35948 36446 35982 36480
rect 36038 36446 36072 36480
rect 36128 36446 36162 36480
rect 36218 36446 36252 36480
rect 36308 36446 36342 36480
rect 37108 36986 37142 37020
rect 37198 36986 37232 37020
rect 37288 36986 37322 37020
rect 37378 36986 37412 37020
rect 37468 36986 37502 37020
rect 37558 36986 37592 37020
rect 37648 36986 37682 37020
rect 37108 36896 37142 36930
rect 37198 36896 37232 36930
rect 37288 36896 37322 36930
rect 37378 36896 37412 36930
rect 37468 36896 37502 36930
rect 37558 36896 37592 36930
rect 37648 36896 37682 36930
rect 37108 36806 37142 36840
rect 37198 36806 37232 36840
rect 37288 36806 37322 36840
rect 37378 36806 37412 36840
rect 37468 36806 37502 36840
rect 37558 36806 37592 36840
rect 37648 36806 37682 36840
rect 37108 36716 37142 36750
rect 37198 36716 37232 36750
rect 37288 36716 37322 36750
rect 37378 36716 37412 36750
rect 37468 36716 37502 36750
rect 37558 36716 37592 36750
rect 37648 36716 37682 36750
rect 37108 36626 37142 36660
rect 37198 36626 37232 36660
rect 37288 36626 37322 36660
rect 37378 36626 37412 36660
rect 37468 36626 37502 36660
rect 37558 36626 37592 36660
rect 37648 36626 37682 36660
rect 37108 36536 37142 36570
rect 37198 36536 37232 36570
rect 37288 36536 37322 36570
rect 37378 36536 37412 36570
rect 37468 36536 37502 36570
rect 37558 36536 37592 36570
rect 37648 36536 37682 36570
rect 37108 36446 37142 36480
rect 37198 36446 37232 36480
rect 37288 36446 37322 36480
rect 37378 36446 37412 36480
rect 37468 36446 37502 36480
rect 37558 36446 37592 36480
rect 37648 36446 37682 36480
rect 38448 36986 38482 37020
rect 38538 36986 38572 37020
rect 38628 36986 38662 37020
rect 38718 36986 38752 37020
rect 38808 36986 38842 37020
rect 38898 36986 38932 37020
rect 38988 36986 39022 37020
rect 38448 36896 38482 36930
rect 38538 36896 38572 36930
rect 38628 36896 38662 36930
rect 38718 36896 38752 36930
rect 38808 36896 38842 36930
rect 38898 36896 38932 36930
rect 38988 36896 39022 36930
rect 38448 36806 38482 36840
rect 38538 36806 38572 36840
rect 38628 36806 38662 36840
rect 38718 36806 38752 36840
rect 38808 36806 38842 36840
rect 38898 36806 38932 36840
rect 38988 36806 39022 36840
rect 38448 36716 38482 36750
rect 38538 36716 38572 36750
rect 38628 36716 38662 36750
rect 38718 36716 38752 36750
rect 38808 36716 38842 36750
rect 38898 36716 38932 36750
rect 38988 36716 39022 36750
rect 38448 36626 38482 36660
rect 38538 36626 38572 36660
rect 38628 36626 38662 36660
rect 38718 36626 38752 36660
rect 38808 36626 38842 36660
rect 38898 36626 38932 36660
rect 38988 36626 39022 36660
rect 38448 36536 38482 36570
rect 38538 36536 38572 36570
rect 38628 36536 38662 36570
rect 38718 36536 38752 36570
rect 38808 36536 38842 36570
rect 38898 36536 38932 36570
rect 38988 36536 39022 36570
rect 38448 36446 38482 36480
rect 38538 36446 38572 36480
rect 38628 36446 38662 36480
rect 38718 36446 38752 36480
rect 38808 36446 38842 36480
rect 38898 36446 38932 36480
rect 38988 36446 39022 36480
rect 14195 33627 14229 33661
rect 14195 33559 14229 33593
rect 14195 33491 14229 33525
rect 14195 33423 14229 33457
rect 14195 33355 14229 33389
rect 14195 33287 14229 33321
rect 14195 33219 14229 33253
rect 14195 33151 14229 33185
rect 14195 33083 14229 33117
rect 14195 33015 14229 33049
rect 14195 32947 14229 32981
rect 14195 32879 14229 32913
rect 14195 32811 14229 32845
rect 14195 32743 14229 32777
rect 14195 32675 14229 32709
rect 14195 32607 14229 32641
rect 14195 32539 14229 32573
rect 14195 32471 14229 32505
rect 14195 32403 14229 32437
rect 14653 33627 14687 33661
rect 14653 33559 14687 33593
rect 14653 33491 14687 33525
rect 14653 33423 14687 33457
rect 14653 33355 14687 33389
rect 14653 33287 14687 33321
rect 14653 33219 14687 33253
rect 14653 33151 14687 33185
rect 14653 33083 14687 33117
rect 14653 33015 14687 33049
rect 14653 32947 14687 32981
rect 14653 32879 14687 32913
rect 14653 32811 14687 32845
rect 14653 32743 14687 32777
rect 14653 32675 14687 32709
rect 14653 32607 14687 32641
rect 14653 32539 14687 32573
rect 14653 32471 14687 32505
rect 14653 32403 14687 32437
rect 15111 33627 15145 33661
rect 15111 33559 15145 33593
rect 15111 33491 15145 33525
rect 15111 33423 15145 33457
rect 15111 33355 15145 33389
rect 15111 33287 15145 33321
rect 15111 33219 15145 33253
rect 15111 33151 15145 33185
rect 15111 33083 15145 33117
rect 15111 33015 15145 33049
rect 15111 32947 15145 32981
rect 15111 32879 15145 32913
rect 15111 32811 15145 32845
rect 15111 32743 15145 32777
rect 15111 32675 15145 32709
rect 15111 32607 15145 32641
rect 15111 32539 15145 32573
rect 15111 32471 15145 32505
rect 15111 32403 15145 32437
rect 15569 33627 15603 33661
rect 15569 33559 15603 33593
rect 15569 33491 15603 33525
rect 15569 33423 15603 33457
rect 15569 33355 15603 33389
rect 15569 33287 15603 33321
rect 15569 33219 15603 33253
rect 15569 33151 15603 33185
rect 15569 33083 15603 33117
rect 15569 33015 15603 33049
rect 15569 32947 15603 32981
rect 15569 32879 15603 32913
rect 15569 32811 15603 32845
rect 15569 32743 15603 32777
rect 15569 32675 15603 32709
rect 15569 32607 15603 32641
rect 15569 32539 15603 32573
rect 15569 32471 15603 32505
rect 15569 32403 15603 32437
rect 16027 33627 16061 33661
rect 16027 33559 16061 33593
rect 16027 33491 16061 33525
rect 16027 33423 16061 33457
rect 16027 33355 16061 33389
rect 16027 33287 16061 33321
rect 16027 33219 16061 33253
rect 16027 33151 16061 33185
rect 16027 33083 16061 33117
rect 16027 33015 16061 33049
rect 16027 32947 16061 32981
rect 16027 32879 16061 32913
rect 16027 32811 16061 32845
rect 16027 32743 16061 32777
rect 16027 32675 16061 32709
rect 16027 32607 16061 32641
rect 16027 32539 16061 32573
rect 16027 32471 16061 32505
rect 16027 32403 16061 32437
rect 16485 33627 16519 33661
rect 16485 33559 16519 33593
rect 16485 33491 16519 33525
rect 16485 33423 16519 33457
rect 16485 33355 16519 33389
rect 16485 33287 16519 33321
rect 16485 33219 16519 33253
rect 16485 33151 16519 33185
rect 16485 33083 16519 33117
rect 16485 33015 16519 33049
rect 16485 32947 16519 32981
rect 16485 32879 16519 32913
rect 16485 32811 16519 32845
rect 16485 32743 16519 32777
rect 16485 32675 16519 32709
rect 16485 32607 16519 32641
rect 16485 32539 16519 32573
rect 16485 32471 16519 32505
rect 16485 32403 16519 32437
rect 16943 33627 16977 33661
rect 16943 33559 16977 33593
rect 16943 33491 16977 33525
rect 16943 33423 16977 33457
rect 16943 33355 16977 33389
rect 16943 33287 16977 33321
rect 16943 33219 16977 33253
rect 16943 33151 16977 33185
rect 16943 33083 16977 33117
rect 16943 33015 16977 33049
rect 16943 32947 16977 32981
rect 16943 32879 16977 32913
rect 16943 32811 16977 32845
rect 16943 32743 16977 32777
rect 16943 32675 16977 32709
rect 16943 32607 16977 32641
rect 16943 32539 16977 32573
rect 16943 32471 16977 32505
rect 16943 32403 16977 32437
rect 17401 33627 17435 33661
rect 17401 33559 17435 33593
rect 17401 33491 17435 33525
rect 17401 33423 17435 33457
rect 17401 33355 17435 33389
rect 17401 33287 17435 33321
rect 17401 33219 17435 33253
rect 17401 33151 17435 33185
rect 17401 33083 17435 33117
rect 17401 33015 17435 33049
rect 17401 32947 17435 32981
rect 17401 32879 17435 32913
rect 17401 32811 17435 32845
rect 17401 32743 17435 32777
rect 17401 32675 17435 32709
rect 17401 32607 17435 32641
rect 17401 32539 17435 32573
rect 17401 32471 17435 32505
rect 17401 32403 17435 32437
rect 17859 33627 17893 33661
rect 17859 33559 17893 33593
rect 17859 33491 17893 33525
rect 17859 33423 17893 33457
rect 17859 33355 17893 33389
rect 17859 33287 17893 33321
rect 17859 33219 17893 33253
rect 17859 33151 17893 33185
rect 17859 33083 17893 33117
rect 17859 33015 17893 33049
rect 17859 32947 17893 32981
rect 17859 32879 17893 32913
rect 17859 32811 17893 32845
rect 17859 32743 17893 32777
rect 17859 32675 17893 32709
rect 17859 32607 17893 32641
rect 17859 32539 17893 32573
rect 17859 32471 17893 32505
rect 17859 32403 17893 32437
rect 18317 33627 18351 33661
rect 18317 33559 18351 33593
rect 18317 33491 18351 33525
rect 18317 33423 18351 33457
rect 18317 33355 18351 33389
rect 18317 33287 18351 33321
rect 18317 33219 18351 33253
rect 18317 33151 18351 33185
rect 18317 33083 18351 33117
rect 18317 33015 18351 33049
rect 18317 32947 18351 32981
rect 18317 32879 18351 32913
rect 18317 32811 18351 32845
rect 18317 32743 18351 32777
rect 18317 32675 18351 32709
rect 18317 32607 18351 32641
rect 18317 32539 18351 32573
rect 18317 32471 18351 32505
rect 18317 32403 18351 32437
rect 18775 33627 18809 33661
rect 18775 33559 18809 33593
rect 18775 33491 18809 33525
rect 18775 33423 18809 33457
rect 18775 33355 18809 33389
rect 18775 33287 18809 33321
rect 18775 33219 18809 33253
rect 18775 33151 18809 33185
rect 18775 33083 18809 33117
rect 18775 33015 18809 33049
rect 18775 32947 18809 32981
rect 18775 32879 18809 32913
rect 18775 32811 18809 32845
rect 18775 32743 18809 32777
rect 18775 32675 18809 32709
rect 18775 32607 18809 32641
rect 18775 32539 18809 32573
rect 18775 32471 18809 32505
rect 18775 32403 18809 32437
rect 19233 33627 19267 33661
rect 19233 33559 19267 33593
rect 19233 33491 19267 33525
rect 19233 33423 19267 33457
rect 19233 33355 19267 33389
rect 19233 33287 19267 33321
rect 19233 33219 19267 33253
rect 19233 33151 19267 33185
rect 19233 33083 19267 33117
rect 19233 33015 19267 33049
rect 19233 32947 19267 32981
rect 19233 32879 19267 32913
rect 19233 32811 19267 32845
rect 19233 32743 19267 32777
rect 19233 32675 19267 32709
rect 19233 32607 19267 32641
rect 19233 32539 19267 32573
rect 19233 32471 19267 32505
rect 19233 32403 19267 32437
rect 19691 33627 19725 33661
rect 19691 33559 19725 33593
rect 19691 33491 19725 33525
rect 19691 33423 19725 33457
rect 19691 33355 19725 33389
rect 19691 33287 19725 33321
rect 19691 33219 19725 33253
rect 19691 33151 19725 33185
rect 19691 33083 19725 33117
rect 19691 33015 19725 33049
rect 19691 32947 19725 32981
rect 19691 32879 19725 32913
rect 19691 32811 19725 32845
rect 19691 32743 19725 32777
rect 19691 32675 19725 32709
rect 19691 32607 19725 32641
rect 19691 32539 19725 32573
rect 19691 32471 19725 32505
rect 19691 32403 19725 32437
rect 20149 33627 20183 33661
rect 20149 33559 20183 33593
rect 20149 33491 20183 33525
rect 20149 33423 20183 33457
rect 20149 33355 20183 33389
rect 20149 33287 20183 33321
rect 20149 33219 20183 33253
rect 20149 33151 20183 33185
rect 20149 33083 20183 33117
rect 20149 33015 20183 33049
rect 20149 32947 20183 32981
rect 20149 32879 20183 32913
rect 20149 32811 20183 32845
rect 20149 32743 20183 32777
rect 20149 32675 20183 32709
rect 20149 32607 20183 32641
rect 20149 32539 20183 32573
rect 20149 32471 20183 32505
rect 20149 32403 20183 32437
rect 20607 33627 20641 33661
rect 20607 33559 20641 33593
rect 20607 33491 20641 33525
rect 20607 33423 20641 33457
rect 20607 33355 20641 33389
rect 20607 33287 20641 33321
rect 20607 33219 20641 33253
rect 20607 33151 20641 33185
rect 20607 33083 20641 33117
rect 20607 33015 20641 33049
rect 20607 32947 20641 32981
rect 20607 32879 20641 32913
rect 20607 32811 20641 32845
rect 20607 32743 20641 32777
rect 20607 32675 20641 32709
rect 20607 32607 20641 32641
rect 20607 32539 20641 32573
rect 20607 32471 20641 32505
rect 20607 32403 20641 32437
rect 21065 33627 21099 33661
rect 21065 33559 21099 33593
rect 21065 33491 21099 33525
rect 21065 33423 21099 33457
rect 21065 33355 21099 33389
rect 21065 33287 21099 33321
rect 21065 33219 21099 33253
rect 21065 33151 21099 33185
rect 21065 33083 21099 33117
rect 21065 33015 21099 33049
rect 21065 32947 21099 32981
rect 21065 32879 21099 32913
rect 21065 32811 21099 32845
rect 21065 32743 21099 32777
rect 21065 32675 21099 32709
rect 21065 32607 21099 32641
rect 21065 32539 21099 32573
rect 21065 32471 21099 32505
rect 21065 32403 21099 32437
rect 21523 33627 21557 33661
rect 21523 33559 21557 33593
rect 21523 33491 21557 33525
rect 21523 33423 21557 33457
rect 21523 33355 21557 33389
rect 21523 33287 21557 33321
rect 21523 33219 21557 33253
rect 21523 33151 21557 33185
rect 21523 33083 21557 33117
rect 21523 33015 21557 33049
rect 21523 32947 21557 32981
rect 21523 32879 21557 32913
rect 21523 32811 21557 32845
rect 21523 32743 21557 32777
rect 21523 32675 21557 32709
rect 21523 32607 21557 32641
rect 21523 32539 21557 32573
rect 21523 32471 21557 32505
rect 21523 32403 21557 32437
rect 21981 33627 22015 33661
rect 21981 33559 22015 33593
rect 21981 33491 22015 33525
rect 21981 33423 22015 33457
rect 21981 33355 22015 33389
rect 21981 33287 22015 33321
rect 21981 33219 22015 33253
rect 21981 33151 22015 33185
rect 21981 33083 22015 33117
rect 21981 33015 22015 33049
rect 21981 32947 22015 32981
rect 21981 32879 22015 32913
rect 21981 32811 22015 32845
rect 21981 32743 22015 32777
rect 21981 32675 22015 32709
rect 21981 32607 22015 32641
rect 21981 32539 22015 32573
rect 21981 32471 22015 32505
rect 21981 32403 22015 32437
rect 22439 33627 22473 33661
rect 22439 33559 22473 33593
rect 22439 33491 22473 33525
rect 22439 33423 22473 33457
rect 22439 33355 22473 33389
rect 22439 33287 22473 33321
rect 22439 33219 22473 33253
rect 22439 33151 22473 33185
rect 22439 33083 22473 33117
rect 22439 33015 22473 33049
rect 22439 32947 22473 32981
rect 22439 32879 22473 32913
rect 22439 32811 22473 32845
rect 22439 32743 22473 32777
rect 22439 32675 22473 32709
rect 22439 32607 22473 32641
rect 22439 32539 22473 32573
rect 22439 32471 22473 32505
rect 22439 32403 22473 32437
rect 22897 33627 22931 33661
rect 22897 33559 22931 33593
rect 22897 33491 22931 33525
rect 22897 33423 22931 33457
rect 22897 33355 22931 33389
rect 22897 33287 22931 33321
rect 22897 33219 22931 33253
rect 22897 33151 22931 33185
rect 22897 33083 22931 33117
rect 22897 33015 22931 33049
rect 22897 32947 22931 32981
rect 22897 32879 22931 32913
rect 22897 32811 22931 32845
rect 22897 32743 22931 32777
rect 22897 32675 22931 32709
rect 22897 32607 22931 32641
rect 22897 32539 22931 32573
rect 22897 32471 22931 32505
rect 22897 32403 22931 32437
rect 23355 33627 23389 33661
rect 23355 33559 23389 33593
rect 23355 33491 23389 33525
rect 23355 33423 23389 33457
rect 23355 33355 23389 33389
rect 23355 33287 23389 33321
rect 23355 33219 23389 33253
rect 23355 33151 23389 33185
rect 23355 33083 23389 33117
rect 23355 33015 23389 33049
rect 23355 32947 23389 32981
rect 23355 32879 23389 32913
rect 23355 32811 23389 32845
rect 23355 32743 23389 32777
rect 23355 32675 23389 32709
rect 23355 32607 23389 32641
rect 23355 32539 23389 32573
rect 23355 32471 23389 32505
rect 23355 32403 23389 32437
rect 23813 33627 23847 33661
rect 23813 33559 23847 33593
rect 23813 33491 23847 33525
rect 23813 33423 23847 33457
rect 23813 33355 23847 33389
rect 23813 33287 23847 33321
rect 23813 33219 23847 33253
rect 23813 33151 23847 33185
rect 23813 33083 23847 33117
rect 23813 33015 23847 33049
rect 23813 32947 23847 32981
rect 23813 32879 23847 32913
rect 23813 32811 23847 32845
rect 23813 32743 23847 32777
rect 23813 32675 23847 32709
rect 23813 32607 23847 32641
rect 23813 32539 23847 32573
rect 23813 32471 23847 32505
rect 23813 32403 23847 32437
rect 24271 33627 24305 33661
rect 24271 33559 24305 33593
rect 24271 33491 24305 33525
rect 24271 33423 24305 33457
rect 24271 33355 24305 33389
rect 24271 33287 24305 33321
rect 24271 33219 24305 33253
rect 24271 33151 24305 33185
rect 24271 33083 24305 33117
rect 24271 33015 24305 33049
rect 24271 32947 24305 32981
rect 24271 32879 24305 32913
rect 24271 32811 24305 32845
rect 24271 32743 24305 32777
rect 24271 32675 24305 32709
rect 24271 32607 24305 32641
rect 24271 32539 24305 32573
rect 24271 32471 24305 32505
rect 24271 32403 24305 32437
rect 24729 33627 24763 33661
rect 24729 33559 24763 33593
rect 24729 33491 24763 33525
rect 24729 33423 24763 33457
rect 24729 33355 24763 33389
rect 24729 33287 24763 33321
rect 24729 33219 24763 33253
rect 24729 33151 24763 33185
rect 24729 33083 24763 33117
rect 24729 33015 24763 33049
rect 24729 32947 24763 32981
rect 24729 32879 24763 32913
rect 24729 32811 24763 32845
rect 24729 32743 24763 32777
rect 24729 32675 24763 32709
rect 24729 32607 24763 32641
rect 24729 32539 24763 32573
rect 24729 32471 24763 32505
rect 24729 32403 24763 32437
rect 25187 33627 25221 33661
rect 25187 33559 25221 33593
rect 25187 33491 25221 33525
rect 25187 33423 25221 33457
rect 25187 33355 25221 33389
rect 25187 33287 25221 33321
rect 25187 33219 25221 33253
rect 25187 33151 25221 33185
rect 25187 33083 25221 33117
rect 25187 33015 25221 33049
rect 25187 32947 25221 32981
rect 25187 32879 25221 32913
rect 25187 32811 25221 32845
rect 25187 32743 25221 32777
rect 25187 32675 25221 32709
rect 25187 32607 25221 32641
rect 25187 32539 25221 32573
rect 25187 32471 25221 32505
rect 25187 32403 25221 32437
rect 25645 33627 25679 33661
rect 25645 33559 25679 33593
rect 25645 33491 25679 33525
rect 25645 33423 25679 33457
rect 25645 33355 25679 33389
rect 25645 33287 25679 33321
rect 25645 33219 25679 33253
rect 25645 33151 25679 33185
rect 25645 33083 25679 33117
rect 25645 33015 25679 33049
rect 25645 32947 25679 32981
rect 25645 32879 25679 32913
rect 25645 32811 25679 32845
rect 25645 32743 25679 32777
rect 25645 32675 25679 32709
rect 25645 32607 25679 32641
rect 25645 32539 25679 32573
rect 25645 32471 25679 32505
rect 25645 32403 25679 32437
rect 26103 33627 26137 33661
rect 26103 33559 26137 33593
rect 26103 33491 26137 33525
rect 26103 33423 26137 33457
rect 26103 33355 26137 33389
rect 26103 33287 26137 33321
rect 26103 33219 26137 33253
rect 26103 33151 26137 33185
rect 26103 33083 26137 33117
rect 26103 33015 26137 33049
rect 26103 32947 26137 32981
rect 26103 32879 26137 32913
rect 26103 32811 26137 32845
rect 26103 32743 26137 32777
rect 26103 32675 26137 32709
rect 26103 32607 26137 32641
rect 26103 32539 26137 32573
rect 26103 32471 26137 32505
rect 26103 32403 26137 32437
rect 26561 33627 26595 33661
rect 26561 33559 26595 33593
rect 26561 33491 26595 33525
rect 26561 33423 26595 33457
rect 26561 33355 26595 33389
rect 26561 33287 26595 33321
rect 26561 33219 26595 33253
rect 26561 33151 26595 33185
rect 26561 33083 26595 33117
rect 26561 33015 26595 33049
rect 26561 32947 26595 32981
rect 26561 32879 26595 32913
rect 26561 32811 26595 32845
rect 26561 32743 26595 32777
rect 26561 32675 26595 32709
rect 26561 32607 26595 32641
rect 26561 32539 26595 32573
rect 26561 32471 26595 32505
rect 26561 32403 26595 32437
rect 27019 33627 27053 33661
rect 27019 33559 27053 33593
rect 27019 33491 27053 33525
rect 27019 33423 27053 33457
rect 27019 33355 27053 33389
rect 27019 33287 27053 33321
rect 27019 33219 27053 33253
rect 27019 33151 27053 33185
rect 27019 33083 27053 33117
rect 27019 33015 27053 33049
rect 27019 32947 27053 32981
rect 27019 32879 27053 32913
rect 27019 32811 27053 32845
rect 27019 32743 27053 32777
rect 27019 32675 27053 32709
rect 27019 32607 27053 32641
rect 27019 32539 27053 32573
rect 27019 32471 27053 32505
rect 27019 32403 27053 32437
rect 27477 33627 27511 33661
rect 27477 33559 27511 33593
rect 27477 33491 27511 33525
rect 27477 33423 27511 33457
rect 27477 33355 27511 33389
rect 27477 33287 27511 33321
rect 27477 33219 27511 33253
rect 27477 33151 27511 33185
rect 27477 33083 27511 33117
rect 27477 33015 27511 33049
rect 27477 32947 27511 32981
rect 27477 32879 27511 32913
rect 27477 32811 27511 32845
rect 27477 32743 27511 32777
rect 27477 32675 27511 32709
rect 27477 32607 27511 32641
rect 27477 32539 27511 32573
rect 27477 32471 27511 32505
rect 27477 32403 27511 32437
rect 27935 33627 27969 33661
rect 27935 33559 27969 33593
rect 27935 33491 27969 33525
rect 27935 33423 27969 33457
rect 27935 33355 27969 33389
rect 27935 33287 27969 33321
rect 27935 33219 27969 33253
rect 27935 33151 27969 33185
rect 27935 33083 27969 33117
rect 27935 33015 27969 33049
rect 27935 32947 27969 32981
rect 27935 32879 27969 32913
rect 27935 32811 27969 32845
rect 27935 32743 27969 32777
rect 27935 32675 27969 32709
rect 27935 32607 27969 32641
rect 27935 32539 27969 32573
rect 27935 32471 27969 32505
rect 27935 32403 27969 32437
rect 28393 33627 28427 33661
rect 28393 33559 28427 33593
rect 28393 33491 28427 33525
rect 28393 33423 28427 33457
rect 28393 33355 28427 33389
rect 28393 33287 28427 33321
rect 28393 33219 28427 33253
rect 28393 33151 28427 33185
rect 28393 33083 28427 33117
rect 28393 33015 28427 33049
rect 28393 32947 28427 32981
rect 28393 32879 28427 32913
rect 28393 32811 28427 32845
rect 28393 32743 28427 32777
rect 28393 32675 28427 32709
rect 28393 32607 28427 32641
rect 28393 32539 28427 32573
rect 28393 32471 28427 32505
rect 28393 32403 28427 32437
rect 28851 33627 28885 33661
rect 28851 33559 28885 33593
rect 28851 33491 28885 33525
rect 28851 33423 28885 33457
rect 28851 33355 28885 33389
rect 28851 33287 28885 33321
rect 28851 33219 28885 33253
rect 28851 33151 28885 33185
rect 28851 33083 28885 33117
rect 28851 33015 28885 33049
rect 28851 32947 28885 32981
rect 28851 32879 28885 32913
rect 28851 32811 28885 32845
rect 28851 32743 28885 32777
rect 28851 32675 28885 32709
rect 28851 32607 28885 32641
rect 28851 32539 28885 32573
rect 28851 32471 28885 32505
rect 28851 32403 28885 32437
rect 29309 33627 29343 33661
rect 29309 33559 29343 33593
rect 29309 33491 29343 33525
rect 29309 33423 29343 33457
rect 29309 33355 29343 33389
rect 29309 33287 29343 33321
rect 29309 33219 29343 33253
rect 29309 33151 29343 33185
rect 29309 33083 29343 33117
rect 29309 33015 29343 33049
rect 29309 32947 29343 32981
rect 29309 32879 29343 32913
rect 29309 32811 29343 32845
rect 29309 32743 29343 32777
rect 29309 32675 29343 32709
rect 29309 32607 29343 32641
rect 29309 32539 29343 32573
rect 29309 32471 29343 32505
rect 29309 32403 29343 32437
rect 29767 33627 29801 33661
rect 29767 33559 29801 33593
rect 29767 33491 29801 33525
rect 29767 33423 29801 33457
rect 29767 33355 29801 33389
rect 29767 33287 29801 33321
rect 29767 33219 29801 33253
rect 29767 33151 29801 33185
rect 29767 33083 29801 33117
rect 29767 33015 29801 33049
rect 29767 32947 29801 32981
rect 29767 32879 29801 32913
rect 29767 32811 29801 32845
rect 29767 32743 29801 32777
rect 29767 32675 29801 32709
rect 29767 32607 29801 32641
rect 29767 32539 29801 32573
rect 29767 32471 29801 32505
rect 29767 32403 29801 32437
rect 30225 33627 30259 33661
rect 30225 33559 30259 33593
rect 30225 33491 30259 33525
rect 30225 33423 30259 33457
rect 30225 33355 30259 33389
rect 30225 33287 30259 33321
rect 30225 33219 30259 33253
rect 30225 33151 30259 33185
rect 30225 33083 30259 33117
rect 30225 33015 30259 33049
rect 30225 32947 30259 32981
rect 30225 32879 30259 32913
rect 30225 32811 30259 32845
rect 30225 32743 30259 32777
rect 30225 32675 30259 32709
rect 30225 32607 30259 32641
rect 30225 32539 30259 32573
rect 30225 32471 30259 32505
rect 30225 32403 30259 32437
rect 30683 33627 30717 33661
rect 30683 33559 30717 33593
rect 30683 33491 30717 33525
rect 30683 33423 30717 33457
rect 30683 33355 30717 33389
rect 30683 33287 30717 33321
rect 30683 33219 30717 33253
rect 30683 33151 30717 33185
rect 30683 33083 30717 33117
rect 30683 33015 30717 33049
rect 30683 32947 30717 32981
rect 30683 32879 30717 32913
rect 30683 32811 30717 32845
rect 30683 32743 30717 32777
rect 30683 32675 30717 32709
rect 30683 32607 30717 32641
rect 30683 32539 30717 32573
rect 30683 32471 30717 32505
rect 30683 32403 30717 32437
rect 31141 33627 31175 33661
rect 31141 33559 31175 33593
rect 31141 33491 31175 33525
rect 31141 33423 31175 33457
rect 31141 33355 31175 33389
rect 31141 33287 31175 33321
rect 31141 33219 31175 33253
rect 31141 33151 31175 33185
rect 31141 33083 31175 33117
rect 31141 33015 31175 33049
rect 31141 32947 31175 32981
rect 31141 32879 31175 32913
rect 31141 32811 31175 32845
rect 31141 32743 31175 32777
rect 31141 32675 31175 32709
rect 31141 32607 31175 32641
rect 31141 32539 31175 32573
rect 31141 32471 31175 32505
rect 31141 32403 31175 32437
rect 31599 33627 31633 33661
rect 31599 33559 31633 33593
rect 31599 33491 31633 33525
rect 31599 33423 31633 33457
rect 31599 33355 31633 33389
rect 31599 33287 31633 33321
rect 31599 33219 31633 33253
rect 31599 33151 31633 33185
rect 31599 33083 31633 33117
rect 31599 33015 31633 33049
rect 31599 32947 31633 32981
rect 31599 32879 31633 32913
rect 31599 32811 31633 32845
rect 31599 32743 31633 32777
rect 31599 32675 31633 32709
rect 31599 32607 31633 32641
rect 31599 32539 31633 32573
rect 31599 32471 31633 32505
rect 31599 32403 31633 32437
rect 32057 33627 32091 33661
rect 32057 33559 32091 33593
rect 32057 33491 32091 33525
rect 32057 33423 32091 33457
rect 32057 33355 32091 33389
rect 32057 33287 32091 33321
rect 32057 33219 32091 33253
rect 32057 33151 32091 33185
rect 32057 33083 32091 33117
rect 32057 33015 32091 33049
rect 32057 32947 32091 32981
rect 32057 32879 32091 32913
rect 32057 32811 32091 32845
rect 32057 32743 32091 32777
rect 32057 32675 32091 32709
rect 32057 32607 32091 32641
rect 32057 32539 32091 32573
rect 32057 32471 32091 32505
rect 32057 32403 32091 32437
rect 32515 33627 32549 33661
rect 32515 33559 32549 33593
rect 32515 33491 32549 33525
rect 32515 33423 32549 33457
rect 32515 33355 32549 33389
rect 32515 33287 32549 33321
rect 32515 33219 32549 33253
rect 32515 33151 32549 33185
rect 32515 33083 32549 33117
rect 32515 33015 32549 33049
rect 32515 32947 32549 32981
rect 32515 32879 32549 32913
rect 32515 32811 32549 32845
rect 32515 32743 32549 32777
rect 32515 32675 32549 32709
rect 32515 32607 32549 32641
rect 32515 32539 32549 32573
rect 32515 32471 32549 32505
rect 32515 32403 32549 32437
rect 32973 33627 33007 33661
rect 32973 33559 33007 33593
rect 32973 33491 33007 33525
rect 32973 33423 33007 33457
rect 32973 33355 33007 33389
rect 32973 33287 33007 33321
rect 32973 33219 33007 33253
rect 32973 33151 33007 33185
rect 32973 33083 33007 33117
rect 32973 33015 33007 33049
rect 32973 32947 33007 32981
rect 32973 32879 33007 32913
rect 32973 32811 33007 32845
rect 32973 32743 33007 32777
rect 32973 32675 33007 32709
rect 32973 32607 33007 32641
rect 32973 32539 33007 32573
rect 32973 32471 33007 32505
rect 32973 32403 33007 32437
rect 33431 33627 33465 33661
rect 33431 33559 33465 33593
rect 33431 33491 33465 33525
rect 33431 33423 33465 33457
rect 33431 33355 33465 33389
rect 33431 33287 33465 33321
rect 33431 33219 33465 33253
rect 33431 33151 33465 33185
rect 33431 33083 33465 33117
rect 33431 33015 33465 33049
rect 33431 32947 33465 32981
rect 33431 32879 33465 32913
rect 33431 32811 33465 32845
rect 33431 32743 33465 32777
rect 33431 32675 33465 32709
rect 33431 32607 33465 32641
rect 33431 32539 33465 32573
rect 33431 32471 33465 32505
rect 33431 32403 33465 32437
rect 33889 33627 33923 33661
rect 33889 33559 33923 33593
rect 33889 33491 33923 33525
rect 33889 33423 33923 33457
rect 33889 33355 33923 33389
rect 33889 33287 33923 33321
rect 33889 33219 33923 33253
rect 33889 33151 33923 33185
rect 33889 33083 33923 33117
rect 33889 33015 33923 33049
rect 33889 32947 33923 32981
rect 33889 32879 33923 32913
rect 33889 32811 33923 32845
rect 33889 32743 33923 32777
rect 33889 32675 33923 32709
rect 33889 32607 33923 32641
rect 33889 32539 33923 32573
rect 33889 32471 33923 32505
rect 33889 32403 33923 32437
rect 34347 33627 34381 33661
rect 34347 33559 34381 33593
rect 34347 33491 34381 33525
rect 34347 33423 34381 33457
rect 34347 33355 34381 33389
rect 34347 33287 34381 33321
rect 34347 33219 34381 33253
rect 34347 33151 34381 33185
rect 34347 33083 34381 33117
rect 34347 33015 34381 33049
rect 34347 32947 34381 32981
rect 34347 32879 34381 32913
rect 34347 32811 34381 32845
rect 34347 32743 34381 32777
rect 34347 32675 34381 32709
rect 34347 32607 34381 32641
rect 34347 32539 34381 32573
rect 34347 32471 34381 32505
rect 34347 32403 34381 32437
rect 34805 33627 34839 33661
rect 34805 33559 34839 33593
rect 34805 33491 34839 33525
rect 34805 33423 34839 33457
rect 34805 33355 34839 33389
rect 34805 33287 34839 33321
rect 34805 33219 34839 33253
rect 34805 33151 34839 33185
rect 34805 33083 34839 33117
rect 34805 33015 34839 33049
rect 34805 32947 34839 32981
rect 34805 32879 34839 32913
rect 34805 32811 34839 32845
rect 34805 32743 34839 32777
rect 34805 32675 34839 32709
rect 34805 32607 34839 32641
rect 34805 32539 34839 32573
rect 34805 32471 34839 32505
rect 34805 32403 34839 32437
rect 35263 33627 35297 33661
rect 35263 33559 35297 33593
rect 35263 33491 35297 33525
rect 35263 33423 35297 33457
rect 35263 33355 35297 33389
rect 35263 33287 35297 33321
rect 35263 33219 35297 33253
rect 35263 33151 35297 33185
rect 35263 33083 35297 33117
rect 35263 33015 35297 33049
rect 35263 32947 35297 32981
rect 35263 32879 35297 32913
rect 35263 32811 35297 32845
rect 35263 32743 35297 32777
rect 35263 32675 35297 32709
rect 35263 32607 35297 32641
rect 35263 32539 35297 32573
rect 35263 32471 35297 32505
rect 35263 32403 35297 32437
rect 35721 33627 35755 33661
rect 35721 33559 35755 33593
rect 35721 33491 35755 33525
rect 35721 33423 35755 33457
rect 35721 33355 35755 33389
rect 35721 33287 35755 33321
rect 35721 33219 35755 33253
rect 35721 33151 35755 33185
rect 35721 33083 35755 33117
rect 35721 33015 35755 33049
rect 35721 32947 35755 32981
rect 35721 32879 35755 32913
rect 35721 32811 35755 32845
rect 35721 32743 35755 32777
rect 35721 32675 35755 32709
rect 35721 32607 35755 32641
rect 35721 32539 35755 32573
rect 35721 32471 35755 32505
rect 35721 32403 35755 32437
rect 36179 33627 36213 33661
rect 36179 33559 36213 33593
rect 36179 33491 36213 33525
rect 36179 33423 36213 33457
rect 36179 33355 36213 33389
rect 36179 33287 36213 33321
rect 36179 33219 36213 33253
rect 36179 33151 36213 33185
rect 36179 33083 36213 33117
rect 36179 33015 36213 33049
rect 36179 32947 36213 32981
rect 36179 32879 36213 32913
rect 36179 32811 36213 32845
rect 36179 32743 36213 32777
rect 36179 32675 36213 32709
rect 36179 32607 36213 32641
rect 36179 32539 36213 32573
rect 36179 32471 36213 32505
rect 36179 32403 36213 32437
rect 36637 33627 36671 33661
rect 36637 33559 36671 33593
rect 36637 33491 36671 33525
rect 36637 33423 36671 33457
rect 36637 33355 36671 33389
rect 36637 33287 36671 33321
rect 36637 33219 36671 33253
rect 36637 33151 36671 33185
rect 36637 33083 36671 33117
rect 36637 33015 36671 33049
rect 36637 32947 36671 32981
rect 36637 32879 36671 32913
rect 36637 32811 36671 32845
rect 36637 32743 36671 32777
rect 36637 32675 36671 32709
rect 36637 32607 36671 32641
rect 36637 32539 36671 32573
rect 36637 32471 36671 32505
rect 36637 32403 36671 32437
rect 37095 33627 37129 33661
rect 37095 33559 37129 33593
rect 37095 33491 37129 33525
rect 37095 33423 37129 33457
rect 37095 33355 37129 33389
rect 37095 33287 37129 33321
rect 37095 33219 37129 33253
rect 37095 33151 37129 33185
rect 37095 33083 37129 33117
rect 37095 33015 37129 33049
rect 37095 32947 37129 32981
rect 37095 32879 37129 32913
rect 37095 32811 37129 32845
rect 37095 32743 37129 32777
rect 37095 32675 37129 32709
rect 37095 32607 37129 32641
rect 37095 32539 37129 32573
rect 37095 32471 37129 32505
rect 37095 32403 37129 32437
rect 37553 33627 37587 33661
rect 37553 33559 37587 33593
rect 37553 33491 37587 33525
rect 37553 33423 37587 33457
rect 37553 33355 37587 33389
rect 37553 33287 37587 33321
rect 37553 33219 37587 33253
rect 37553 33151 37587 33185
rect 37553 33083 37587 33117
rect 37553 33015 37587 33049
rect 37553 32947 37587 32981
rect 37553 32879 37587 32913
rect 37553 32811 37587 32845
rect 37553 32743 37587 32777
rect 37553 32675 37587 32709
rect 37553 32607 37587 32641
rect 37553 32539 37587 32573
rect 37553 32471 37587 32505
rect 37553 32403 37587 32437
rect 38011 33627 38045 33661
rect 38011 33559 38045 33593
rect 38011 33491 38045 33525
rect 38011 33423 38045 33457
rect 38011 33355 38045 33389
rect 38011 33287 38045 33321
rect 38011 33219 38045 33253
rect 38011 33151 38045 33185
rect 38011 33083 38045 33117
rect 38011 33015 38045 33049
rect 38011 32947 38045 32981
rect 38011 32879 38045 32913
rect 38011 32811 38045 32845
rect 38011 32743 38045 32777
rect 38011 32675 38045 32709
rect 38011 32607 38045 32641
rect 38011 32539 38045 32573
rect 38011 32471 38045 32505
rect 38011 32403 38045 32437
rect 38469 33627 38503 33661
rect 38469 33559 38503 33593
rect 38469 33491 38503 33525
rect 38469 33423 38503 33457
rect 38469 33355 38503 33389
rect 38469 33287 38503 33321
rect 38469 33219 38503 33253
rect 38469 33151 38503 33185
rect 38469 33083 38503 33117
rect 38469 33015 38503 33049
rect 38469 32947 38503 32981
rect 38469 32879 38503 32913
rect 38469 32811 38503 32845
rect 38469 32743 38503 32777
rect 38469 32675 38503 32709
rect 38469 32607 38503 32641
rect 38469 32539 38503 32573
rect 38469 32471 38503 32505
rect 38469 32403 38503 32437
rect 38927 33627 38961 33661
rect 38927 33559 38961 33593
rect 38927 33491 38961 33525
rect 38927 33423 38961 33457
rect 38927 33355 38961 33389
rect 38927 33287 38961 33321
rect 38927 33219 38961 33253
rect 38927 33151 38961 33185
rect 38927 33083 38961 33117
rect 38927 33015 38961 33049
rect 38927 32947 38961 32981
rect 38927 32879 38961 32913
rect 38927 32811 38961 32845
rect 38927 32743 38961 32777
rect 38927 32675 38961 32709
rect 38927 32607 38961 32641
rect 38927 32539 38961 32573
rect 38927 32471 38961 32505
rect 38927 32403 38961 32437
rect 39385 33627 39419 33661
rect 39385 33559 39419 33593
rect 39385 33491 39419 33525
rect 39385 33423 39419 33457
rect 39385 33355 39419 33389
rect 39385 33287 39419 33321
rect 39385 33219 39419 33253
rect 39385 33151 39419 33185
rect 39385 33083 39419 33117
rect 39385 33015 39419 33049
rect 39385 32947 39419 32981
rect 39385 32879 39419 32913
rect 39385 32811 39419 32845
rect 39385 32743 39419 32777
rect 39385 32675 39419 32709
rect 39385 32607 39419 32641
rect 39385 32539 39419 32573
rect 39385 32471 39419 32505
rect 39385 32403 39419 32437
rect 39843 33627 39877 33661
rect 39843 33559 39877 33593
rect 39843 33491 39877 33525
rect 39843 33423 39877 33457
rect 39843 33355 39877 33389
rect 39843 33287 39877 33321
rect 39843 33219 39877 33253
rect 39843 33151 39877 33185
rect 39843 33083 39877 33117
rect 39843 33015 39877 33049
rect 39843 32947 39877 32981
rect 39843 32879 39877 32913
rect 39843 32811 39877 32845
rect 39843 32743 39877 32777
rect 39843 32675 39877 32709
rect 39843 32607 39877 32641
rect 39843 32539 39877 32573
rect 39843 32471 39877 32505
rect 39843 32403 39877 32437
rect 40301 33627 40335 33661
rect 40301 33559 40335 33593
rect 40301 33491 40335 33525
rect 40301 33423 40335 33457
rect 40301 33355 40335 33389
rect 40301 33287 40335 33321
rect 40301 33219 40335 33253
rect 40301 33151 40335 33185
rect 40301 33083 40335 33117
rect 40301 33015 40335 33049
rect 40301 32947 40335 32981
rect 40301 32879 40335 32913
rect 40301 32811 40335 32845
rect 40301 32743 40335 32777
rect 40301 32675 40335 32709
rect 40301 32607 40335 32641
rect 40301 32539 40335 32573
rect 40301 32471 40335 32505
rect 40301 32403 40335 32437
rect 40759 33627 40793 33661
rect 40759 33559 40793 33593
rect 40759 33491 40793 33525
rect 40759 33423 40793 33457
rect 40759 33355 40793 33389
rect 40759 33287 40793 33321
rect 40759 33219 40793 33253
rect 40759 33151 40793 33185
rect 40759 33083 40793 33117
rect 40759 33015 40793 33049
rect 40759 32947 40793 32981
rect 40759 32879 40793 32913
rect 40759 32811 40793 32845
rect 40759 32743 40793 32777
rect 40759 32675 40793 32709
rect 40759 32607 40793 32641
rect 40759 32539 40793 32573
rect 40759 32471 40793 32505
rect 40759 32403 40793 32437
rect 41217 33627 41251 33661
rect 41217 33559 41251 33593
rect 41217 33491 41251 33525
rect 41217 33423 41251 33457
rect 41217 33355 41251 33389
rect 41217 33287 41251 33321
rect 41217 33219 41251 33253
rect 41217 33151 41251 33185
rect 41217 33083 41251 33117
rect 41217 33015 41251 33049
rect 41217 32947 41251 32981
rect 41217 32879 41251 32913
rect 41217 32811 41251 32845
rect 41217 32743 41251 32777
rect 41217 32675 41251 32709
rect 41217 32607 41251 32641
rect 41217 32539 41251 32573
rect 41217 32471 41251 32505
rect 41217 32403 41251 32437
rect 41675 33627 41709 33661
rect 41675 33559 41709 33593
rect 41675 33491 41709 33525
rect 41675 33423 41709 33457
rect 41675 33355 41709 33389
rect 41675 33287 41709 33321
rect 41675 33219 41709 33253
rect 41675 33151 41709 33185
rect 41675 33083 41709 33117
rect 41675 33015 41709 33049
rect 41675 32947 41709 32981
rect 41675 32879 41709 32913
rect 41675 32811 41709 32845
rect 41675 32743 41709 32777
rect 41675 32675 41709 32709
rect 41675 32607 41709 32641
rect 41675 32539 41709 32573
rect 41675 32471 41709 32505
rect 41675 32403 41709 32437
rect 6061 29867 6095 29901
rect 6061 29799 6095 29833
rect 6061 29731 6095 29765
rect 6061 29663 6095 29697
rect 6061 29595 6095 29629
rect 6061 29527 6095 29561
rect 6061 29459 6095 29493
rect 6061 29391 6095 29425
rect 6061 29323 6095 29357
rect 6061 29255 6095 29289
rect 6061 29187 6095 29221
rect 6061 29119 6095 29153
rect 6061 29051 6095 29085
rect 6061 28983 6095 29017
rect 6061 28915 6095 28949
rect 6061 28847 6095 28881
rect 6061 28779 6095 28813
rect 6061 28711 6095 28745
rect 6061 28643 6095 28677
rect 6519 29867 6553 29901
rect 6519 29799 6553 29833
rect 6519 29731 6553 29765
rect 6519 29663 6553 29697
rect 6519 29595 6553 29629
rect 6519 29527 6553 29561
rect 6519 29459 6553 29493
rect 6519 29391 6553 29425
rect 6519 29323 6553 29357
rect 6519 29255 6553 29289
rect 6519 29187 6553 29221
rect 6519 29119 6553 29153
rect 6519 29051 6553 29085
rect 6519 28983 6553 29017
rect 6519 28915 6553 28949
rect 6519 28847 6553 28881
rect 6519 28779 6553 28813
rect 6519 28711 6553 28745
rect 6519 28643 6553 28677
rect 6977 29867 7011 29901
rect 6977 29799 7011 29833
rect 6977 29731 7011 29765
rect 6977 29663 7011 29697
rect 6977 29595 7011 29629
rect 6977 29527 7011 29561
rect 6977 29459 7011 29493
rect 6977 29391 7011 29425
rect 6977 29323 7011 29357
rect 6977 29255 7011 29289
rect 6977 29187 7011 29221
rect 6977 29119 7011 29153
rect 6977 29051 7011 29085
rect 6977 28983 7011 29017
rect 6977 28915 7011 28949
rect 6977 28847 7011 28881
rect 6977 28779 7011 28813
rect 6977 28711 7011 28745
rect 6977 28643 7011 28677
rect 7435 29867 7469 29901
rect 7435 29799 7469 29833
rect 7435 29731 7469 29765
rect 7435 29663 7469 29697
rect 7435 29595 7469 29629
rect 7435 29527 7469 29561
rect 7435 29459 7469 29493
rect 7435 29391 7469 29425
rect 7435 29323 7469 29357
rect 7435 29255 7469 29289
rect 7435 29187 7469 29221
rect 7435 29119 7469 29153
rect 7435 29051 7469 29085
rect 7435 28983 7469 29017
rect 7435 28915 7469 28949
rect 7435 28847 7469 28881
rect 7435 28779 7469 28813
rect 7435 28711 7469 28745
rect 7435 28643 7469 28677
rect 7893 29867 7927 29901
rect 7893 29799 7927 29833
rect 7893 29731 7927 29765
rect 7893 29663 7927 29697
rect 7893 29595 7927 29629
rect 7893 29527 7927 29561
rect 7893 29459 7927 29493
rect 7893 29391 7927 29425
rect 7893 29323 7927 29357
rect 7893 29255 7927 29289
rect 7893 29187 7927 29221
rect 7893 29119 7927 29153
rect 7893 29051 7927 29085
rect 7893 28983 7927 29017
rect 7893 28915 7927 28949
rect 7893 28847 7927 28881
rect 7893 28779 7927 28813
rect 7893 28711 7927 28745
rect 7893 28643 7927 28677
rect 8351 29867 8385 29901
rect 8351 29799 8385 29833
rect 8351 29731 8385 29765
rect 8351 29663 8385 29697
rect 8351 29595 8385 29629
rect 8351 29527 8385 29561
rect 8351 29459 8385 29493
rect 8351 29391 8385 29425
rect 8351 29323 8385 29357
rect 8351 29255 8385 29289
rect 8351 29187 8385 29221
rect 8351 29119 8385 29153
rect 8351 29051 8385 29085
rect 8351 28983 8385 29017
rect 8351 28915 8385 28949
rect 8351 28847 8385 28881
rect 8351 28779 8385 28813
rect 8351 28711 8385 28745
rect 8351 28643 8385 28677
rect 8809 29867 8843 29901
rect 8809 29799 8843 29833
rect 8809 29731 8843 29765
rect 8809 29663 8843 29697
rect 8809 29595 8843 29629
rect 8809 29527 8843 29561
rect 8809 29459 8843 29493
rect 8809 29391 8843 29425
rect 8809 29323 8843 29357
rect 8809 29255 8843 29289
rect 8809 29187 8843 29221
rect 8809 29119 8843 29153
rect 8809 29051 8843 29085
rect 8809 28983 8843 29017
rect 8809 28915 8843 28949
rect 8809 28847 8843 28881
rect 8809 28779 8843 28813
rect 8809 28711 8843 28745
rect 8809 28643 8843 28677
rect 9267 29867 9301 29901
rect 9267 29799 9301 29833
rect 9267 29731 9301 29765
rect 9267 29663 9301 29697
rect 9267 29595 9301 29629
rect 9267 29527 9301 29561
rect 9267 29459 9301 29493
rect 9267 29391 9301 29425
rect 9267 29323 9301 29357
rect 9267 29255 9301 29289
rect 9267 29187 9301 29221
rect 9267 29119 9301 29153
rect 9267 29051 9301 29085
rect 9267 28983 9301 29017
rect 9267 28915 9301 28949
rect 9267 28847 9301 28881
rect 9267 28779 9301 28813
rect 9267 28711 9301 28745
rect 9267 28643 9301 28677
rect 9725 29867 9759 29901
rect 9725 29799 9759 29833
rect 9725 29731 9759 29765
rect 9725 29663 9759 29697
rect 9725 29595 9759 29629
rect 9725 29527 9759 29561
rect 9725 29459 9759 29493
rect 9725 29391 9759 29425
rect 9725 29323 9759 29357
rect 9725 29255 9759 29289
rect 9725 29187 9759 29221
rect 9725 29119 9759 29153
rect 9725 29051 9759 29085
rect 9725 28983 9759 29017
rect 9725 28915 9759 28949
rect 9725 28847 9759 28881
rect 9725 28779 9759 28813
rect 9725 28711 9759 28745
rect 9725 28643 9759 28677
rect 10183 29867 10217 29901
rect 10183 29799 10217 29833
rect 10183 29731 10217 29765
rect 10183 29663 10217 29697
rect 10183 29595 10217 29629
rect 10183 29527 10217 29561
rect 10183 29459 10217 29493
rect 10183 29391 10217 29425
rect 10183 29323 10217 29357
rect 10183 29255 10217 29289
rect 10183 29187 10217 29221
rect 10183 29119 10217 29153
rect 10183 29051 10217 29085
rect 10183 28983 10217 29017
rect 10183 28915 10217 28949
rect 10183 28847 10217 28881
rect 10183 28779 10217 28813
rect 10183 28711 10217 28745
rect 10183 28643 10217 28677
rect 10641 29867 10675 29901
rect 10641 29799 10675 29833
rect 10641 29731 10675 29765
rect 10641 29663 10675 29697
rect 10641 29595 10675 29629
rect 10641 29527 10675 29561
rect 10641 29459 10675 29493
rect 10641 29391 10675 29425
rect 10641 29323 10675 29357
rect 10641 29255 10675 29289
rect 10641 29187 10675 29221
rect 10641 29119 10675 29153
rect 10641 29051 10675 29085
rect 10641 28983 10675 29017
rect 10641 28915 10675 28949
rect 10641 28847 10675 28881
rect 10641 28779 10675 28813
rect 10641 28711 10675 28745
rect 10641 28643 10675 28677
rect 11099 29867 11133 29901
rect 11099 29799 11133 29833
rect 11099 29731 11133 29765
rect 11099 29663 11133 29697
rect 11099 29595 11133 29629
rect 11099 29527 11133 29561
rect 11099 29459 11133 29493
rect 11099 29391 11133 29425
rect 11099 29323 11133 29357
rect 11099 29255 11133 29289
rect 11099 29187 11133 29221
rect 11099 29119 11133 29153
rect 11099 29051 11133 29085
rect 11099 28983 11133 29017
rect 11099 28915 11133 28949
rect 11099 28847 11133 28881
rect 11099 28779 11133 28813
rect 11099 28711 11133 28745
rect 11099 28643 11133 28677
rect 11557 29867 11591 29901
rect 11557 29799 11591 29833
rect 11557 29731 11591 29765
rect 11557 29663 11591 29697
rect 11557 29595 11591 29629
rect 11557 29527 11591 29561
rect 11557 29459 11591 29493
rect 11557 29391 11591 29425
rect 11557 29323 11591 29357
rect 11557 29255 11591 29289
rect 11557 29187 11591 29221
rect 11557 29119 11591 29153
rect 11557 29051 11591 29085
rect 11557 28983 11591 29017
rect 11557 28915 11591 28949
rect 11557 28847 11591 28881
rect 11557 28779 11591 28813
rect 11557 28711 11591 28745
rect 11557 28643 11591 28677
rect 12015 29867 12049 29901
rect 12015 29799 12049 29833
rect 12015 29731 12049 29765
rect 12015 29663 12049 29697
rect 12015 29595 12049 29629
rect 12015 29527 12049 29561
rect 12015 29459 12049 29493
rect 12015 29391 12049 29425
rect 12015 29323 12049 29357
rect 12015 29255 12049 29289
rect 12015 29187 12049 29221
rect 12015 29119 12049 29153
rect 12015 29051 12049 29085
rect 12015 28983 12049 29017
rect 12015 28915 12049 28949
rect 12015 28847 12049 28881
rect 12015 28779 12049 28813
rect 12015 28711 12049 28745
rect 12015 28643 12049 28677
rect 12473 29867 12507 29901
rect 12473 29799 12507 29833
rect 12473 29731 12507 29765
rect 12473 29663 12507 29697
rect 12473 29595 12507 29629
rect 12473 29527 12507 29561
rect 12473 29459 12507 29493
rect 12473 29391 12507 29425
rect 12473 29323 12507 29357
rect 12473 29255 12507 29289
rect 12473 29187 12507 29221
rect 12473 29119 12507 29153
rect 12473 29051 12507 29085
rect 12473 28983 12507 29017
rect 12473 28915 12507 28949
rect 12473 28847 12507 28881
rect 12473 28779 12507 28813
rect 12473 28711 12507 28745
rect 12473 28643 12507 28677
rect 12931 29867 12965 29901
rect 12931 29799 12965 29833
rect 12931 29731 12965 29765
rect 12931 29663 12965 29697
rect 12931 29595 12965 29629
rect 12931 29527 12965 29561
rect 12931 29459 12965 29493
rect 12931 29391 12965 29425
rect 12931 29323 12965 29357
rect 12931 29255 12965 29289
rect 12931 29187 12965 29221
rect 12931 29119 12965 29153
rect 12931 29051 12965 29085
rect 12931 28983 12965 29017
rect 12931 28915 12965 28949
rect 12931 28847 12965 28881
rect 12931 28779 12965 28813
rect 12931 28711 12965 28745
rect 12931 28643 12965 28677
rect 13389 29867 13423 29901
rect 13389 29799 13423 29833
rect 13389 29731 13423 29765
rect 13389 29663 13423 29697
rect 13389 29595 13423 29629
rect 13389 29527 13423 29561
rect 13389 29459 13423 29493
rect 13389 29391 13423 29425
rect 13389 29323 13423 29357
rect 13389 29255 13423 29289
rect 13389 29187 13423 29221
rect 13389 29119 13423 29153
rect 13389 29051 13423 29085
rect 13389 28983 13423 29017
rect 13389 28915 13423 28949
rect 13389 28847 13423 28881
rect 13389 28779 13423 28813
rect 13389 28711 13423 28745
rect 13389 28643 13423 28677
rect 13847 29867 13881 29901
rect 13847 29799 13881 29833
rect 13847 29731 13881 29765
rect 13847 29663 13881 29697
rect 13847 29595 13881 29629
rect 13847 29527 13881 29561
rect 13847 29459 13881 29493
rect 13847 29391 13881 29425
rect 13847 29323 13881 29357
rect 13847 29255 13881 29289
rect 13847 29187 13881 29221
rect 13847 29119 13881 29153
rect 13847 29051 13881 29085
rect 13847 28983 13881 29017
rect 13847 28915 13881 28949
rect 13847 28847 13881 28881
rect 13847 28779 13881 28813
rect 13847 28711 13881 28745
rect 13847 28643 13881 28677
rect 14305 29867 14339 29901
rect 14305 29799 14339 29833
rect 14305 29731 14339 29765
rect 14305 29663 14339 29697
rect 14305 29595 14339 29629
rect 14305 29527 14339 29561
rect 14305 29459 14339 29493
rect 14305 29391 14339 29425
rect 14305 29323 14339 29357
rect 14305 29255 14339 29289
rect 14305 29187 14339 29221
rect 14305 29119 14339 29153
rect 14305 29051 14339 29085
rect 14305 28983 14339 29017
rect 14305 28915 14339 28949
rect 14305 28847 14339 28881
rect 14305 28779 14339 28813
rect 14305 28711 14339 28745
rect 14305 28643 14339 28677
rect 14763 29867 14797 29901
rect 14763 29799 14797 29833
rect 14763 29731 14797 29765
rect 14763 29663 14797 29697
rect 14763 29595 14797 29629
rect 14763 29527 14797 29561
rect 14763 29459 14797 29493
rect 14763 29391 14797 29425
rect 14763 29323 14797 29357
rect 14763 29255 14797 29289
rect 14763 29187 14797 29221
rect 14763 29119 14797 29153
rect 14763 29051 14797 29085
rect 14763 28983 14797 29017
rect 14763 28915 14797 28949
rect 14763 28847 14797 28881
rect 14763 28779 14797 28813
rect 14763 28711 14797 28745
rect 14763 28643 14797 28677
rect 15221 29867 15255 29901
rect 15221 29799 15255 29833
rect 15221 29731 15255 29765
rect 15221 29663 15255 29697
rect 15221 29595 15255 29629
rect 15221 29527 15255 29561
rect 15221 29459 15255 29493
rect 15221 29391 15255 29425
rect 15221 29323 15255 29357
rect 15221 29255 15255 29289
rect 15221 29187 15255 29221
rect 15221 29119 15255 29153
rect 15221 29051 15255 29085
rect 15221 28983 15255 29017
rect 15221 28915 15255 28949
rect 15221 28847 15255 28881
rect 15221 28779 15255 28813
rect 15221 28711 15255 28745
rect 15221 28643 15255 28677
rect 15679 29867 15713 29901
rect 15679 29799 15713 29833
rect 15679 29731 15713 29765
rect 15679 29663 15713 29697
rect 15679 29595 15713 29629
rect 15679 29527 15713 29561
rect 15679 29459 15713 29493
rect 15679 29391 15713 29425
rect 15679 29323 15713 29357
rect 15679 29255 15713 29289
rect 15679 29187 15713 29221
rect 15679 29119 15713 29153
rect 15679 29051 15713 29085
rect 15679 28983 15713 29017
rect 15679 28915 15713 28949
rect 15679 28847 15713 28881
rect 15679 28779 15713 28813
rect 15679 28711 15713 28745
rect 15679 28643 15713 28677
rect 16137 29867 16171 29901
rect 16137 29799 16171 29833
rect 16137 29731 16171 29765
rect 16137 29663 16171 29697
rect 16137 29595 16171 29629
rect 16137 29527 16171 29561
rect 16137 29459 16171 29493
rect 16137 29391 16171 29425
rect 16137 29323 16171 29357
rect 16137 29255 16171 29289
rect 16137 29187 16171 29221
rect 16137 29119 16171 29153
rect 16137 29051 16171 29085
rect 16137 28983 16171 29017
rect 16137 28915 16171 28949
rect 16137 28847 16171 28881
rect 16137 28779 16171 28813
rect 16137 28711 16171 28745
rect 16137 28643 16171 28677
rect 16595 29867 16629 29901
rect 16595 29799 16629 29833
rect 16595 29731 16629 29765
rect 16595 29663 16629 29697
rect 16595 29595 16629 29629
rect 16595 29527 16629 29561
rect 16595 29459 16629 29493
rect 16595 29391 16629 29425
rect 16595 29323 16629 29357
rect 16595 29255 16629 29289
rect 16595 29187 16629 29221
rect 16595 29119 16629 29153
rect 16595 29051 16629 29085
rect 16595 28983 16629 29017
rect 16595 28915 16629 28949
rect 16595 28847 16629 28881
rect 16595 28779 16629 28813
rect 16595 28711 16629 28745
rect 16595 28643 16629 28677
rect 17053 29867 17087 29901
rect 17053 29799 17087 29833
rect 17053 29731 17087 29765
rect 17053 29663 17087 29697
rect 17053 29595 17087 29629
rect 17053 29527 17087 29561
rect 17053 29459 17087 29493
rect 17053 29391 17087 29425
rect 17053 29323 17087 29357
rect 17053 29255 17087 29289
rect 17053 29187 17087 29221
rect 17053 29119 17087 29153
rect 17053 29051 17087 29085
rect 17053 28983 17087 29017
rect 17053 28915 17087 28949
rect 17053 28847 17087 28881
rect 17053 28779 17087 28813
rect 17053 28711 17087 28745
rect 17053 28643 17087 28677
rect 17511 29867 17545 29901
rect 17511 29799 17545 29833
rect 17511 29731 17545 29765
rect 17511 29663 17545 29697
rect 17511 29595 17545 29629
rect 17511 29527 17545 29561
rect 17511 29459 17545 29493
rect 17511 29391 17545 29425
rect 17511 29323 17545 29357
rect 17511 29255 17545 29289
rect 17511 29187 17545 29221
rect 17511 29119 17545 29153
rect 17511 29051 17545 29085
rect 17511 28983 17545 29017
rect 17511 28915 17545 28949
rect 17511 28847 17545 28881
rect 17511 28779 17545 28813
rect 17511 28711 17545 28745
rect 17511 28643 17545 28677
rect 17969 29867 18003 29901
rect 17969 29799 18003 29833
rect 17969 29731 18003 29765
rect 17969 29663 18003 29697
rect 17969 29595 18003 29629
rect 17969 29527 18003 29561
rect 17969 29459 18003 29493
rect 17969 29391 18003 29425
rect 17969 29323 18003 29357
rect 17969 29255 18003 29289
rect 17969 29187 18003 29221
rect 17969 29119 18003 29153
rect 17969 29051 18003 29085
rect 17969 28983 18003 29017
rect 17969 28915 18003 28949
rect 17969 28847 18003 28881
rect 17969 28779 18003 28813
rect 17969 28711 18003 28745
rect 17969 28643 18003 28677
rect 18427 29867 18461 29901
rect 18427 29799 18461 29833
rect 18427 29731 18461 29765
rect 18427 29663 18461 29697
rect 18427 29595 18461 29629
rect 18427 29527 18461 29561
rect 18427 29459 18461 29493
rect 18427 29391 18461 29425
rect 18427 29323 18461 29357
rect 18427 29255 18461 29289
rect 18427 29187 18461 29221
rect 18427 29119 18461 29153
rect 18427 29051 18461 29085
rect 18427 28983 18461 29017
rect 18427 28915 18461 28949
rect 18427 28847 18461 28881
rect 18427 28779 18461 28813
rect 18427 28711 18461 28745
rect 18427 28643 18461 28677
rect 18885 29867 18919 29901
rect 18885 29799 18919 29833
rect 18885 29731 18919 29765
rect 18885 29663 18919 29697
rect 18885 29595 18919 29629
rect 18885 29527 18919 29561
rect 18885 29459 18919 29493
rect 18885 29391 18919 29425
rect 18885 29323 18919 29357
rect 18885 29255 18919 29289
rect 18885 29187 18919 29221
rect 18885 29119 18919 29153
rect 18885 29051 18919 29085
rect 18885 28983 18919 29017
rect 18885 28915 18919 28949
rect 18885 28847 18919 28881
rect 18885 28779 18919 28813
rect 18885 28711 18919 28745
rect 18885 28643 18919 28677
rect 19343 29867 19377 29901
rect 19343 29799 19377 29833
rect 19343 29731 19377 29765
rect 19343 29663 19377 29697
rect 19343 29595 19377 29629
rect 19343 29527 19377 29561
rect 19343 29459 19377 29493
rect 19343 29391 19377 29425
rect 19343 29323 19377 29357
rect 19343 29255 19377 29289
rect 19343 29187 19377 29221
rect 19343 29119 19377 29153
rect 19343 29051 19377 29085
rect 19343 28983 19377 29017
rect 19343 28915 19377 28949
rect 19343 28847 19377 28881
rect 19343 28779 19377 28813
rect 19343 28711 19377 28745
rect 19343 28643 19377 28677
rect 19801 29867 19835 29901
rect 19801 29799 19835 29833
rect 19801 29731 19835 29765
rect 19801 29663 19835 29697
rect 19801 29595 19835 29629
rect 19801 29527 19835 29561
rect 19801 29459 19835 29493
rect 19801 29391 19835 29425
rect 19801 29323 19835 29357
rect 19801 29255 19835 29289
rect 19801 29187 19835 29221
rect 19801 29119 19835 29153
rect 19801 29051 19835 29085
rect 19801 28983 19835 29017
rect 19801 28915 19835 28949
rect 19801 28847 19835 28881
rect 19801 28779 19835 28813
rect 19801 28711 19835 28745
rect 19801 28643 19835 28677
rect 20259 29867 20293 29901
rect 20259 29799 20293 29833
rect 20259 29731 20293 29765
rect 20259 29663 20293 29697
rect 20259 29595 20293 29629
rect 20259 29527 20293 29561
rect 20259 29459 20293 29493
rect 20259 29391 20293 29425
rect 20259 29323 20293 29357
rect 20259 29255 20293 29289
rect 20259 29187 20293 29221
rect 20259 29119 20293 29153
rect 20259 29051 20293 29085
rect 20259 28983 20293 29017
rect 20259 28915 20293 28949
rect 20259 28847 20293 28881
rect 20259 28779 20293 28813
rect 20259 28711 20293 28745
rect 20259 28643 20293 28677
rect 20717 29867 20751 29901
rect 20717 29799 20751 29833
rect 20717 29731 20751 29765
rect 20717 29663 20751 29697
rect 20717 29595 20751 29629
rect 20717 29527 20751 29561
rect 20717 29459 20751 29493
rect 20717 29391 20751 29425
rect 20717 29323 20751 29357
rect 20717 29255 20751 29289
rect 20717 29187 20751 29221
rect 20717 29119 20751 29153
rect 20717 29051 20751 29085
rect 20717 28983 20751 29017
rect 20717 28915 20751 28949
rect 20717 28847 20751 28881
rect 20717 28779 20751 28813
rect 20717 28711 20751 28745
rect 20717 28643 20751 28677
rect 21175 29867 21209 29901
rect 21175 29799 21209 29833
rect 21175 29731 21209 29765
rect 21175 29663 21209 29697
rect 21175 29595 21209 29629
rect 21175 29527 21209 29561
rect 21175 29459 21209 29493
rect 21175 29391 21209 29425
rect 21175 29323 21209 29357
rect 21175 29255 21209 29289
rect 21175 29187 21209 29221
rect 21175 29119 21209 29153
rect 21175 29051 21209 29085
rect 21175 28983 21209 29017
rect 21175 28915 21209 28949
rect 21175 28847 21209 28881
rect 21175 28779 21209 28813
rect 21175 28711 21209 28745
rect 21175 28643 21209 28677
rect 21633 29867 21667 29901
rect 21633 29799 21667 29833
rect 21633 29731 21667 29765
rect 21633 29663 21667 29697
rect 21633 29595 21667 29629
rect 21633 29527 21667 29561
rect 21633 29459 21667 29493
rect 21633 29391 21667 29425
rect 21633 29323 21667 29357
rect 21633 29255 21667 29289
rect 21633 29187 21667 29221
rect 21633 29119 21667 29153
rect 21633 29051 21667 29085
rect 21633 28983 21667 29017
rect 21633 28915 21667 28949
rect 21633 28847 21667 28881
rect 21633 28779 21667 28813
rect 21633 28711 21667 28745
rect 21633 28643 21667 28677
rect 22091 29867 22125 29901
rect 22091 29799 22125 29833
rect 22091 29731 22125 29765
rect 22091 29663 22125 29697
rect 22091 29595 22125 29629
rect 22091 29527 22125 29561
rect 22091 29459 22125 29493
rect 22091 29391 22125 29425
rect 22091 29323 22125 29357
rect 22091 29255 22125 29289
rect 22091 29187 22125 29221
rect 22091 29119 22125 29153
rect 22091 29051 22125 29085
rect 22091 28983 22125 29017
rect 22091 28915 22125 28949
rect 22091 28847 22125 28881
rect 22091 28779 22125 28813
rect 22091 28711 22125 28745
rect 22091 28643 22125 28677
rect 22549 29867 22583 29901
rect 22549 29799 22583 29833
rect 22549 29731 22583 29765
rect 22549 29663 22583 29697
rect 22549 29595 22583 29629
rect 22549 29527 22583 29561
rect 22549 29459 22583 29493
rect 22549 29391 22583 29425
rect 22549 29323 22583 29357
rect 22549 29255 22583 29289
rect 22549 29187 22583 29221
rect 22549 29119 22583 29153
rect 22549 29051 22583 29085
rect 22549 28983 22583 29017
rect 22549 28915 22583 28949
rect 22549 28847 22583 28881
rect 22549 28779 22583 28813
rect 22549 28711 22583 28745
rect 22549 28643 22583 28677
rect 23007 29867 23041 29901
rect 23007 29799 23041 29833
rect 23007 29731 23041 29765
rect 23007 29663 23041 29697
rect 23007 29595 23041 29629
rect 23007 29527 23041 29561
rect 23007 29459 23041 29493
rect 23007 29391 23041 29425
rect 23007 29323 23041 29357
rect 23007 29255 23041 29289
rect 23007 29187 23041 29221
rect 23007 29119 23041 29153
rect 23007 29051 23041 29085
rect 23007 28983 23041 29017
rect 23007 28915 23041 28949
rect 23007 28847 23041 28881
rect 23007 28779 23041 28813
rect 23007 28711 23041 28745
rect 23007 28643 23041 28677
rect 23465 29867 23499 29901
rect 23465 29799 23499 29833
rect 23465 29731 23499 29765
rect 23465 29663 23499 29697
rect 23465 29595 23499 29629
rect 23465 29527 23499 29561
rect 23465 29459 23499 29493
rect 23465 29391 23499 29425
rect 23465 29323 23499 29357
rect 23465 29255 23499 29289
rect 23465 29187 23499 29221
rect 23465 29119 23499 29153
rect 23465 29051 23499 29085
rect 23465 28983 23499 29017
rect 23465 28915 23499 28949
rect 23465 28847 23499 28881
rect 23465 28779 23499 28813
rect 23465 28711 23499 28745
rect 23465 28643 23499 28677
rect 23923 29867 23957 29901
rect 23923 29799 23957 29833
rect 23923 29731 23957 29765
rect 23923 29663 23957 29697
rect 23923 29595 23957 29629
rect 23923 29527 23957 29561
rect 23923 29459 23957 29493
rect 23923 29391 23957 29425
rect 23923 29323 23957 29357
rect 23923 29255 23957 29289
rect 23923 29187 23957 29221
rect 23923 29119 23957 29153
rect 23923 29051 23957 29085
rect 23923 28983 23957 29017
rect 23923 28915 23957 28949
rect 23923 28847 23957 28881
rect 23923 28779 23957 28813
rect 23923 28711 23957 28745
rect 23923 28643 23957 28677
rect 24381 29867 24415 29901
rect 24381 29799 24415 29833
rect 24381 29731 24415 29765
rect 24381 29663 24415 29697
rect 24381 29595 24415 29629
rect 24381 29527 24415 29561
rect 24381 29459 24415 29493
rect 24381 29391 24415 29425
rect 24381 29323 24415 29357
rect 24381 29255 24415 29289
rect 24381 29187 24415 29221
rect 24381 29119 24415 29153
rect 24381 29051 24415 29085
rect 24381 28983 24415 29017
rect 24381 28915 24415 28949
rect 24381 28847 24415 28881
rect 24381 28779 24415 28813
rect 24381 28711 24415 28745
rect 24381 28643 24415 28677
rect 24839 29867 24873 29901
rect 24839 29799 24873 29833
rect 24839 29731 24873 29765
rect 24839 29663 24873 29697
rect 24839 29595 24873 29629
rect 24839 29527 24873 29561
rect 24839 29459 24873 29493
rect 24839 29391 24873 29425
rect 24839 29323 24873 29357
rect 24839 29255 24873 29289
rect 24839 29187 24873 29221
rect 24839 29119 24873 29153
rect 24839 29051 24873 29085
rect 24839 28983 24873 29017
rect 24839 28915 24873 28949
rect 24839 28847 24873 28881
rect 24839 28779 24873 28813
rect 24839 28711 24873 28745
rect 24839 28643 24873 28677
rect 25297 29867 25331 29901
rect 25297 29799 25331 29833
rect 25297 29731 25331 29765
rect 25297 29663 25331 29697
rect 25297 29595 25331 29629
rect 25297 29527 25331 29561
rect 25297 29459 25331 29493
rect 25297 29391 25331 29425
rect 25297 29323 25331 29357
rect 25297 29255 25331 29289
rect 25297 29187 25331 29221
rect 25297 29119 25331 29153
rect 25297 29051 25331 29085
rect 25297 28983 25331 29017
rect 25297 28915 25331 28949
rect 25297 28847 25331 28881
rect 25297 28779 25331 28813
rect 25297 28711 25331 28745
rect 25297 28643 25331 28677
rect 25755 29867 25789 29901
rect 25755 29799 25789 29833
rect 25755 29731 25789 29765
rect 25755 29663 25789 29697
rect 25755 29595 25789 29629
rect 25755 29527 25789 29561
rect 25755 29459 25789 29493
rect 25755 29391 25789 29425
rect 25755 29323 25789 29357
rect 25755 29255 25789 29289
rect 25755 29187 25789 29221
rect 25755 29119 25789 29153
rect 25755 29051 25789 29085
rect 25755 28983 25789 29017
rect 25755 28915 25789 28949
rect 25755 28847 25789 28881
rect 25755 28779 25789 28813
rect 25755 28711 25789 28745
rect 25755 28643 25789 28677
rect 26213 29867 26247 29901
rect 26213 29799 26247 29833
rect 26213 29731 26247 29765
rect 26213 29663 26247 29697
rect 26213 29595 26247 29629
rect 26213 29527 26247 29561
rect 26213 29459 26247 29493
rect 26213 29391 26247 29425
rect 26213 29323 26247 29357
rect 26213 29255 26247 29289
rect 26213 29187 26247 29221
rect 26213 29119 26247 29153
rect 26213 29051 26247 29085
rect 26213 28983 26247 29017
rect 26213 28915 26247 28949
rect 26213 28847 26247 28881
rect 26213 28779 26247 28813
rect 26213 28711 26247 28745
rect 26213 28643 26247 28677
rect 26671 29867 26705 29901
rect 26671 29799 26705 29833
rect 26671 29731 26705 29765
rect 26671 29663 26705 29697
rect 26671 29595 26705 29629
rect 26671 29527 26705 29561
rect 26671 29459 26705 29493
rect 26671 29391 26705 29425
rect 26671 29323 26705 29357
rect 26671 29255 26705 29289
rect 26671 29187 26705 29221
rect 26671 29119 26705 29153
rect 26671 29051 26705 29085
rect 26671 28983 26705 29017
rect 26671 28915 26705 28949
rect 26671 28847 26705 28881
rect 26671 28779 26705 28813
rect 26671 28711 26705 28745
rect 26671 28643 26705 28677
rect 27129 29867 27163 29901
rect 27129 29799 27163 29833
rect 27129 29731 27163 29765
rect 27129 29663 27163 29697
rect 27129 29595 27163 29629
rect 27129 29527 27163 29561
rect 27129 29459 27163 29493
rect 27129 29391 27163 29425
rect 27129 29323 27163 29357
rect 27129 29255 27163 29289
rect 27129 29187 27163 29221
rect 27129 29119 27163 29153
rect 27129 29051 27163 29085
rect 27129 28983 27163 29017
rect 27129 28915 27163 28949
rect 27129 28847 27163 28881
rect 27129 28779 27163 28813
rect 27129 28711 27163 28745
rect 27129 28643 27163 28677
rect 27587 29867 27621 29901
rect 27587 29799 27621 29833
rect 27587 29731 27621 29765
rect 27587 29663 27621 29697
rect 27587 29595 27621 29629
rect 27587 29527 27621 29561
rect 27587 29459 27621 29493
rect 27587 29391 27621 29425
rect 27587 29323 27621 29357
rect 27587 29255 27621 29289
rect 27587 29187 27621 29221
rect 27587 29119 27621 29153
rect 27587 29051 27621 29085
rect 27587 28983 27621 29017
rect 27587 28915 27621 28949
rect 27587 28847 27621 28881
rect 27587 28779 27621 28813
rect 27587 28711 27621 28745
rect 27587 28643 27621 28677
rect 28045 29867 28079 29901
rect 28045 29799 28079 29833
rect 28045 29731 28079 29765
rect 28045 29663 28079 29697
rect 28045 29595 28079 29629
rect 28045 29527 28079 29561
rect 28045 29459 28079 29493
rect 28045 29391 28079 29425
rect 28045 29323 28079 29357
rect 28045 29255 28079 29289
rect 28045 29187 28079 29221
rect 28045 29119 28079 29153
rect 28045 29051 28079 29085
rect 28045 28983 28079 29017
rect 28045 28915 28079 28949
rect 28045 28847 28079 28881
rect 28045 28779 28079 28813
rect 28045 28711 28079 28745
rect 28045 28643 28079 28677
rect 28503 29867 28537 29901
rect 28503 29799 28537 29833
rect 28503 29731 28537 29765
rect 28503 29663 28537 29697
rect 28503 29595 28537 29629
rect 28503 29527 28537 29561
rect 28503 29459 28537 29493
rect 28503 29391 28537 29425
rect 28503 29323 28537 29357
rect 28503 29255 28537 29289
rect 28503 29187 28537 29221
rect 28503 29119 28537 29153
rect 28503 29051 28537 29085
rect 28503 28983 28537 29017
rect 28503 28915 28537 28949
rect 28503 28847 28537 28881
rect 28503 28779 28537 28813
rect 28503 28711 28537 28745
rect 28503 28643 28537 28677
rect 28961 29867 28995 29901
rect 28961 29799 28995 29833
rect 28961 29731 28995 29765
rect 28961 29663 28995 29697
rect 28961 29595 28995 29629
rect 28961 29527 28995 29561
rect 28961 29459 28995 29493
rect 28961 29391 28995 29425
rect 28961 29323 28995 29357
rect 28961 29255 28995 29289
rect 28961 29187 28995 29221
rect 28961 29119 28995 29153
rect 28961 29051 28995 29085
rect 28961 28983 28995 29017
rect 28961 28915 28995 28949
rect 28961 28847 28995 28881
rect 28961 28779 28995 28813
rect 28961 28711 28995 28745
rect 28961 28643 28995 28677
rect 29419 29867 29453 29901
rect 29419 29799 29453 29833
rect 29419 29731 29453 29765
rect 29419 29663 29453 29697
rect 29419 29595 29453 29629
rect 29419 29527 29453 29561
rect 29419 29459 29453 29493
rect 29419 29391 29453 29425
rect 29419 29323 29453 29357
rect 29419 29255 29453 29289
rect 29419 29187 29453 29221
rect 29419 29119 29453 29153
rect 29419 29051 29453 29085
rect 29419 28983 29453 29017
rect 29419 28915 29453 28949
rect 29419 28847 29453 28881
rect 29419 28779 29453 28813
rect 29419 28711 29453 28745
rect 29419 28643 29453 28677
rect 29877 29867 29911 29901
rect 29877 29799 29911 29833
rect 29877 29731 29911 29765
rect 29877 29663 29911 29697
rect 29877 29595 29911 29629
rect 29877 29527 29911 29561
rect 29877 29459 29911 29493
rect 29877 29391 29911 29425
rect 29877 29323 29911 29357
rect 29877 29255 29911 29289
rect 29877 29187 29911 29221
rect 29877 29119 29911 29153
rect 29877 29051 29911 29085
rect 29877 28983 29911 29017
rect 29877 28915 29911 28949
rect 29877 28847 29911 28881
rect 29877 28779 29911 28813
rect 29877 28711 29911 28745
rect 29877 28643 29911 28677
rect 30335 29867 30369 29901
rect 30335 29799 30369 29833
rect 30335 29731 30369 29765
rect 30335 29663 30369 29697
rect 30335 29595 30369 29629
rect 30335 29527 30369 29561
rect 30335 29459 30369 29493
rect 30335 29391 30369 29425
rect 30335 29323 30369 29357
rect 30335 29255 30369 29289
rect 30335 29187 30369 29221
rect 30335 29119 30369 29153
rect 30335 29051 30369 29085
rect 30335 28983 30369 29017
rect 30335 28915 30369 28949
rect 30335 28847 30369 28881
rect 30335 28779 30369 28813
rect 30335 28711 30369 28745
rect 30335 28643 30369 28677
rect 30793 29867 30827 29901
rect 30793 29799 30827 29833
rect 30793 29731 30827 29765
rect 30793 29663 30827 29697
rect 30793 29595 30827 29629
rect 30793 29527 30827 29561
rect 30793 29459 30827 29493
rect 30793 29391 30827 29425
rect 30793 29323 30827 29357
rect 30793 29255 30827 29289
rect 30793 29187 30827 29221
rect 30793 29119 30827 29153
rect 30793 29051 30827 29085
rect 30793 28983 30827 29017
rect 30793 28915 30827 28949
rect 30793 28847 30827 28881
rect 30793 28779 30827 28813
rect 30793 28711 30827 28745
rect 30793 28643 30827 28677
rect 31251 29867 31285 29901
rect 31251 29799 31285 29833
rect 31251 29731 31285 29765
rect 31251 29663 31285 29697
rect 31251 29595 31285 29629
rect 31251 29527 31285 29561
rect 31251 29459 31285 29493
rect 31251 29391 31285 29425
rect 31251 29323 31285 29357
rect 31251 29255 31285 29289
rect 31251 29187 31285 29221
rect 31251 29119 31285 29153
rect 31251 29051 31285 29085
rect 31251 28983 31285 29017
rect 31251 28915 31285 28949
rect 31251 28847 31285 28881
rect 31251 28779 31285 28813
rect 31251 28711 31285 28745
rect 31251 28643 31285 28677
rect 31709 29867 31743 29901
rect 31709 29799 31743 29833
rect 31709 29731 31743 29765
rect 31709 29663 31743 29697
rect 31709 29595 31743 29629
rect 31709 29527 31743 29561
rect 31709 29459 31743 29493
rect 31709 29391 31743 29425
rect 31709 29323 31743 29357
rect 31709 29255 31743 29289
rect 31709 29187 31743 29221
rect 31709 29119 31743 29153
rect 31709 29051 31743 29085
rect 31709 28983 31743 29017
rect 31709 28915 31743 28949
rect 31709 28847 31743 28881
rect 31709 28779 31743 28813
rect 31709 28711 31743 28745
rect 31709 28643 31743 28677
rect 32167 29867 32201 29901
rect 32167 29799 32201 29833
rect 32167 29731 32201 29765
rect 32167 29663 32201 29697
rect 32167 29595 32201 29629
rect 32167 29527 32201 29561
rect 32167 29459 32201 29493
rect 32167 29391 32201 29425
rect 32167 29323 32201 29357
rect 32167 29255 32201 29289
rect 32167 29187 32201 29221
rect 32167 29119 32201 29153
rect 32167 29051 32201 29085
rect 32167 28983 32201 29017
rect 32167 28915 32201 28949
rect 32167 28847 32201 28881
rect 32167 28779 32201 28813
rect 32167 28711 32201 28745
rect 32167 28643 32201 28677
rect 32625 29867 32659 29901
rect 32625 29799 32659 29833
rect 32625 29731 32659 29765
rect 32625 29663 32659 29697
rect 32625 29595 32659 29629
rect 32625 29527 32659 29561
rect 32625 29459 32659 29493
rect 32625 29391 32659 29425
rect 32625 29323 32659 29357
rect 32625 29255 32659 29289
rect 32625 29187 32659 29221
rect 32625 29119 32659 29153
rect 32625 29051 32659 29085
rect 32625 28983 32659 29017
rect 32625 28915 32659 28949
rect 32625 28847 32659 28881
rect 32625 28779 32659 28813
rect 32625 28711 32659 28745
rect 32625 28643 32659 28677
rect 33083 29867 33117 29901
rect 33083 29799 33117 29833
rect 33083 29731 33117 29765
rect 33083 29663 33117 29697
rect 33083 29595 33117 29629
rect 33083 29527 33117 29561
rect 33083 29459 33117 29493
rect 33083 29391 33117 29425
rect 33083 29323 33117 29357
rect 33083 29255 33117 29289
rect 33083 29187 33117 29221
rect 33083 29119 33117 29153
rect 33083 29051 33117 29085
rect 33083 28983 33117 29017
rect 33083 28915 33117 28949
rect 33083 28847 33117 28881
rect 33083 28779 33117 28813
rect 33083 28711 33117 28745
rect 33083 28643 33117 28677
rect 33541 29867 33575 29901
rect 33541 29799 33575 29833
rect 33541 29731 33575 29765
rect 33541 29663 33575 29697
rect 33541 29595 33575 29629
rect 33541 29527 33575 29561
rect 33541 29459 33575 29493
rect 33541 29391 33575 29425
rect 33541 29323 33575 29357
rect 33541 29255 33575 29289
rect 33541 29187 33575 29221
rect 33541 29119 33575 29153
rect 33541 29051 33575 29085
rect 33541 28983 33575 29017
rect 33541 28915 33575 28949
rect 33541 28847 33575 28881
rect 33541 28779 33575 28813
rect 33541 28711 33575 28745
rect 33541 28643 33575 28677
rect 34089 29867 34123 29901
rect 34089 29799 34123 29833
rect 34089 29731 34123 29765
rect 34089 29663 34123 29697
rect 34089 29595 34123 29629
rect 34089 29527 34123 29561
rect 34089 29459 34123 29493
rect 34089 29391 34123 29425
rect 34089 29323 34123 29357
rect 34089 29255 34123 29289
rect 34089 29187 34123 29221
rect 34089 29119 34123 29153
rect 34089 29051 34123 29085
rect 34089 28983 34123 29017
rect 34089 28915 34123 28949
rect 34089 28847 34123 28881
rect 34089 28779 34123 28813
rect 34089 28711 34123 28745
rect 34089 28643 34123 28677
rect 34547 29867 34581 29901
rect 34547 29799 34581 29833
rect 34547 29731 34581 29765
rect 34547 29663 34581 29697
rect 34547 29595 34581 29629
rect 34547 29527 34581 29561
rect 34547 29459 34581 29493
rect 34547 29391 34581 29425
rect 34547 29323 34581 29357
rect 34547 29255 34581 29289
rect 34547 29187 34581 29221
rect 34547 29119 34581 29153
rect 34547 29051 34581 29085
rect 34547 28983 34581 29017
rect 34547 28915 34581 28949
rect 34547 28847 34581 28881
rect 34547 28779 34581 28813
rect 34547 28711 34581 28745
rect 34547 28643 34581 28677
rect 35005 29867 35039 29901
rect 35005 29799 35039 29833
rect 35005 29731 35039 29765
rect 35005 29663 35039 29697
rect 35005 29595 35039 29629
rect 35005 29527 35039 29561
rect 35005 29459 35039 29493
rect 35005 29391 35039 29425
rect 35005 29323 35039 29357
rect 35005 29255 35039 29289
rect 35005 29187 35039 29221
rect 35005 29119 35039 29153
rect 35005 29051 35039 29085
rect 35005 28983 35039 29017
rect 35005 28915 35039 28949
rect 35005 28847 35039 28881
rect 35005 28779 35039 28813
rect 35005 28711 35039 28745
rect 35005 28643 35039 28677
rect 35463 29867 35497 29901
rect 35463 29799 35497 29833
rect 35463 29731 35497 29765
rect 35463 29663 35497 29697
rect 35463 29595 35497 29629
rect 35463 29527 35497 29561
rect 35463 29459 35497 29493
rect 35463 29391 35497 29425
rect 35463 29323 35497 29357
rect 35463 29255 35497 29289
rect 35463 29187 35497 29221
rect 35463 29119 35497 29153
rect 35463 29051 35497 29085
rect 35463 28983 35497 29017
rect 35463 28915 35497 28949
rect 35463 28847 35497 28881
rect 35463 28779 35497 28813
rect 35463 28711 35497 28745
rect 35463 28643 35497 28677
rect 35921 29867 35955 29901
rect 35921 29799 35955 29833
rect 35921 29731 35955 29765
rect 35921 29663 35955 29697
rect 35921 29595 35955 29629
rect 35921 29527 35955 29561
rect 35921 29459 35955 29493
rect 35921 29391 35955 29425
rect 35921 29323 35955 29357
rect 35921 29255 35955 29289
rect 35921 29187 35955 29221
rect 35921 29119 35955 29153
rect 35921 29051 35955 29085
rect 35921 28983 35955 29017
rect 35921 28915 35955 28949
rect 35921 28847 35955 28881
rect 35921 28779 35955 28813
rect 35921 28711 35955 28745
rect 35921 28643 35955 28677
rect 36379 29867 36413 29901
rect 36379 29799 36413 29833
rect 36379 29731 36413 29765
rect 36379 29663 36413 29697
rect 36379 29595 36413 29629
rect 36379 29527 36413 29561
rect 36379 29459 36413 29493
rect 36379 29391 36413 29425
rect 36379 29323 36413 29357
rect 36379 29255 36413 29289
rect 36379 29187 36413 29221
rect 36379 29119 36413 29153
rect 36379 29051 36413 29085
rect 36379 28983 36413 29017
rect 36379 28915 36413 28949
rect 36379 28847 36413 28881
rect 36379 28779 36413 28813
rect 36379 28711 36413 28745
rect 36379 28643 36413 28677
rect 36837 29867 36871 29901
rect 36837 29799 36871 29833
rect 36837 29731 36871 29765
rect 36837 29663 36871 29697
rect 36837 29595 36871 29629
rect 36837 29527 36871 29561
rect 36837 29459 36871 29493
rect 36837 29391 36871 29425
rect 36837 29323 36871 29357
rect 36837 29255 36871 29289
rect 36837 29187 36871 29221
rect 36837 29119 36871 29153
rect 36837 29051 36871 29085
rect 36837 28983 36871 29017
rect 36837 28915 36871 28949
rect 36837 28847 36871 28881
rect 36837 28779 36871 28813
rect 36837 28711 36871 28745
rect 36837 28643 36871 28677
rect 9589 26107 9623 26141
rect 9589 26039 9623 26073
rect 9589 25971 9623 26005
rect 9589 25903 9623 25937
rect 9589 25835 9623 25869
rect 9589 25767 9623 25801
rect 9589 25699 9623 25733
rect 9589 25631 9623 25665
rect 9589 25563 9623 25597
rect 9589 25495 9623 25529
rect 9589 25427 9623 25461
rect 9589 25359 9623 25393
rect 9589 25291 9623 25325
rect 9589 25223 9623 25257
rect 9589 25155 9623 25189
rect 9589 25087 9623 25121
rect 9589 25019 9623 25053
rect 9589 24951 9623 24985
rect 9589 24883 9623 24917
rect 10047 26107 10081 26141
rect 10047 26039 10081 26073
rect 10047 25971 10081 26005
rect 10047 25903 10081 25937
rect 10047 25835 10081 25869
rect 10047 25767 10081 25801
rect 10047 25699 10081 25733
rect 10047 25631 10081 25665
rect 10047 25563 10081 25597
rect 10047 25495 10081 25529
rect 10047 25427 10081 25461
rect 10047 25359 10081 25393
rect 10047 25291 10081 25325
rect 10047 25223 10081 25257
rect 10047 25155 10081 25189
rect 10047 25087 10081 25121
rect 10047 25019 10081 25053
rect 10047 24951 10081 24985
rect 10047 24883 10081 24917
rect 10505 26107 10539 26141
rect 10505 26039 10539 26073
rect 10505 25971 10539 26005
rect 10505 25903 10539 25937
rect 10505 25835 10539 25869
rect 10505 25767 10539 25801
rect 10505 25699 10539 25733
rect 10505 25631 10539 25665
rect 10505 25563 10539 25597
rect 10505 25495 10539 25529
rect 10505 25427 10539 25461
rect 10505 25359 10539 25393
rect 10505 25291 10539 25325
rect 10505 25223 10539 25257
rect 10505 25155 10539 25189
rect 10505 25087 10539 25121
rect 10505 25019 10539 25053
rect 10505 24951 10539 24985
rect 10505 24883 10539 24917
rect 10963 26107 10997 26141
rect 10963 26039 10997 26073
rect 10963 25971 10997 26005
rect 10963 25903 10997 25937
rect 10963 25835 10997 25869
rect 10963 25767 10997 25801
rect 10963 25699 10997 25733
rect 10963 25631 10997 25665
rect 10963 25563 10997 25597
rect 10963 25495 10997 25529
rect 10963 25427 10997 25461
rect 10963 25359 10997 25393
rect 10963 25291 10997 25325
rect 10963 25223 10997 25257
rect 10963 25155 10997 25189
rect 10963 25087 10997 25121
rect 10963 25019 10997 25053
rect 10963 24951 10997 24985
rect 10963 24883 10997 24917
rect 11421 26107 11455 26141
rect 11421 26039 11455 26073
rect 11421 25971 11455 26005
rect 11421 25903 11455 25937
rect 11421 25835 11455 25869
rect 11421 25767 11455 25801
rect 11421 25699 11455 25733
rect 11421 25631 11455 25665
rect 11421 25563 11455 25597
rect 11421 25495 11455 25529
rect 11421 25427 11455 25461
rect 11421 25359 11455 25393
rect 11421 25291 11455 25325
rect 11421 25223 11455 25257
rect 11421 25155 11455 25189
rect 11421 25087 11455 25121
rect 11421 25019 11455 25053
rect 11421 24951 11455 24985
rect 11421 24883 11455 24917
rect 11879 26107 11913 26141
rect 11879 26039 11913 26073
rect 11879 25971 11913 26005
rect 11879 25903 11913 25937
rect 11879 25835 11913 25869
rect 11879 25767 11913 25801
rect 11879 25699 11913 25733
rect 11879 25631 11913 25665
rect 11879 25563 11913 25597
rect 11879 25495 11913 25529
rect 11879 25427 11913 25461
rect 11879 25359 11913 25393
rect 11879 25291 11913 25325
rect 11879 25223 11913 25257
rect 11879 25155 11913 25189
rect 11879 25087 11913 25121
rect 11879 25019 11913 25053
rect 11879 24951 11913 24985
rect 11879 24883 11913 24917
rect 12337 26107 12371 26141
rect 12337 26039 12371 26073
rect 12337 25971 12371 26005
rect 12337 25903 12371 25937
rect 12337 25835 12371 25869
rect 12337 25767 12371 25801
rect 12337 25699 12371 25733
rect 12337 25631 12371 25665
rect 12337 25563 12371 25597
rect 12337 25495 12371 25529
rect 12337 25427 12371 25461
rect 12337 25359 12371 25393
rect 12337 25291 12371 25325
rect 12337 25223 12371 25257
rect 12337 25155 12371 25189
rect 12337 25087 12371 25121
rect 12337 25019 12371 25053
rect 12337 24951 12371 24985
rect 12337 24883 12371 24917
rect 12795 26107 12829 26141
rect 12795 26039 12829 26073
rect 12795 25971 12829 26005
rect 12795 25903 12829 25937
rect 12795 25835 12829 25869
rect 12795 25767 12829 25801
rect 12795 25699 12829 25733
rect 12795 25631 12829 25665
rect 12795 25563 12829 25597
rect 12795 25495 12829 25529
rect 12795 25427 12829 25461
rect 12795 25359 12829 25393
rect 12795 25291 12829 25325
rect 12795 25223 12829 25257
rect 12795 25155 12829 25189
rect 12795 25087 12829 25121
rect 12795 25019 12829 25053
rect 12795 24951 12829 24985
rect 12795 24883 12829 24917
rect 13253 26107 13287 26141
rect 13253 26039 13287 26073
rect 13253 25971 13287 26005
rect 13253 25903 13287 25937
rect 13253 25835 13287 25869
rect 13253 25767 13287 25801
rect 13253 25699 13287 25733
rect 13253 25631 13287 25665
rect 13253 25563 13287 25597
rect 13253 25495 13287 25529
rect 13253 25427 13287 25461
rect 13253 25359 13287 25393
rect 13253 25291 13287 25325
rect 13253 25223 13287 25257
rect 13253 25155 13287 25189
rect 13253 25087 13287 25121
rect 13253 25019 13287 25053
rect 13253 24951 13287 24985
rect 13253 24883 13287 24917
rect 13711 26107 13745 26141
rect 13711 26039 13745 26073
rect 13711 25971 13745 26005
rect 13711 25903 13745 25937
rect 13711 25835 13745 25869
rect 13711 25767 13745 25801
rect 13711 25699 13745 25733
rect 13711 25631 13745 25665
rect 13711 25563 13745 25597
rect 13711 25495 13745 25529
rect 13711 25427 13745 25461
rect 13711 25359 13745 25393
rect 13711 25291 13745 25325
rect 13711 25223 13745 25257
rect 13711 25155 13745 25189
rect 13711 25087 13745 25121
rect 13711 25019 13745 25053
rect 13711 24951 13745 24985
rect 13711 24883 13745 24917
rect 14169 26107 14203 26141
rect 14169 26039 14203 26073
rect 14169 25971 14203 26005
rect 14169 25903 14203 25937
rect 14169 25835 14203 25869
rect 14169 25767 14203 25801
rect 14169 25699 14203 25733
rect 14169 25631 14203 25665
rect 14169 25563 14203 25597
rect 14169 25495 14203 25529
rect 14169 25427 14203 25461
rect 14169 25359 14203 25393
rect 14169 25291 14203 25325
rect 14169 25223 14203 25257
rect 14169 25155 14203 25189
rect 14169 25087 14203 25121
rect 14169 25019 14203 25053
rect 14169 24951 14203 24985
rect 14169 24883 14203 24917
rect 14627 26107 14661 26141
rect 14627 26039 14661 26073
rect 14627 25971 14661 26005
rect 14627 25903 14661 25937
rect 14627 25835 14661 25869
rect 14627 25767 14661 25801
rect 14627 25699 14661 25733
rect 14627 25631 14661 25665
rect 14627 25563 14661 25597
rect 14627 25495 14661 25529
rect 14627 25427 14661 25461
rect 14627 25359 14661 25393
rect 14627 25291 14661 25325
rect 14627 25223 14661 25257
rect 14627 25155 14661 25189
rect 14627 25087 14661 25121
rect 14627 25019 14661 25053
rect 14627 24951 14661 24985
rect 14627 24883 14661 24917
rect 15085 26107 15119 26141
rect 15085 26039 15119 26073
rect 15085 25971 15119 26005
rect 15085 25903 15119 25937
rect 15085 25835 15119 25869
rect 15085 25767 15119 25801
rect 15085 25699 15119 25733
rect 15085 25631 15119 25665
rect 15085 25563 15119 25597
rect 15085 25495 15119 25529
rect 15085 25427 15119 25461
rect 15085 25359 15119 25393
rect 15085 25291 15119 25325
rect 15085 25223 15119 25257
rect 15085 25155 15119 25189
rect 15085 25087 15119 25121
rect 15085 25019 15119 25053
rect 15085 24951 15119 24985
rect 15085 24883 15119 24917
rect 28644 25706 28678 25740
rect 28734 25706 28768 25740
rect 28824 25706 28858 25740
rect 28914 25706 28948 25740
rect 29004 25706 29038 25740
rect 29094 25706 29128 25740
rect 29184 25706 29218 25740
rect 28644 25616 28678 25650
rect 28734 25616 28768 25650
rect 28824 25616 28858 25650
rect 28914 25616 28948 25650
rect 29004 25616 29038 25650
rect 29094 25616 29128 25650
rect 29184 25616 29218 25650
rect 28644 25526 28678 25560
rect 28734 25526 28768 25560
rect 28824 25526 28858 25560
rect 28914 25526 28948 25560
rect 29004 25526 29038 25560
rect 29094 25526 29128 25560
rect 29184 25526 29218 25560
rect 28644 25436 28678 25470
rect 28734 25436 28768 25470
rect 28824 25436 28858 25470
rect 28914 25436 28948 25470
rect 29004 25436 29038 25470
rect 29094 25436 29128 25470
rect 29184 25436 29218 25470
rect 28644 25346 28678 25380
rect 28734 25346 28768 25380
rect 28824 25346 28858 25380
rect 28914 25346 28948 25380
rect 29004 25346 29038 25380
rect 29094 25346 29128 25380
rect 29184 25346 29218 25380
rect 28644 25256 28678 25290
rect 28734 25256 28768 25290
rect 28824 25256 28858 25290
rect 28914 25256 28948 25290
rect 29004 25256 29038 25290
rect 29094 25256 29128 25290
rect 29184 25256 29218 25290
rect 28644 25166 28678 25200
rect 28734 25166 28768 25200
rect 28824 25166 28858 25200
rect 28914 25166 28948 25200
rect 29004 25166 29038 25200
rect 29094 25166 29128 25200
rect 29184 25166 29218 25200
rect 29984 25706 30018 25740
rect 30074 25706 30108 25740
rect 30164 25706 30198 25740
rect 30254 25706 30288 25740
rect 30344 25706 30378 25740
rect 30434 25706 30468 25740
rect 30524 25706 30558 25740
rect 29984 25616 30018 25650
rect 30074 25616 30108 25650
rect 30164 25616 30198 25650
rect 30254 25616 30288 25650
rect 30344 25616 30378 25650
rect 30434 25616 30468 25650
rect 30524 25616 30558 25650
rect 29984 25526 30018 25560
rect 30074 25526 30108 25560
rect 30164 25526 30198 25560
rect 30254 25526 30288 25560
rect 30344 25526 30378 25560
rect 30434 25526 30468 25560
rect 30524 25526 30558 25560
rect 29984 25436 30018 25470
rect 30074 25436 30108 25470
rect 30164 25436 30198 25470
rect 30254 25436 30288 25470
rect 30344 25436 30378 25470
rect 30434 25436 30468 25470
rect 30524 25436 30558 25470
rect 29984 25346 30018 25380
rect 30074 25346 30108 25380
rect 30164 25346 30198 25380
rect 30254 25346 30288 25380
rect 30344 25346 30378 25380
rect 30434 25346 30468 25380
rect 30524 25346 30558 25380
rect 29984 25256 30018 25290
rect 30074 25256 30108 25290
rect 30164 25256 30198 25290
rect 30254 25256 30288 25290
rect 30344 25256 30378 25290
rect 30434 25256 30468 25290
rect 30524 25256 30558 25290
rect 29984 25166 30018 25200
rect 30074 25166 30108 25200
rect 30164 25166 30198 25200
rect 30254 25166 30288 25200
rect 30344 25166 30378 25200
rect 30434 25166 30468 25200
rect 30524 25166 30558 25200
rect 31324 25706 31358 25740
rect 31414 25706 31448 25740
rect 31504 25706 31538 25740
rect 31594 25706 31628 25740
rect 31684 25706 31718 25740
rect 31774 25706 31808 25740
rect 31864 25706 31898 25740
rect 31324 25616 31358 25650
rect 31414 25616 31448 25650
rect 31504 25616 31538 25650
rect 31594 25616 31628 25650
rect 31684 25616 31718 25650
rect 31774 25616 31808 25650
rect 31864 25616 31898 25650
rect 31324 25526 31358 25560
rect 31414 25526 31448 25560
rect 31504 25526 31538 25560
rect 31594 25526 31628 25560
rect 31684 25526 31718 25560
rect 31774 25526 31808 25560
rect 31864 25526 31898 25560
rect 31324 25436 31358 25470
rect 31414 25436 31448 25470
rect 31504 25436 31538 25470
rect 31594 25436 31628 25470
rect 31684 25436 31718 25470
rect 31774 25436 31808 25470
rect 31864 25436 31898 25470
rect 31324 25346 31358 25380
rect 31414 25346 31448 25380
rect 31504 25346 31538 25380
rect 31594 25346 31628 25380
rect 31684 25346 31718 25380
rect 31774 25346 31808 25380
rect 31864 25346 31898 25380
rect 31324 25256 31358 25290
rect 31414 25256 31448 25290
rect 31504 25256 31538 25290
rect 31594 25256 31628 25290
rect 31684 25256 31718 25290
rect 31774 25256 31808 25290
rect 31864 25256 31898 25290
rect 31324 25166 31358 25200
rect 31414 25166 31448 25200
rect 31504 25166 31538 25200
rect 31594 25166 31628 25200
rect 31684 25166 31718 25200
rect 31774 25166 31808 25200
rect 31864 25166 31898 25200
rect 32664 25706 32698 25740
rect 32754 25706 32788 25740
rect 32844 25706 32878 25740
rect 32934 25706 32968 25740
rect 33024 25706 33058 25740
rect 33114 25706 33148 25740
rect 33204 25706 33238 25740
rect 32664 25616 32698 25650
rect 32754 25616 32788 25650
rect 32844 25616 32878 25650
rect 32934 25616 32968 25650
rect 33024 25616 33058 25650
rect 33114 25616 33148 25650
rect 33204 25616 33238 25650
rect 32664 25526 32698 25560
rect 32754 25526 32788 25560
rect 32844 25526 32878 25560
rect 32934 25526 32968 25560
rect 33024 25526 33058 25560
rect 33114 25526 33148 25560
rect 33204 25526 33238 25560
rect 32664 25436 32698 25470
rect 32754 25436 32788 25470
rect 32844 25436 32878 25470
rect 32934 25436 32968 25470
rect 33024 25436 33058 25470
rect 33114 25436 33148 25470
rect 33204 25436 33238 25470
rect 32664 25346 32698 25380
rect 32754 25346 32788 25380
rect 32844 25346 32878 25380
rect 32934 25346 32968 25380
rect 33024 25346 33058 25380
rect 33114 25346 33148 25380
rect 33204 25346 33238 25380
rect 32664 25256 32698 25290
rect 32754 25256 32788 25290
rect 32844 25256 32878 25290
rect 32934 25256 32968 25290
rect 33024 25256 33058 25290
rect 33114 25256 33148 25290
rect 33204 25256 33238 25290
rect 32664 25166 32698 25200
rect 32754 25166 32788 25200
rect 32844 25166 32878 25200
rect 32934 25166 32968 25200
rect 33024 25166 33058 25200
rect 33114 25166 33148 25200
rect 33204 25166 33238 25200
rect 34004 25706 34038 25740
rect 34094 25706 34128 25740
rect 34184 25706 34218 25740
rect 34274 25706 34308 25740
rect 34364 25706 34398 25740
rect 34454 25706 34488 25740
rect 34544 25706 34578 25740
rect 34004 25616 34038 25650
rect 34094 25616 34128 25650
rect 34184 25616 34218 25650
rect 34274 25616 34308 25650
rect 34364 25616 34398 25650
rect 34454 25616 34488 25650
rect 34544 25616 34578 25650
rect 34004 25526 34038 25560
rect 34094 25526 34128 25560
rect 34184 25526 34218 25560
rect 34274 25526 34308 25560
rect 34364 25526 34398 25560
rect 34454 25526 34488 25560
rect 34544 25526 34578 25560
rect 34004 25436 34038 25470
rect 34094 25436 34128 25470
rect 34184 25436 34218 25470
rect 34274 25436 34308 25470
rect 34364 25436 34398 25470
rect 34454 25436 34488 25470
rect 34544 25436 34578 25470
rect 34004 25346 34038 25380
rect 34094 25346 34128 25380
rect 34184 25346 34218 25380
rect 34274 25346 34308 25380
rect 34364 25346 34398 25380
rect 34454 25346 34488 25380
rect 34544 25346 34578 25380
rect 34004 25256 34038 25290
rect 34094 25256 34128 25290
rect 34184 25256 34218 25290
rect 34274 25256 34308 25290
rect 34364 25256 34398 25290
rect 34454 25256 34488 25290
rect 34544 25256 34578 25290
rect 34004 25166 34038 25200
rect 34094 25166 34128 25200
rect 34184 25166 34218 25200
rect 34274 25166 34308 25200
rect 34364 25166 34398 25200
rect 34454 25166 34488 25200
rect 34544 25166 34578 25200
rect 35344 25706 35378 25740
rect 35434 25706 35468 25740
rect 35524 25706 35558 25740
rect 35614 25706 35648 25740
rect 35704 25706 35738 25740
rect 35794 25706 35828 25740
rect 35884 25706 35918 25740
rect 35344 25616 35378 25650
rect 35434 25616 35468 25650
rect 35524 25616 35558 25650
rect 35614 25616 35648 25650
rect 35704 25616 35738 25650
rect 35794 25616 35828 25650
rect 35884 25616 35918 25650
rect 35344 25526 35378 25560
rect 35434 25526 35468 25560
rect 35524 25526 35558 25560
rect 35614 25526 35648 25560
rect 35704 25526 35738 25560
rect 35794 25526 35828 25560
rect 35884 25526 35918 25560
rect 35344 25436 35378 25470
rect 35434 25436 35468 25470
rect 35524 25436 35558 25470
rect 35614 25436 35648 25470
rect 35704 25436 35738 25470
rect 35794 25436 35828 25470
rect 35884 25436 35918 25470
rect 35344 25346 35378 25380
rect 35434 25346 35468 25380
rect 35524 25346 35558 25380
rect 35614 25346 35648 25380
rect 35704 25346 35738 25380
rect 35794 25346 35828 25380
rect 35884 25346 35918 25380
rect 35344 25256 35378 25290
rect 35434 25256 35468 25290
rect 35524 25256 35558 25290
rect 35614 25256 35648 25290
rect 35704 25256 35738 25290
rect 35794 25256 35828 25290
rect 35884 25256 35918 25290
rect 35344 25166 35378 25200
rect 35434 25166 35468 25200
rect 35524 25166 35558 25200
rect 35614 25166 35648 25200
rect 35704 25166 35738 25200
rect 35794 25166 35828 25200
rect 35884 25166 35918 25200
rect 36684 25706 36718 25740
rect 36774 25706 36808 25740
rect 36864 25706 36898 25740
rect 36954 25706 36988 25740
rect 37044 25706 37078 25740
rect 37134 25706 37168 25740
rect 37224 25706 37258 25740
rect 36684 25616 36718 25650
rect 36774 25616 36808 25650
rect 36864 25616 36898 25650
rect 36954 25616 36988 25650
rect 37044 25616 37078 25650
rect 37134 25616 37168 25650
rect 37224 25616 37258 25650
rect 36684 25526 36718 25560
rect 36774 25526 36808 25560
rect 36864 25526 36898 25560
rect 36954 25526 36988 25560
rect 37044 25526 37078 25560
rect 37134 25526 37168 25560
rect 37224 25526 37258 25560
rect 36684 25436 36718 25470
rect 36774 25436 36808 25470
rect 36864 25436 36898 25470
rect 36954 25436 36988 25470
rect 37044 25436 37078 25470
rect 37134 25436 37168 25470
rect 37224 25436 37258 25470
rect 36684 25346 36718 25380
rect 36774 25346 36808 25380
rect 36864 25346 36898 25380
rect 36954 25346 36988 25380
rect 37044 25346 37078 25380
rect 37134 25346 37168 25380
rect 37224 25346 37258 25380
rect 36684 25256 36718 25290
rect 36774 25256 36808 25290
rect 36864 25256 36898 25290
rect 36954 25256 36988 25290
rect 37044 25256 37078 25290
rect 37134 25256 37168 25290
rect 37224 25256 37258 25290
rect 36684 25166 36718 25200
rect 36774 25166 36808 25200
rect 36864 25166 36898 25200
rect 36954 25166 36988 25200
rect 37044 25166 37078 25200
rect 37134 25166 37168 25200
rect 37224 25166 37258 25200
rect 38024 25706 38058 25740
rect 38114 25706 38148 25740
rect 38204 25706 38238 25740
rect 38294 25706 38328 25740
rect 38384 25706 38418 25740
rect 38474 25706 38508 25740
rect 38564 25706 38598 25740
rect 38024 25616 38058 25650
rect 38114 25616 38148 25650
rect 38204 25616 38238 25650
rect 38294 25616 38328 25650
rect 38384 25616 38418 25650
rect 38474 25616 38508 25650
rect 38564 25616 38598 25650
rect 38024 25526 38058 25560
rect 38114 25526 38148 25560
rect 38204 25526 38238 25560
rect 38294 25526 38328 25560
rect 38384 25526 38418 25560
rect 38474 25526 38508 25560
rect 38564 25526 38598 25560
rect 38024 25436 38058 25470
rect 38114 25436 38148 25470
rect 38204 25436 38238 25470
rect 38294 25436 38328 25470
rect 38384 25436 38418 25470
rect 38474 25436 38508 25470
rect 38564 25436 38598 25470
rect 38024 25346 38058 25380
rect 38114 25346 38148 25380
rect 38204 25346 38238 25380
rect 38294 25346 38328 25380
rect 38384 25346 38418 25380
rect 38474 25346 38508 25380
rect 38564 25346 38598 25380
rect 38024 25256 38058 25290
rect 38114 25256 38148 25290
rect 38204 25256 38238 25290
rect 38294 25256 38328 25290
rect 38384 25256 38418 25290
rect 38474 25256 38508 25290
rect 38564 25256 38598 25290
rect 38024 25166 38058 25200
rect 38114 25166 38148 25200
rect 38204 25166 38238 25200
rect 38294 25166 38328 25200
rect 38384 25166 38418 25200
rect 38474 25166 38508 25200
rect 38564 25166 38598 25200
rect 7727 22347 7761 22381
rect 7727 22279 7761 22313
rect 7727 22211 7761 22245
rect 7727 22143 7761 22177
rect 7727 22075 7761 22109
rect 7727 22007 7761 22041
rect 7727 21939 7761 21973
rect 7727 21871 7761 21905
rect 7727 21803 7761 21837
rect 7727 21735 7761 21769
rect 7727 21667 7761 21701
rect 7727 21599 7761 21633
rect 7727 21531 7761 21565
rect 7727 21463 7761 21497
rect 7727 21395 7761 21429
rect 7727 21327 7761 21361
rect 7727 21259 7761 21293
rect 7727 21191 7761 21225
rect 7727 21123 7761 21157
rect 8185 22347 8219 22381
rect 8185 22279 8219 22313
rect 8185 22211 8219 22245
rect 8185 22143 8219 22177
rect 8185 22075 8219 22109
rect 8185 22007 8219 22041
rect 8185 21939 8219 21973
rect 8185 21871 8219 21905
rect 8185 21803 8219 21837
rect 8185 21735 8219 21769
rect 8185 21667 8219 21701
rect 8185 21599 8219 21633
rect 8185 21531 8219 21565
rect 8185 21463 8219 21497
rect 8185 21395 8219 21429
rect 8185 21327 8219 21361
rect 8185 21259 8219 21293
rect 8185 21191 8219 21225
rect 8185 21123 8219 21157
rect 8643 22347 8677 22381
rect 8643 22279 8677 22313
rect 8643 22211 8677 22245
rect 8643 22143 8677 22177
rect 8643 22075 8677 22109
rect 8643 22007 8677 22041
rect 8643 21939 8677 21973
rect 8643 21871 8677 21905
rect 8643 21803 8677 21837
rect 8643 21735 8677 21769
rect 8643 21667 8677 21701
rect 8643 21599 8677 21633
rect 8643 21531 8677 21565
rect 8643 21463 8677 21497
rect 8643 21395 8677 21429
rect 8643 21327 8677 21361
rect 8643 21259 8677 21293
rect 8643 21191 8677 21225
rect 8643 21123 8677 21157
rect 9101 22347 9135 22381
rect 9101 22279 9135 22313
rect 9101 22211 9135 22245
rect 9101 22143 9135 22177
rect 9101 22075 9135 22109
rect 9101 22007 9135 22041
rect 9101 21939 9135 21973
rect 9101 21871 9135 21905
rect 9101 21803 9135 21837
rect 9101 21735 9135 21769
rect 9101 21667 9135 21701
rect 9101 21599 9135 21633
rect 9101 21531 9135 21565
rect 9101 21463 9135 21497
rect 9101 21395 9135 21429
rect 9101 21327 9135 21361
rect 9101 21259 9135 21293
rect 9101 21191 9135 21225
rect 9101 21123 9135 21157
rect 9559 22347 9593 22381
rect 9559 22279 9593 22313
rect 9559 22211 9593 22245
rect 9559 22143 9593 22177
rect 9559 22075 9593 22109
rect 9559 22007 9593 22041
rect 9559 21939 9593 21973
rect 9559 21871 9593 21905
rect 9559 21803 9593 21837
rect 9559 21735 9593 21769
rect 9559 21667 9593 21701
rect 9559 21599 9593 21633
rect 9559 21531 9593 21565
rect 9559 21463 9593 21497
rect 9559 21395 9593 21429
rect 9559 21327 9593 21361
rect 9559 21259 9593 21293
rect 9559 21191 9593 21225
rect 9559 21123 9593 21157
rect 10017 22347 10051 22381
rect 10017 22279 10051 22313
rect 10017 22211 10051 22245
rect 10017 22143 10051 22177
rect 10017 22075 10051 22109
rect 10017 22007 10051 22041
rect 10017 21939 10051 21973
rect 10017 21871 10051 21905
rect 10017 21803 10051 21837
rect 10017 21735 10051 21769
rect 10017 21667 10051 21701
rect 10017 21599 10051 21633
rect 10017 21531 10051 21565
rect 10017 21463 10051 21497
rect 10017 21395 10051 21429
rect 10017 21327 10051 21361
rect 10017 21259 10051 21293
rect 10017 21191 10051 21225
rect 10017 21123 10051 21157
rect 10475 22347 10509 22381
rect 10475 22279 10509 22313
rect 10475 22211 10509 22245
rect 10475 22143 10509 22177
rect 10475 22075 10509 22109
rect 10475 22007 10509 22041
rect 10475 21939 10509 21973
rect 10475 21871 10509 21905
rect 10475 21803 10509 21837
rect 10475 21735 10509 21769
rect 10475 21667 10509 21701
rect 10475 21599 10509 21633
rect 10475 21531 10509 21565
rect 10475 21463 10509 21497
rect 10475 21395 10509 21429
rect 10475 21327 10509 21361
rect 10475 21259 10509 21293
rect 10475 21191 10509 21225
rect 10475 21123 10509 21157
rect 10933 22347 10967 22381
rect 10933 22279 10967 22313
rect 10933 22211 10967 22245
rect 10933 22143 10967 22177
rect 10933 22075 10967 22109
rect 10933 22007 10967 22041
rect 10933 21939 10967 21973
rect 10933 21871 10967 21905
rect 10933 21803 10967 21837
rect 10933 21735 10967 21769
rect 10933 21667 10967 21701
rect 10933 21599 10967 21633
rect 10933 21531 10967 21565
rect 10933 21463 10967 21497
rect 10933 21395 10967 21429
rect 10933 21327 10967 21361
rect 10933 21259 10967 21293
rect 10933 21191 10967 21225
rect 10933 21123 10967 21157
rect 11391 22347 11425 22381
rect 11391 22279 11425 22313
rect 11391 22211 11425 22245
rect 11391 22143 11425 22177
rect 11391 22075 11425 22109
rect 11391 22007 11425 22041
rect 11391 21939 11425 21973
rect 11391 21871 11425 21905
rect 11391 21803 11425 21837
rect 11391 21735 11425 21769
rect 11391 21667 11425 21701
rect 11391 21599 11425 21633
rect 11391 21531 11425 21565
rect 11391 21463 11425 21497
rect 11391 21395 11425 21429
rect 11391 21327 11425 21361
rect 11391 21259 11425 21293
rect 11391 21191 11425 21225
rect 11391 21123 11425 21157
rect 11849 22347 11883 22381
rect 11849 22279 11883 22313
rect 11849 22211 11883 22245
rect 11849 22143 11883 22177
rect 11849 22075 11883 22109
rect 11849 22007 11883 22041
rect 11849 21939 11883 21973
rect 11849 21871 11883 21905
rect 11849 21803 11883 21837
rect 11849 21735 11883 21769
rect 11849 21667 11883 21701
rect 11849 21599 11883 21633
rect 11849 21531 11883 21565
rect 11849 21463 11883 21497
rect 11849 21395 11883 21429
rect 11849 21327 11883 21361
rect 11849 21259 11883 21293
rect 11849 21191 11883 21225
rect 11849 21123 11883 21157
rect 12307 22347 12341 22381
rect 12307 22279 12341 22313
rect 12307 22211 12341 22245
rect 12307 22143 12341 22177
rect 12307 22075 12341 22109
rect 12307 22007 12341 22041
rect 12307 21939 12341 21973
rect 12307 21871 12341 21905
rect 12307 21803 12341 21837
rect 12307 21735 12341 21769
rect 12307 21667 12341 21701
rect 12307 21599 12341 21633
rect 12307 21531 12341 21565
rect 12307 21463 12341 21497
rect 12307 21395 12341 21429
rect 12307 21327 12341 21361
rect 12307 21259 12341 21293
rect 12307 21191 12341 21225
rect 12307 21123 12341 21157
rect 12765 22347 12799 22381
rect 12765 22279 12799 22313
rect 12765 22211 12799 22245
rect 12765 22143 12799 22177
rect 12765 22075 12799 22109
rect 12765 22007 12799 22041
rect 12765 21939 12799 21973
rect 12765 21871 12799 21905
rect 12765 21803 12799 21837
rect 12765 21735 12799 21769
rect 12765 21667 12799 21701
rect 12765 21599 12799 21633
rect 12765 21531 12799 21565
rect 12765 21463 12799 21497
rect 12765 21395 12799 21429
rect 12765 21327 12799 21361
rect 12765 21259 12799 21293
rect 12765 21191 12799 21225
rect 12765 21123 12799 21157
rect 13223 22347 13257 22381
rect 13223 22279 13257 22313
rect 13223 22211 13257 22245
rect 13223 22143 13257 22177
rect 13223 22075 13257 22109
rect 13223 22007 13257 22041
rect 13223 21939 13257 21973
rect 13223 21871 13257 21905
rect 13223 21803 13257 21837
rect 13223 21735 13257 21769
rect 13223 21667 13257 21701
rect 13223 21599 13257 21633
rect 13223 21531 13257 21565
rect 13223 21463 13257 21497
rect 13223 21395 13257 21429
rect 13223 21327 13257 21361
rect 13223 21259 13257 21293
rect 13223 21191 13257 21225
rect 13223 21123 13257 21157
rect 21392 21946 21426 21980
rect 21482 21946 21516 21980
rect 21572 21946 21606 21980
rect 21662 21946 21696 21980
rect 21752 21946 21786 21980
rect 21842 21946 21876 21980
rect 21932 21946 21966 21980
rect 21392 21856 21426 21890
rect 21482 21856 21516 21890
rect 21572 21856 21606 21890
rect 21662 21856 21696 21890
rect 21752 21856 21786 21890
rect 21842 21856 21876 21890
rect 21932 21856 21966 21890
rect 21392 21766 21426 21800
rect 21482 21766 21516 21800
rect 21572 21766 21606 21800
rect 21662 21766 21696 21800
rect 21752 21766 21786 21800
rect 21842 21766 21876 21800
rect 21932 21766 21966 21800
rect 21392 21676 21426 21710
rect 21482 21676 21516 21710
rect 21572 21676 21606 21710
rect 21662 21676 21696 21710
rect 21752 21676 21786 21710
rect 21842 21676 21876 21710
rect 21932 21676 21966 21710
rect 21392 21586 21426 21620
rect 21482 21586 21516 21620
rect 21572 21586 21606 21620
rect 21662 21586 21696 21620
rect 21752 21586 21786 21620
rect 21842 21586 21876 21620
rect 21932 21586 21966 21620
rect 21392 21496 21426 21530
rect 21482 21496 21516 21530
rect 21572 21496 21606 21530
rect 21662 21496 21696 21530
rect 21752 21496 21786 21530
rect 21842 21496 21876 21530
rect 21932 21496 21966 21530
rect 21392 21406 21426 21440
rect 21482 21406 21516 21440
rect 21572 21406 21606 21440
rect 21662 21406 21696 21440
rect 21752 21406 21786 21440
rect 21842 21406 21876 21440
rect 21932 21406 21966 21440
rect 28644 21946 28678 21980
rect 28734 21946 28768 21980
rect 28824 21946 28858 21980
rect 28914 21946 28948 21980
rect 29004 21946 29038 21980
rect 29094 21946 29128 21980
rect 29184 21946 29218 21980
rect 28644 21856 28678 21890
rect 28734 21856 28768 21890
rect 28824 21856 28858 21890
rect 28914 21856 28948 21890
rect 29004 21856 29038 21890
rect 29094 21856 29128 21890
rect 29184 21856 29218 21890
rect 28644 21766 28678 21800
rect 28734 21766 28768 21800
rect 28824 21766 28858 21800
rect 28914 21766 28948 21800
rect 29004 21766 29038 21800
rect 29094 21766 29128 21800
rect 29184 21766 29218 21800
rect 28644 21676 28678 21710
rect 28734 21676 28768 21710
rect 28824 21676 28858 21710
rect 28914 21676 28948 21710
rect 29004 21676 29038 21710
rect 29094 21676 29128 21710
rect 29184 21676 29218 21710
rect 28644 21586 28678 21620
rect 28734 21586 28768 21620
rect 28824 21586 28858 21620
rect 28914 21586 28948 21620
rect 29004 21586 29038 21620
rect 29094 21586 29128 21620
rect 29184 21586 29218 21620
rect 28644 21496 28678 21530
rect 28734 21496 28768 21530
rect 28824 21496 28858 21530
rect 28914 21496 28948 21530
rect 29004 21496 29038 21530
rect 29094 21496 29128 21530
rect 29184 21496 29218 21530
rect 28644 21406 28678 21440
rect 28734 21406 28768 21440
rect 28824 21406 28858 21440
rect 28914 21406 28948 21440
rect 29004 21406 29038 21440
rect 29094 21406 29128 21440
rect 29184 21406 29218 21440
rect 29984 21946 30018 21980
rect 30074 21946 30108 21980
rect 30164 21946 30198 21980
rect 30254 21946 30288 21980
rect 30344 21946 30378 21980
rect 30434 21946 30468 21980
rect 30524 21946 30558 21980
rect 29984 21856 30018 21890
rect 30074 21856 30108 21890
rect 30164 21856 30198 21890
rect 30254 21856 30288 21890
rect 30344 21856 30378 21890
rect 30434 21856 30468 21890
rect 30524 21856 30558 21890
rect 29984 21766 30018 21800
rect 30074 21766 30108 21800
rect 30164 21766 30198 21800
rect 30254 21766 30288 21800
rect 30344 21766 30378 21800
rect 30434 21766 30468 21800
rect 30524 21766 30558 21800
rect 29984 21676 30018 21710
rect 30074 21676 30108 21710
rect 30164 21676 30198 21710
rect 30254 21676 30288 21710
rect 30344 21676 30378 21710
rect 30434 21676 30468 21710
rect 30524 21676 30558 21710
rect 29984 21586 30018 21620
rect 30074 21586 30108 21620
rect 30164 21586 30198 21620
rect 30254 21586 30288 21620
rect 30344 21586 30378 21620
rect 30434 21586 30468 21620
rect 30524 21586 30558 21620
rect 29984 21496 30018 21530
rect 30074 21496 30108 21530
rect 30164 21496 30198 21530
rect 30254 21496 30288 21530
rect 30344 21496 30378 21530
rect 30434 21496 30468 21530
rect 30524 21496 30558 21530
rect 29984 21406 30018 21440
rect 30074 21406 30108 21440
rect 30164 21406 30198 21440
rect 30254 21406 30288 21440
rect 30344 21406 30378 21440
rect 30434 21406 30468 21440
rect 30524 21406 30558 21440
rect 31324 21946 31358 21980
rect 31414 21946 31448 21980
rect 31504 21946 31538 21980
rect 31594 21946 31628 21980
rect 31684 21946 31718 21980
rect 31774 21946 31808 21980
rect 31864 21946 31898 21980
rect 31324 21856 31358 21890
rect 31414 21856 31448 21890
rect 31504 21856 31538 21890
rect 31594 21856 31628 21890
rect 31684 21856 31718 21890
rect 31774 21856 31808 21890
rect 31864 21856 31898 21890
rect 31324 21766 31358 21800
rect 31414 21766 31448 21800
rect 31504 21766 31538 21800
rect 31594 21766 31628 21800
rect 31684 21766 31718 21800
rect 31774 21766 31808 21800
rect 31864 21766 31898 21800
rect 31324 21676 31358 21710
rect 31414 21676 31448 21710
rect 31504 21676 31538 21710
rect 31594 21676 31628 21710
rect 31684 21676 31718 21710
rect 31774 21676 31808 21710
rect 31864 21676 31898 21710
rect 31324 21586 31358 21620
rect 31414 21586 31448 21620
rect 31504 21586 31538 21620
rect 31594 21586 31628 21620
rect 31684 21586 31718 21620
rect 31774 21586 31808 21620
rect 31864 21586 31898 21620
rect 31324 21496 31358 21530
rect 31414 21496 31448 21530
rect 31504 21496 31538 21530
rect 31594 21496 31628 21530
rect 31684 21496 31718 21530
rect 31774 21496 31808 21530
rect 31864 21496 31898 21530
rect 31324 21406 31358 21440
rect 31414 21406 31448 21440
rect 31504 21406 31538 21440
rect 31594 21406 31628 21440
rect 31684 21406 31718 21440
rect 31774 21406 31808 21440
rect 31864 21406 31898 21440
rect 32664 21946 32698 21980
rect 32754 21946 32788 21980
rect 32844 21946 32878 21980
rect 32934 21946 32968 21980
rect 33024 21946 33058 21980
rect 33114 21946 33148 21980
rect 33204 21946 33238 21980
rect 32664 21856 32698 21890
rect 32754 21856 32788 21890
rect 32844 21856 32878 21890
rect 32934 21856 32968 21890
rect 33024 21856 33058 21890
rect 33114 21856 33148 21890
rect 33204 21856 33238 21890
rect 32664 21766 32698 21800
rect 32754 21766 32788 21800
rect 32844 21766 32878 21800
rect 32934 21766 32968 21800
rect 33024 21766 33058 21800
rect 33114 21766 33148 21800
rect 33204 21766 33238 21800
rect 32664 21676 32698 21710
rect 32754 21676 32788 21710
rect 32844 21676 32878 21710
rect 32934 21676 32968 21710
rect 33024 21676 33058 21710
rect 33114 21676 33148 21710
rect 33204 21676 33238 21710
rect 32664 21586 32698 21620
rect 32754 21586 32788 21620
rect 32844 21586 32878 21620
rect 32934 21586 32968 21620
rect 33024 21586 33058 21620
rect 33114 21586 33148 21620
rect 33204 21586 33238 21620
rect 32664 21496 32698 21530
rect 32754 21496 32788 21530
rect 32844 21496 32878 21530
rect 32934 21496 32968 21530
rect 33024 21496 33058 21530
rect 33114 21496 33148 21530
rect 33204 21496 33238 21530
rect 32664 21406 32698 21440
rect 32754 21406 32788 21440
rect 32844 21406 32878 21440
rect 32934 21406 32968 21440
rect 33024 21406 33058 21440
rect 33114 21406 33148 21440
rect 33204 21406 33238 21440
rect 34004 21946 34038 21980
rect 34094 21946 34128 21980
rect 34184 21946 34218 21980
rect 34274 21946 34308 21980
rect 34364 21946 34398 21980
rect 34454 21946 34488 21980
rect 34544 21946 34578 21980
rect 34004 21856 34038 21890
rect 34094 21856 34128 21890
rect 34184 21856 34218 21890
rect 34274 21856 34308 21890
rect 34364 21856 34398 21890
rect 34454 21856 34488 21890
rect 34544 21856 34578 21890
rect 34004 21766 34038 21800
rect 34094 21766 34128 21800
rect 34184 21766 34218 21800
rect 34274 21766 34308 21800
rect 34364 21766 34398 21800
rect 34454 21766 34488 21800
rect 34544 21766 34578 21800
rect 34004 21676 34038 21710
rect 34094 21676 34128 21710
rect 34184 21676 34218 21710
rect 34274 21676 34308 21710
rect 34364 21676 34398 21710
rect 34454 21676 34488 21710
rect 34544 21676 34578 21710
rect 34004 21586 34038 21620
rect 34094 21586 34128 21620
rect 34184 21586 34218 21620
rect 34274 21586 34308 21620
rect 34364 21586 34398 21620
rect 34454 21586 34488 21620
rect 34544 21586 34578 21620
rect 34004 21496 34038 21530
rect 34094 21496 34128 21530
rect 34184 21496 34218 21530
rect 34274 21496 34308 21530
rect 34364 21496 34398 21530
rect 34454 21496 34488 21530
rect 34544 21496 34578 21530
rect 34004 21406 34038 21440
rect 34094 21406 34128 21440
rect 34184 21406 34218 21440
rect 34274 21406 34308 21440
rect 34364 21406 34398 21440
rect 34454 21406 34488 21440
rect 34544 21406 34578 21440
rect 35344 21946 35378 21980
rect 35434 21946 35468 21980
rect 35524 21946 35558 21980
rect 35614 21946 35648 21980
rect 35704 21946 35738 21980
rect 35794 21946 35828 21980
rect 35884 21946 35918 21980
rect 35344 21856 35378 21890
rect 35434 21856 35468 21890
rect 35524 21856 35558 21890
rect 35614 21856 35648 21890
rect 35704 21856 35738 21890
rect 35794 21856 35828 21890
rect 35884 21856 35918 21890
rect 35344 21766 35378 21800
rect 35434 21766 35468 21800
rect 35524 21766 35558 21800
rect 35614 21766 35648 21800
rect 35704 21766 35738 21800
rect 35794 21766 35828 21800
rect 35884 21766 35918 21800
rect 35344 21676 35378 21710
rect 35434 21676 35468 21710
rect 35524 21676 35558 21710
rect 35614 21676 35648 21710
rect 35704 21676 35738 21710
rect 35794 21676 35828 21710
rect 35884 21676 35918 21710
rect 35344 21586 35378 21620
rect 35434 21586 35468 21620
rect 35524 21586 35558 21620
rect 35614 21586 35648 21620
rect 35704 21586 35738 21620
rect 35794 21586 35828 21620
rect 35884 21586 35918 21620
rect 35344 21496 35378 21530
rect 35434 21496 35468 21530
rect 35524 21496 35558 21530
rect 35614 21496 35648 21530
rect 35704 21496 35738 21530
rect 35794 21496 35828 21530
rect 35884 21496 35918 21530
rect 35344 21406 35378 21440
rect 35434 21406 35468 21440
rect 35524 21406 35558 21440
rect 35614 21406 35648 21440
rect 35704 21406 35738 21440
rect 35794 21406 35828 21440
rect 35884 21406 35918 21440
rect 36684 21946 36718 21980
rect 36774 21946 36808 21980
rect 36864 21946 36898 21980
rect 36954 21946 36988 21980
rect 37044 21946 37078 21980
rect 37134 21946 37168 21980
rect 37224 21946 37258 21980
rect 36684 21856 36718 21890
rect 36774 21856 36808 21890
rect 36864 21856 36898 21890
rect 36954 21856 36988 21890
rect 37044 21856 37078 21890
rect 37134 21856 37168 21890
rect 37224 21856 37258 21890
rect 36684 21766 36718 21800
rect 36774 21766 36808 21800
rect 36864 21766 36898 21800
rect 36954 21766 36988 21800
rect 37044 21766 37078 21800
rect 37134 21766 37168 21800
rect 37224 21766 37258 21800
rect 36684 21676 36718 21710
rect 36774 21676 36808 21710
rect 36864 21676 36898 21710
rect 36954 21676 36988 21710
rect 37044 21676 37078 21710
rect 37134 21676 37168 21710
rect 37224 21676 37258 21710
rect 36684 21586 36718 21620
rect 36774 21586 36808 21620
rect 36864 21586 36898 21620
rect 36954 21586 36988 21620
rect 37044 21586 37078 21620
rect 37134 21586 37168 21620
rect 37224 21586 37258 21620
rect 36684 21496 36718 21530
rect 36774 21496 36808 21530
rect 36864 21496 36898 21530
rect 36954 21496 36988 21530
rect 37044 21496 37078 21530
rect 37134 21496 37168 21530
rect 37224 21496 37258 21530
rect 36684 21406 36718 21440
rect 36774 21406 36808 21440
rect 36864 21406 36898 21440
rect 36954 21406 36988 21440
rect 37044 21406 37078 21440
rect 37134 21406 37168 21440
rect 37224 21406 37258 21440
rect 38024 21946 38058 21980
rect 38114 21946 38148 21980
rect 38204 21946 38238 21980
rect 38294 21946 38328 21980
rect 38384 21946 38418 21980
rect 38474 21946 38508 21980
rect 38564 21946 38598 21980
rect 38024 21856 38058 21890
rect 38114 21856 38148 21890
rect 38204 21856 38238 21890
rect 38294 21856 38328 21890
rect 38384 21856 38418 21890
rect 38474 21856 38508 21890
rect 38564 21856 38598 21890
rect 38024 21766 38058 21800
rect 38114 21766 38148 21800
rect 38204 21766 38238 21800
rect 38294 21766 38328 21800
rect 38384 21766 38418 21800
rect 38474 21766 38508 21800
rect 38564 21766 38598 21800
rect 38024 21676 38058 21710
rect 38114 21676 38148 21710
rect 38204 21676 38238 21710
rect 38294 21676 38328 21710
rect 38384 21676 38418 21710
rect 38474 21676 38508 21710
rect 38564 21676 38598 21710
rect 38024 21586 38058 21620
rect 38114 21586 38148 21620
rect 38204 21586 38238 21620
rect 38294 21586 38328 21620
rect 38384 21586 38418 21620
rect 38474 21586 38508 21620
rect 38564 21586 38598 21620
rect 38024 21496 38058 21530
rect 38114 21496 38148 21530
rect 38204 21496 38238 21530
rect 38294 21496 38328 21530
rect 38384 21496 38418 21530
rect 38474 21496 38508 21530
rect 38564 21496 38598 21530
rect 38024 21406 38058 21440
rect 38114 21406 38148 21440
rect 38204 21406 38238 21440
rect 38294 21406 38328 21440
rect 38384 21406 38418 21440
rect 38474 21406 38508 21440
rect 38564 21406 38598 21440
rect 23995 18587 24029 18621
rect 23995 18519 24029 18553
rect 23995 18451 24029 18485
rect 23995 18383 24029 18417
rect 23995 18315 24029 18349
rect 23995 18247 24029 18281
rect 23995 18179 24029 18213
rect 23995 18111 24029 18145
rect 23995 18043 24029 18077
rect 23995 17975 24029 18009
rect 23995 17907 24029 17941
rect 23995 17839 24029 17873
rect 23995 17771 24029 17805
rect 23995 17703 24029 17737
rect 23995 17635 24029 17669
rect 23995 17567 24029 17601
rect 23995 17499 24029 17533
rect 23995 17431 24029 17465
rect 23995 17363 24029 17397
rect 24453 18587 24487 18621
rect 24453 18519 24487 18553
rect 24453 18451 24487 18485
rect 24453 18383 24487 18417
rect 24453 18315 24487 18349
rect 24453 18247 24487 18281
rect 24453 18179 24487 18213
rect 24453 18111 24487 18145
rect 24453 18043 24487 18077
rect 24453 17975 24487 18009
rect 24453 17907 24487 17941
rect 24453 17839 24487 17873
rect 24453 17771 24487 17805
rect 24453 17703 24487 17737
rect 24453 17635 24487 17669
rect 24453 17567 24487 17601
rect 24453 17499 24487 17533
rect 24453 17431 24487 17465
rect 24453 17363 24487 17397
rect 24911 18587 24945 18621
rect 24911 18519 24945 18553
rect 24911 18451 24945 18485
rect 24911 18383 24945 18417
rect 24911 18315 24945 18349
rect 24911 18247 24945 18281
rect 24911 18179 24945 18213
rect 24911 18111 24945 18145
rect 24911 18043 24945 18077
rect 24911 17975 24945 18009
rect 24911 17907 24945 17941
rect 24911 17839 24945 17873
rect 24911 17771 24945 17805
rect 24911 17703 24945 17737
rect 24911 17635 24945 17669
rect 24911 17567 24945 17601
rect 24911 17499 24945 17533
rect 24911 17431 24945 17465
rect 24911 17363 24945 17397
rect 25369 18587 25403 18621
rect 25369 18519 25403 18553
rect 25369 18451 25403 18485
rect 25369 18383 25403 18417
rect 25369 18315 25403 18349
rect 25369 18247 25403 18281
rect 25369 18179 25403 18213
rect 25369 18111 25403 18145
rect 25369 18043 25403 18077
rect 25369 17975 25403 18009
rect 25369 17907 25403 17941
rect 25369 17839 25403 17873
rect 25369 17771 25403 17805
rect 25369 17703 25403 17737
rect 25369 17635 25403 17669
rect 25369 17567 25403 17601
rect 25369 17499 25403 17533
rect 25369 17431 25403 17465
rect 25369 17363 25403 17397
rect 25827 18587 25861 18621
rect 25827 18519 25861 18553
rect 25827 18451 25861 18485
rect 25827 18383 25861 18417
rect 25827 18315 25861 18349
rect 25827 18247 25861 18281
rect 25827 18179 25861 18213
rect 25827 18111 25861 18145
rect 25827 18043 25861 18077
rect 25827 17975 25861 18009
rect 25827 17907 25861 17941
rect 25827 17839 25861 17873
rect 25827 17771 25861 17805
rect 25827 17703 25861 17737
rect 25827 17635 25861 17669
rect 25827 17567 25861 17601
rect 25827 17499 25861 17533
rect 25827 17431 25861 17465
rect 25827 17363 25861 17397
rect 26285 18587 26319 18621
rect 26285 18519 26319 18553
rect 26285 18451 26319 18485
rect 26285 18383 26319 18417
rect 26285 18315 26319 18349
rect 26285 18247 26319 18281
rect 26285 18179 26319 18213
rect 26285 18111 26319 18145
rect 26285 18043 26319 18077
rect 26285 17975 26319 18009
rect 26285 17907 26319 17941
rect 26285 17839 26319 17873
rect 26285 17771 26319 17805
rect 26285 17703 26319 17737
rect 26285 17635 26319 17669
rect 26285 17567 26319 17601
rect 26285 17499 26319 17533
rect 26285 17431 26319 17465
rect 26285 17363 26319 17397
rect 26743 18587 26777 18621
rect 26743 18519 26777 18553
rect 26743 18451 26777 18485
rect 26743 18383 26777 18417
rect 26743 18315 26777 18349
rect 26743 18247 26777 18281
rect 26743 18179 26777 18213
rect 26743 18111 26777 18145
rect 26743 18043 26777 18077
rect 26743 17975 26777 18009
rect 26743 17907 26777 17941
rect 26743 17839 26777 17873
rect 26743 17771 26777 17805
rect 26743 17703 26777 17737
rect 26743 17635 26777 17669
rect 26743 17567 26777 17601
rect 26743 17499 26777 17533
rect 26743 17431 26777 17465
rect 26743 17363 26777 17397
rect 28644 18186 28678 18220
rect 28734 18186 28768 18220
rect 28824 18186 28858 18220
rect 28914 18186 28948 18220
rect 29004 18186 29038 18220
rect 29094 18186 29128 18220
rect 29184 18186 29218 18220
rect 28644 18096 28678 18130
rect 28734 18096 28768 18130
rect 28824 18096 28858 18130
rect 28914 18096 28948 18130
rect 29004 18096 29038 18130
rect 29094 18096 29128 18130
rect 29184 18096 29218 18130
rect 28644 18006 28678 18040
rect 28734 18006 28768 18040
rect 28824 18006 28858 18040
rect 28914 18006 28948 18040
rect 29004 18006 29038 18040
rect 29094 18006 29128 18040
rect 29184 18006 29218 18040
rect 28644 17916 28678 17950
rect 28734 17916 28768 17950
rect 28824 17916 28858 17950
rect 28914 17916 28948 17950
rect 29004 17916 29038 17950
rect 29094 17916 29128 17950
rect 29184 17916 29218 17950
rect 28644 17826 28678 17860
rect 28734 17826 28768 17860
rect 28824 17826 28858 17860
rect 28914 17826 28948 17860
rect 29004 17826 29038 17860
rect 29094 17826 29128 17860
rect 29184 17826 29218 17860
rect 28644 17736 28678 17770
rect 28734 17736 28768 17770
rect 28824 17736 28858 17770
rect 28914 17736 28948 17770
rect 29004 17736 29038 17770
rect 29094 17736 29128 17770
rect 29184 17736 29218 17770
rect 28644 17646 28678 17680
rect 28734 17646 28768 17680
rect 28824 17646 28858 17680
rect 28914 17646 28948 17680
rect 29004 17646 29038 17680
rect 29094 17646 29128 17680
rect 29184 17646 29218 17680
rect 29984 18186 30018 18220
rect 30074 18186 30108 18220
rect 30164 18186 30198 18220
rect 30254 18186 30288 18220
rect 30344 18186 30378 18220
rect 30434 18186 30468 18220
rect 30524 18186 30558 18220
rect 29984 18096 30018 18130
rect 30074 18096 30108 18130
rect 30164 18096 30198 18130
rect 30254 18096 30288 18130
rect 30344 18096 30378 18130
rect 30434 18096 30468 18130
rect 30524 18096 30558 18130
rect 29984 18006 30018 18040
rect 30074 18006 30108 18040
rect 30164 18006 30198 18040
rect 30254 18006 30288 18040
rect 30344 18006 30378 18040
rect 30434 18006 30468 18040
rect 30524 18006 30558 18040
rect 29984 17916 30018 17950
rect 30074 17916 30108 17950
rect 30164 17916 30198 17950
rect 30254 17916 30288 17950
rect 30344 17916 30378 17950
rect 30434 17916 30468 17950
rect 30524 17916 30558 17950
rect 29984 17826 30018 17860
rect 30074 17826 30108 17860
rect 30164 17826 30198 17860
rect 30254 17826 30288 17860
rect 30344 17826 30378 17860
rect 30434 17826 30468 17860
rect 30524 17826 30558 17860
rect 29984 17736 30018 17770
rect 30074 17736 30108 17770
rect 30164 17736 30198 17770
rect 30254 17736 30288 17770
rect 30344 17736 30378 17770
rect 30434 17736 30468 17770
rect 30524 17736 30558 17770
rect 29984 17646 30018 17680
rect 30074 17646 30108 17680
rect 30164 17646 30198 17680
rect 30254 17646 30288 17680
rect 30344 17646 30378 17680
rect 30434 17646 30468 17680
rect 30524 17646 30558 17680
rect 31324 18186 31358 18220
rect 31414 18186 31448 18220
rect 31504 18186 31538 18220
rect 31594 18186 31628 18220
rect 31684 18186 31718 18220
rect 31774 18186 31808 18220
rect 31864 18186 31898 18220
rect 31324 18096 31358 18130
rect 31414 18096 31448 18130
rect 31504 18096 31538 18130
rect 31594 18096 31628 18130
rect 31684 18096 31718 18130
rect 31774 18096 31808 18130
rect 31864 18096 31898 18130
rect 31324 18006 31358 18040
rect 31414 18006 31448 18040
rect 31504 18006 31538 18040
rect 31594 18006 31628 18040
rect 31684 18006 31718 18040
rect 31774 18006 31808 18040
rect 31864 18006 31898 18040
rect 31324 17916 31358 17950
rect 31414 17916 31448 17950
rect 31504 17916 31538 17950
rect 31594 17916 31628 17950
rect 31684 17916 31718 17950
rect 31774 17916 31808 17950
rect 31864 17916 31898 17950
rect 31324 17826 31358 17860
rect 31414 17826 31448 17860
rect 31504 17826 31538 17860
rect 31594 17826 31628 17860
rect 31684 17826 31718 17860
rect 31774 17826 31808 17860
rect 31864 17826 31898 17860
rect 31324 17736 31358 17770
rect 31414 17736 31448 17770
rect 31504 17736 31538 17770
rect 31594 17736 31628 17770
rect 31684 17736 31718 17770
rect 31774 17736 31808 17770
rect 31864 17736 31898 17770
rect 31324 17646 31358 17680
rect 31414 17646 31448 17680
rect 31504 17646 31538 17680
rect 31594 17646 31628 17680
rect 31684 17646 31718 17680
rect 31774 17646 31808 17680
rect 31864 17646 31898 17680
rect 32664 18186 32698 18220
rect 32754 18186 32788 18220
rect 32844 18186 32878 18220
rect 32934 18186 32968 18220
rect 33024 18186 33058 18220
rect 33114 18186 33148 18220
rect 33204 18186 33238 18220
rect 32664 18096 32698 18130
rect 32754 18096 32788 18130
rect 32844 18096 32878 18130
rect 32934 18096 32968 18130
rect 33024 18096 33058 18130
rect 33114 18096 33148 18130
rect 33204 18096 33238 18130
rect 32664 18006 32698 18040
rect 32754 18006 32788 18040
rect 32844 18006 32878 18040
rect 32934 18006 32968 18040
rect 33024 18006 33058 18040
rect 33114 18006 33148 18040
rect 33204 18006 33238 18040
rect 32664 17916 32698 17950
rect 32754 17916 32788 17950
rect 32844 17916 32878 17950
rect 32934 17916 32968 17950
rect 33024 17916 33058 17950
rect 33114 17916 33148 17950
rect 33204 17916 33238 17950
rect 32664 17826 32698 17860
rect 32754 17826 32788 17860
rect 32844 17826 32878 17860
rect 32934 17826 32968 17860
rect 33024 17826 33058 17860
rect 33114 17826 33148 17860
rect 33204 17826 33238 17860
rect 32664 17736 32698 17770
rect 32754 17736 32788 17770
rect 32844 17736 32878 17770
rect 32934 17736 32968 17770
rect 33024 17736 33058 17770
rect 33114 17736 33148 17770
rect 33204 17736 33238 17770
rect 32664 17646 32698 17680
rect 32754 17646 32788 17680
rect 32844 17646 32878 17680
rect 32934 17646 32968 17680
rect 33024 17646 33058 17680
rect 33114 17646 33148 17680
rect 33204 17646 33238 17680
rect 34004 18186 34038 18220
rect 34094 18186 34128 18220
rect 34184 18186 34218 18220
rect 34274 18186 34308 18220
rect 34364 18186 34398 18220
rect 34454 18186 34488 18220
rect 34544 18186 34578 18220
rect 34004 18096 34038 18130
rect 34094 18096 34128 18130
rect 34184 18096 34218 18130
rect 34274 18096 34308 18130
rect 34364 18096 34398 18130
rect 34454 18096 34488 18130
rect 34544 18096 34578 18130
rect 34004 18006 34038 18040
rect 34094 18006 34128 18040
rect 34184 18006 34218 18040
rect 34274 18006 34308 18040
rect 34364 18006 34398 18040
rect 34454 18006 34488 18040
rect 34544 18006 34578 18040
rect 34004 17916 34038 17950
rect 34094 17916 34128 17950
rect 34184 17916 34218 17950
rect 34274 17916 34308 17950
rect 34364 17916 34398 17950
rect 34454 17916 34488 17950
rect 34544 17916 34578 17950
rect 34004 17826 34038 17860
rect 34094 17826 34128 17860
rect 34184 17826 34218 17860
rect 34274 17826 34308 17860
rect 34364 17826 34398 17860
rect 34454 17826 34488 17860
rect 34544 17826 34578 17860
rect 34004 17736 34038 17770
rect 34094 17736 34128 17770
rect 34184 17736 34218 17770
rect 34274 17736 34308 17770
rect 34364 17736 34398 17770
rect 34454 17736 34488 17770
rect 34544 17736 34578 17770
rect 34004 17646 34038 17680
rect 34094 17646 34128 17680
rect 34184 17646 34218 17680
rect 34274 17646 34308 17680
rect 34364 17646 34398 17680
rect 34454 17646 34488 17680
rect 34544 17646 34578 17680
rect 35344 18186 35378 18220
rect 35434 18186 35468 18220
rect 35524 18186 35558 18220
rect 35614 18186 35648 18220
rect 35704 18186 35738 18220
rect 35794 18186 35828 18220
rect 35884 18186 35918 18220
rect 35344 18096 35378 18130
rect 35434 18096 35468 18130
rect 35524 18096 35558 18130
rect 35614 18096 35648 18130
rect 35704 18096 35738 18130
rect 35794 18096 35828 18130
rect 35884 18096 35918 18130
rect 35344 18006 35378 18040
rect 35434 18006 35468 18040
rect 35524 18006 35558 18040
rect 35614 18006 35648 18040
rect 35704 18006 35738 18040
rect 35794 18006 35828 18040
rect 35884 18006 35918 18040
rect 35344 17916 35378 17950
rect 35434 17916 35468 17950
rect 35524 17916 35558 17950
rect 35614 17916 35648 17950
rect 35704 17916 35738 17950
rect 35794 17916 35828 17950
rect 35884 17916 35918 17950
rect 35344 17826 35378 17860
rect 35434 17826 35468 17860
rect 35524 17826 35558 17860
rect 35614 17826 35648 17860
rect 35704 17826 35738 17860
rect 35794 17826 35828 17860
rect 35884 17826 35918 17860
rect 35344 17736 35378 17770
rect 35434 17736 35468 17770
rect 35524 17736 35558 17770
rect 35614 17736 35648 17770
rect 35704 17736 35738 17770
rect 35794 17736 35828 17770
rect 35884 17736 35918 17770
rect 35344 17646 35378 17680
rect 35434 17646 35468 17680
rect 35524 17646 35558 17680
rect 35614 17646 35648 17680
rect 35704 17646 35738 17680
rect 35794 17646 35828 17680
rect 35884 17646 35918 17680
rect 36684 18186 36718 18220
rect 36774 18186 36808 18220
rect 36864 18186 36898 18220
rect 36954 18186 36988 18220
rect 37044 18186 37078 18220
rect 37134 18186 37168 18220
rect 37224 18186 37258 18220
rect 36684 18096 36718 18130
rect 36774 18096 36808 18130
rect 36864 18096 36898 18130
rect 36954 18096 36988 18130
rect 37044 18096 37078 18130
rect 37134 18096 37168 18130
rect 37224 18096 37258 18130
rect 36684 18006 36718 18040
rect 36774 18006 36808 18040
rect 36864 18006 36898 18040
rect 36954 18006 36988 18040
rect 37044 18006 37078 18040
rect 37134 18006 37168 18040
rect 37224 18006 37258 18040
rect 36684 17916 36718 17950
rect 36774 17916 36808 17950
rect 36864 17916 36898 17950
rect 36954 17916 36988 17950
rect 37044 17916 37078 17950
rect 37134 17916 37168 17950
rect 37224 17916 37258 17950
rect 36684 17826 36718 17860
rect 36774 17826 36808 17860
rect 36864 17826 36898 17860
rect 36954 17826 36988 17860
rect 37044 17826 37078 17860
rect 37134 17826 37168 17860
rect 37224 17826 37258 17860
rect 36684 17736 36718 17770
rect 36774 17736 36808 17770
rect 36864 17736 36898 17770
rect 36954 17736 36988 17770
rect 37044 17736 37078 17770
rect 37134 17736 37168 17770
rect 37224 17736 37258 17770
rect 36684 17646 36718 17680
rect 36774 17646 36808 17680
rect 36864 17646 36898 17680
rect 36954 17646 36988 17680
rect 37044 17646 37078 17680
rect 37134 17646 37168 17680
rect 37224 17646 37258 17680
rect 38024 18186 38058 18220
rect 38114 18186 38148 18220
rect 38204 18186 38238 18220
rect 38294 18186 38328 18220
rect 38384 18186 38418 18220
rect 38474 18186 38508 18220
rect 38564 18186 38598 18220
rect 38024 18096 38058 18130
rect 38114 18096 38148 18130
rect 38204 18096 38238 18130
rect 38294 18096 38328 18130
rect 38384 18096 38418 18130
rect 38474 18096 38508 18130
rect 38564 18096 38598 18130
rect 38024 18006 38058 18040
rect 38114 18006 38148 18040
rect 38204 18006 38238 18040
rect 38294 18006 38328 18040
rect 38384 18006 38418 18040
rect 38474 18006 38508 18040
rect 38564 18006 38598 18040
rect 38024 17916 38058 17950
rect 38114 17916 38148 17950
rect 38204 17916 38238 17950
rect 38294 17916 38328 17950
rect 38384 17916 38418 17950
rect 38474 17916 38508 17950
rect 38564 17916 38598 17950
rect 38024 17826 38058 17860
rect 38114 17826 38148 17860
rect 38204 17826 38238 17860
rect 38294 17826 38328 17860
rect 38384 17826 38418 17860
rect 38474 17826 38508 17860
rect 38564 17826 38598 17860
rect 38024 17736 38058 17770
rect 38114 17736 38148 17770
rect 38204 17736 38238 17770
rect 38294 17736 38328 17770
rect 38384 17736 38418 17770
rect 38474 17736 38508 17770
rect 38564 17736 38598 17770
rect 38024 17646 38058 17680
rect 38114 17646 38148 17680
rect 38204 17646 38238 17680
rect 38294 17646 38328 17680
rect 38384 17646 38418 17680
rect 38474 17646 38508 17680
rect 38564 17646 38598 17680
rect 28644 14426 28678 14460
rect 28734 14426 28768 14460
rect 28824 14426 28858 14460
rect 28914 14426 28948 14460
rect 29004 14426 29038 14460
rect 29094 14426 29128 14460
rect 29184 14426 29218 14460
rect 28644 14336 28678 14370
rect 28734 14336 28768 14370
rect 28824 14336 28858 14370
rect 28914 14336 28948 14370
rect 29004 14336 29038 14370
rect 29094 14336 29128 14370
rect 29184 14336 29218 14370
rect 28644 14246 28678 14280
rect 28734 14246 28768 14280
rect 28824 14246 28858 14280
rect 28914 14246 28948 14280
rect 29004 14246 29038 14280
rect 29094 14246 29128 14280
rect 29184 14246 29218 14280
rect 28644 14156 28678 14190
rect 28734 14156 28768 14190
rect 28824 14156 28858 14190
rect 28914 14156 28948 14190
rect 29004 14156 29038 14190
rect 29094 14156 29128 14190
rect 29184 14156 29218 14190
rect 28644 14066 28678 14100
rect 28734 14066 28768 14100
rect 28824 14066 28858 14100
rect 28914 14066 28948 14100
rect 29004 14066 29038 14100
rect 29094 14066 29128 14100
rect 29184 14066 29218 14100
rect 28644 13976 28678 14010
rect 28734 13976 28768 14010
rect 28824 13976 28858 14010
rect 28914 13976 28948 14010
rect 29004 13976 29038 14010
rect 29094 13976 29128 14010
rect 29184 13976 29218 14010
rect 28644 13886 28678 13920
rect 28734 13886 28768 13920
rect 28824 13886 28858 13920
rect 28914 13886 28948 13920
rect 29004 13886 29038 13920
rect 29094 13886 29128 13920
rect 29184 13886 29218 13920
rect 29984 14426 30018 14460
rect 30074 14426 30108 14460
rect 30164 14426 30198 14460
rect 30254 14426 30288 14460
rect 30344 14426 30378 14460
rect 30434 14426 30468 14460
rect 30524 14426 30558 14460
rect 29984 14336 30018 14370
rect 30074 14336 30108 14370
rect 30164 14336 30198 14370
rect 30254 14336 30288 14370
rect 30344 14336 30378 14370
rect 30434 14336 30468 14370
rect 30524 14336 30558 14370
rect 29984 14246 30018 14280
rect 30074 14246 30108 14280
rect 30164 14246 30198 14280
rect 30254 14246 30288 14280
rect 30344 14246 30378 14280
rect 30434 14246 30468 14280
rect 30524 14246 30558 14280
rect 29984 14156 30018 14190
rect 30074 14156 30108 14190
rect 30164 14156 30198 14190
rect 30254 14156 30288 14190
rect 30344 14156 30378 14190
rect 30434 14156 30468 14190
rect 30524 14156 30558 14190
rect 29984 14066 30018 14100
rect 30074 14066 30108 14100
rect 30164 14066 30198 14100
rect 30254 14066 30288 14100
rect 30344 14066 30378 14100
rect 30434 14066 30468 14100
rect 30524 14066 30558 14100
rect 29984 13976 30018 14010
rect 30074 13976 30108 14010
rect 30164 13976 30198 14010
rect 30254 13976 30288 14010
rect 30344 13976 30378 14010
rect 30434 13976 30468 14010
rect 30524 13976 30558 14010
rect 29984 13886 30018 13920
rect 30074 13886 30108 13920
rect 30164 13886 30198 13920
rect 30254 13886 30288 13920
rect 30344 13886 30378 13920
rect 30434 13886 30468 13920
rect 30524 13886 30558 13920
rect 31324 14426 31358 14460
rect 31414 14426 31448 14460
rect 31504 14426 31538 14460
rect 31594 14426 31628 14460
rect 31684 14426 31718 14460
rect 31774 14426 31808 14460
rect 31864 14426 31898 14460
rect 31324 14336 31358 14370
rect 31414 14336 31448 14370
rect 31504 14336 31538 14370
rect 31594 14336 31628 14370
rect 31684 14336 31718 14370
rect 31774 14336 31808 14370
rect 31864 14336 31898 14370
rect 31324 14246 31358 14280
rect 31414 14246 31448 14280
rect 31504 14246 31538 14280
rect 31594 14246 31628 14280
rect 31684 14246 31718 14280
rect 31774 14246 31808 14280
rect 31864 14246 31898 14280
rect 31324 14156 31358 14190
rect 31414 14156 31448 14190
rect 31504 14156 31538 14190
rect 31594 14156 31628 14190
rect 31684 14156 31718 14190
rect 31774 14156 31808 14190
rect 31864 14156 31898 14190
rect 31324 14066 31358 14100
rect 31414 14066 31448 14100
rect 31504 14066 31538 14100
rect 31594 14066 31628 14100
rect 31684 14066 31718 14100
rect 31774 14066 31808 14100
rect 31864 14066 31898 14100
rect 31324 13976 31358 14010
rect 31414 13976 31448 14010
rect 31504 13976 31538 14010
rect 31594 13976 31628 14010
rect 31684 13976 31718 14010
rect 31774 13976 31808 14010
rect 31864 13976 31898 14010
rect 31324 13886 31358 13920
rect 31414 13886 31448 13920
rect 31504 13886 31538 13920
rect 31594 13886 31628 13920
rect 31684 13886 31718 13920
rect 31774 13886 31808 13920
rect 31864 13886 31898 13920
rect 32664 14426 32698 14460
rect 32754 14426 32788 14460
rect 32844 14426 32878 14460
rect 32934 14426 32968 14460
rect 33024 14426 33058 14460
rect 33114 14426 33148 14460
rect 33204 14426 33238 14460
rect 32664 14336 32698 14370
rect 32754 14336 32788 14370
rect 32844 14336 32878 14370
rect 32934 14336 32968 14370
rect 33024 14336 33058 14370
rect 33114 14336 33148 14370
rect 33204 14336 33238 14370
rect 32664 14246 32698 14280
rect 32754 14246 32788 14280
rect 32844 14246 32878 14280
rect 32934 14246 32968 14280
rect 33024 14246 33058 14280
rect 33114 14246 33148 14280
rect 33204 14246 33238 14280
rect 32664 14156 32698 14190
rect 32754 14156 32788 14190
rect 32844 14156 32878 14190
rect 32934 14156 32968 14190
rect 33024 14156 33058 14190
rect 33114 14156 33148 14190
rect 33204 14156 33238 14190
rect 32664 14066 32698 14100
rect 32754 14066 32788 14100
rect 32844 14066 32878 14100
rect 32934 14066 32968 14100
rect 33024 14066 33058 14100
rect 33114 14066 33148 14100
rect 33204 14066 33238 14100
rect 32664 13976 32698 14010
rect 32754 13976 32788 14010
rect 32844 13976 32878 14010
rect 32934 13976 32968 14010
rect 33024 13976 33058 14010
rect 33114 13976 33148 14010
rect 33204 13976 33238 14010
rect 32664 13886 32698 13920
rect 32754 13886 32788 13920
rect 32844 13886 32878 13920
rect 32934 13886 32968 13920
rect 33024 13886 33058 13920
rect 33114 13886 33148 13920
rect 33204 13886 33238 13920
rect 34004 14426 34038 14460
rect 34094 14426 34128 14460
rect 34184 14426 34218 14460
rect 34274 14426 34308 14460
rect 34364 14426 34398 14460
rect 34454 14426 34488 14460
rect 34544 14426 34578 14460
rect 34004 14336 34038 14370
rect 34094 14336 34128 14370
rect 34184 14336 34218 14370
rect 34274 14336 34308 14370
rect 34364 14336 34398 14370
rect 34454 14336 34488 14370
rect 34544 14336 34578 14370
rect 34004 14246 34038 14280
rect 34094 14246 34128 14280
rect 34184 14246 34218 14280
rect 34274 14246 34308 14280
rect 34364 14246 34398 14280
rect 34454 14246 34488 14280
rect 34544 14246 34578 14280
rect 34004 14156 34038 14190
rect 34094 14156 34128 14190
rect 34184 14156 34218 14190
rect 34274 14156 34308 14190
rect 34364 14156 34398 14190
rect 34454 14156 34488 14190
rect 34544 14156 34578 14190
rect 34004 14066 34038 14100
rect 34094 14066 34128 14100
rect 34184 14066 34218 14100
rect 34274 14066 34308 14100
rect 34364 14066 34398 14100
rect 34454 14066 34488 14100
rect 34544 14066 34578 14100
rect 34004 13976 34038 14010
rect 34094 13976 34128 14010
rect 34184 13976 34218 14010
rect 34274 13976 34308 14010
rect 34364 13976 34398 14010
rect 34454 13976 34488 14010
rect 34544 13976 34578 14010
rect 34004 13886 34038 13920
rect 34094 13886 34128 13920
rect 34184 13886 34218 13920
rect 34274 13886 34308 13920
rect 34364 13886 34398 13920
rect 34454 13886 34488 13920
rect 34544 13886 34578 13920
rect 35344 14426 35378 14460
rect 35434 14426 35468 14460
rect 35524 14426 35558 14460
rect 35614 14426 35648 14460
rect 35704 14426 35738 14460
rect 35794 14426 35828 14460
rect 35884 14426 35918 14460
rect 35344 14336 35378 14370
rect 35434 14336 35468 14370
rect 35524 14336 35558 14370
rect 35614 14336 35648 14370
rect 35704 14336 35738 14370
rect 35794 14336 35828 14370
rect 35884 14336 35918 14370
rect 35344 14246 35378 14280
rect 35434 14246 35468 14280
rect 35524 14246 35558 14280
rect 35614 14246 35648 14280
rect 35704 14246 35738 14280
rect 35794 14246 35828 14280
rect 35884 14246 35918 14280
rect 35344 14156 35378 14190
rect 35434 14156 35468 14190
rect 35524 14156 35558 14190
rect 35614 14156 35648 14190
rect 35704 14156 35738 14190
rect 35794 14156 35828 14190
rect 35884 14156 35918 14190
rect 35344 14066 35378 14100
rect 35434 14066 35468 14100
rect 35524 14066 35558 14100
rect 35614 14066 35648 14100
rect 35704 14066 35738 14100
rect 35794 14066 35828 14100
rect 35884 14066 35918 14100
rect 35344 13976 35378 14010
rect 35434 13976 35468 14010
rect 35524 13976 35558 14010
rect 35614 13976 35648 14010
rect 35704 13976 35738 14010
rect 35794 13976 35828 14010
rect 35884 13976 35918 14010
rect 35344 13886 35378 13920
rect 35434 13886 35468 13920
rect 35524 13886 35558 13920
rect 35614 13886 35648 13920
rect 35704 13886 35738 13920
rect 35794 13886 35828 13920
rect 35884 13886 35918 13920
rect 36684 14426 36718 14460
rect 36774 14426 36808 14460
rect 36864 14426 36898 14460
rect 36954 14426 36988 14460
rect 37044 14426 37078 14460
rect 37134 14426 37168 14460
rect 37224 14426 37258 14460
rect 36684 14336 36718 14370
rect 36774 14336 36808 14370
rect 36864 14336 36898 14370
rect 36954 14336 36988 14370
rect 37044 14336 37078 14370
rect 37134 14336 37168 14370
rect 37224 14336 37258 14370
rect 36684 14246 36718 14280
rect 36774 14246 36808 14280
rect 36864 14246 36898 14280
rect 36954 14246 36988 14280
rect 37044 14246 37078 14280
rect 37134 14246 37168 14280
rect 37224 14246 37258 14280
rect 36684 14156 36718 14190
rect 36774 14156 36808 14190
rect 36864 14156 36898 14190
rect 36954 14156 36988 14190
rect 37044 14156 37078 14190
rect 37134 14156 37168 14190
rect 37224 14156 37258 14190
rect 36684 14066 36718 14100
rect 36774 14066 36808 14100
rect 36864 14066 36898 14100
rect 36954 14066 36988 14100
rect 37044 14066 37078 14100
rect 37134 14066 37168 14100
rect 37224 14066 37258 14100
rect 36684 13976 36718 14010
rect 36774 13976 36808 14010
rect 36864 13976 36898 14010
rect 36954 13976 36988 14010
rect 37044 13976 37078 14010
rect 37134 13976 37168 14010
rect 37224 13976 37258 14010
rect 36684 13886 36718 13920
rect 36774 13886 36808 13920
rect 36864 13886 36898 13920
rect 36954 13886 36988 13920
rect 37044 13886 37078 13920
rect 37134 13886 37168 13920
rect 37224 13886 37258 13920
rect 38024 14426 38058 14460
rect 38114 14426 38148 14460
rect 38204 14426 38238 14460
rect 38294 14426 38328 14460
rect 38384 14426 38418 14460
rect 38474 14426 38508 14460
rect 38564 14426 38598 14460
rect 38024 14336 38058 14370
rect 38114 14336 38148 14370
rect 38204 14336 38238 14370
rect 38294 14336 38328 14370
rect 38384 14336 38418 14370
rect 38474 14336 38508 14370
rect 38564 14336 38598 14370
rect 38024 14246 38058 14280
rect 38114 14246 38148 14280
rect 38204 14246 38238 14280
rect 38294 14246 38328 14280
rect 38384 14246 38418 14280
rect 38474 14246 38508 14280
rect 38564 14246 38598 14280
rect 38024 14156 38058 14190
rect 38114 14156 38148 14190
rect 38204 14156 38238 14190
rect 38294 14156 38328 14190
rect 38384 14156 38418 14190
rect 38474 14156 38508 14190
rect 38564 14156 38598 14190
rect 38024 14066 38058 14100
rect 38114 14066 38148 14100
rect 38204 14066 38238 14100
rect 38294 14066 38328 14100
rect 38384 14066 38418 14100
rect 38474 14066 38508 14100
rect 38564 14066 38598 14100
rect 38024 13976 38058 14010
rect 38114 13976 38148 14010
rect 38204 13976 38238 14010
rect 38294 13976 38328 14010
rect 38384 13976 38418 14010
rect 38474 13976 38508 14010
rect 38564 13976 38598 14010
rect 38024 13886 38058 13920
rect 38114 13886 38148 13920
rect 38204 13886 38238 13920
rect 38294 13886 38328 13920
rect 38384 13886 38418 13920
rect 38474 13886 38508 13920
rect 38564 13886 38598 13920
<< psubdiff >>
rect 5924 39709 5964 39752
rect 5924 39675 5927 39709
rect 5961 39675 5964 39709
rect 5924 39632 5964 39675
rect 30050 37341 39378 37376
rect 30050 37318 30180 37341
rect 30050 37284 30084 37318
rect 30118 37307 30180 37318
rect 30214 37307 30270 37341
rect 30304 37307 30360 37341
rect 30394 37307 30450 37341
rect 30484 37307 30540 37341
rect 30574 37307 30630 37341
rect 30664 37307 30720 37341
rect 30754 37307 30810 37341
rect 30844 37307 30900 37341
rect 30934 37307 30990 37341
rect 31024 37307 31080 37341
rect 31114 37307 31170 37341
rect 31204 37318 31520 37341
rect 31204 37307 31271 37318
rect 30118 37284 31271 37307
rect 31305 37284 31424 37318
rect 31458 37307 31520 37318
rect 31554 37307 31610 37341
rect 31644 37307 31700 37341
rect 31734 37307 31790 37341
rect 31824 37307 31880 37341
rect 31914 37307 31970 37341
rect 32004 37307 32060 37341
rect 32094 37307 32150 37341
rect 32184 37307 32240 37341
rect 32274 37307 32330 37341
rect 32364 37307 32420 37341
rect 32454 37307 32510 37341
rect 32544 37318 32860 37341
rect 32544 37307 32611 37318
rect 31458 37284 32611 37307
rect 32645 37284 32764 37318
rect 32798 37307 32860 37318
rect 32894 37307 32950 37341
rect 32984 37307 33040 37341
rect 33074 37307 33130 37341
rect 33164 37307 33220 37341
rect 33254 37307 33310 37341
rect 33344 37307 33400 37341
rect 33434 37307 33490 37341
rect 33524 37307 33580 37341
rect 33614 37307 33670 37341
rect 33704 37307 33760 37341
rect 33794 37307 33850 37341
rect 33884 37318 34200 37341
rect 33884 37307 33951 37318
rect 32798 37284 33951 37307
rect 33985 37284 34104 37318
rect 34138 37307 34200 37318
rect 34234 37307 34290 37341
rect 34324 37307 34380 37341
rect 34414 37307 34470 37341
rect 34504 37307 34560 37341
rect 34594 37307 34650 37341
rect 34684 37307 34740 37341
rect 34774 37307 34830 37341
rect 34864 37307 34920 37341
rect 34954 37307 35010 37341
rect 35044 37307 35100 37341
rect 35134 37307 35190 37341
rect 35224 37318 35540 37341
rect 35224 37307 35291 37318
rect 34138 37284 35291 37307
rect 35325 37284 35444 37318
rect 35478 37307 35540 37318
rect 35574 37307 35630 37341
rect 35664 37307 35720 37341
rect 35754 37307 35810 37341
rect 35844 37307 35900 37341
rect 35934 37307 35990 37341
rect 36024 37307 36080 37341
rect 36114 37307 36170 37341
rect 36204 37307 36260 37341
rect 36294 37307 36350 37341
rect 36384 37307 36440 37341
rect 36474 37307 36530 37341
rect 36564 37318 36880 37341
rect 36564 37307 36631 37318
rect 35478 37284 36631 37307
rect 36665 37284 36784 37318
rect 36818 37307 36880 37318
rect 36914 37307 36970 37341
rect 37004 37307 37060 37341
rect 37094 37307 37150 37341
rect 37184 37307 37240 37341
rect 37274 37307 37330 37341
rect 37364 37307 37420 37341
rect 37454 37307 37510 37341
rect 37544 37307 37600 37341
rect 37634 37307 37690 37341
rect 37724 37307 37780 37341
rect 37814 37307 37870 37341
rect 37904 37318 38220 37341
rect 37904 37307 37971 37318
rect 36818 37284 37971 37307
rect 38005 37284 38124 37318
rect 38158 37307 38220 37318
rect 38254 37307 38310 37341
rect 38344 37307 38400 37341
rect 38434 37307 38490 37341
rect 38524 37307 38580 37341
rect 38614 37307 38670 37341
rect 38704 37307 38760 37341
rect 38794 37307 38850 37341
rect 38884 37307 38940 37341
rect 38974 37307 39030 37341
rect 39064 37307 39120 37341
rect 39154 37307 39210 37341
rect 39244 37318 39378 37341
rect 39244 37307 39311 37318
rect 38158 37284 39311 37307
rect 39345 37284 39378 37318
rect 30050 37275 39378 37284
rect 30050 37228 30151 37275
rect 30050 37194 30084 37228
rect 30118 37194 30151 37228
rect 31237 37228 31491 37275
rect 30050 37138 30151 37194
rect 30050 37104 30084 37138
rect 30118 37104 30151 37138
rect 30050 37048 30151 37104
rect 30050 37014 30084 37048
rect 30118 37014 30151 37048
rect 30050 36958 30151 37014
rect 30050 36924 30084 36958
rect 30118 36924 30151 36958
rect 30050 36868 30151 36924
rect 30050 36834 30084 36868
rect 30118 36834 30151 36868
rect 30050 36778 30151 36834
rect 30050 36744 30084 36778
rect 30118 36744 30151 36778
rect 30050 36688 30151 36744
rect 30050 36654 30084 36688
rect 30118 36654 30151 36688
rect 30050 36598 30151 36654
rect 30050 36564 30084 36598
rect 30118 36564 30151 36598
rect 30050 36508 30151 36564
rect 30050 36474 30084 36508
rect 30118 36474 30151 36508
rect 30050 36418 30151 36474
rect 30050 36384 30084 36418
rect 30118 36384 30151 36418
rect 30050 36328 30151 36384
rect 30050 36294 30084 36328
rect 30118 36294 30151 36328
rect 30050 36238 30151 36294
rect 31237 37194 31271 37228
rect 31305 37194 31424 37228
rect 31458 37194 31491 37228
rect 32577 37228 32831 37275
rect 31237 37138 31491 37194
rect 31237 37104 31271 37138
rect 31305 37104 31424 37138
rect 31458 37104 31491 37138
rect 31237 37048 31491 37104
rect 31237 37014 31271 37048
rect 31305 37014 31424 37048
rect 31458 37014 31491 37048
rect 31237 36958 31491 37014
rect 31237 36924 31271 36958
rect 31305 36924 31424 36958
rect 31458 36924 31491 36958
rect 31237 36868 31491 36924
rect 31237 36834 31271 36868
rect 31305 36834 31424 36868
rect 31458 36834 31491 36868
rect 31237 36778 31491 36834
rect 31237 36744 31271 36778
rect 31305 36744 31424 36778
rect 31458 36744 31491 36778
rect 31237 36688 31491 36744
rect 31237 36654 31271 36688
rect 31305 36654 31424 36688
rect 31458 36654 31491 36688
rect 31237 36598 31491 36654
rect 31237 36564 31271 36598
rect 31305 36564 31424 36598
rect 31458 36564 31491 36598
rect 31237 36508 31491 36564
rect 31237 36474 31271 36508
rect 31305 36474 31424 36508
rect 31458 36474 31491 36508
rect 31237 36418 31491 36474
rect 31237 36384 31271 36418
rect 31305 36384 31424 36418
rect 31458 36384 31491 36418
rect 31237 36328 31491 36384
rect 31237 36294 31271 36328
rect 31305 36294 31424 36328
rect 31458 36294 31491 36328
rect 30050 36204 30084 36238
rect 30118 36204 30151 36238
rect 30050 36189 30151 36204
rect 31237 36238 31491 36294
rect 32577 37194 32611 37228
rect 32645 37194 32764 37228
rect 32798 37194 32831 37228
rect 33917 37228 34171 37275
rect 32577 37138 32831 37194
rect 32577 37104 32611 37138
rect 32645 37104 32764 37138
rect 32798 37104 32831 37138
rect 32577 37048 32831 37104
rect 32577 37014 32611 37048
rect 32645 37014 32764 37048
rect 32798 37014 32831 37048
rect 32577 36958 32831 37014
rect 32577 36924 32611 36958
rect 32645 36924 32764 36958
rect 32798 36924 32831 36958
rect 32577 36868 32831 36924
rect 32577 36834 32611 36868
rect 32645 36834 32764 36868
rect 32798 36834 32831 36868
rect 32577 36778 32831 36834
rect 32577 36744 32611 36778
rect 32645 36744 32764 36778
rect 32798 36744 32831 36778
rect 32577 36688 32831 36744
rect 32577 36654 32611 36688
rect 32645 36654 32764 36688
rect 32798 36654 32831 36688
rect 32577 36598 32831 36654
rect 32577 36564 32611 36598
rect 32645 36564 32764 36598
rect 32798 36564 32831 36598
rect 32577 36508 32831 36564
rect 32577 36474 32611 36508
rect 32645 36474 32764 36508
rect 32798 36474 32831 36508
rect 32577 36418 32831 36474
rect 32577 36384 32611 36418
rect 32645 36384 32764 36418
rect 32798 36384 32831 36418
rect 32577 36328 32831 36384
rect 32577 36294 32611 36328
rect 32645 36294 32764 36328
rect 32798 36294 32831 36328
rect 31237 36204 31271 36238
rect 31305 36204 31424 36238
rect 31458 36204 31491 36238
rect 31237 36189 31491 36204
rect 32577 36238 32831 36294
rect 33917 37194 33951 37228
rect 33985 37194 34104 37228
rect 34138 37194 34171 37228
rect 35257 37228 35511 37275
rect 33917 37138 34171 37194
rect 33917 37104 33951 37138
rect 33985 37104 34104 37138
rect 34138 37104 34171 37138
rect 33917 37048 34171 37104
rect 33917 37014 33951 37048
rect 33985 37014 34104 37048
rect 34138 37014 34171 37048
rect 33917 36958 34171 37014
rect 33917 36924 33951 36958
rect 33985 36924 34104 36958
rect 34138 36924 34171 36958
rect 33917 36868 34171 36924
rect 33917 36834 33951 36868
rect 33985 36834 34104 36868
rect 34138 36834 34171 36868
rect 33917 36778 34171 36834
rect 33917 36744 33951 36778
rect 33985 36744 34104 36778
rect 34138 36744 34171 36778
rect 33917 36688 34171 36744
rect 33917 36654 33951 36688
rect 33985 36654 34104 36688
rect 34138 36654 34171 36688
rect 33917 36598 34171 36654
rect 33917 36564 33951 36598
rect 33985 36564 34104 36598
rect 34138 36564 34171 36598
rect 33917 36508 34171 36564
rect 33917 36474 33951 36508
rect 33985 36474 34104 36508
rect 34138 36474 34171 36508
rect 33917 36418 34171 36474
rect 33917 36384 33951 36418
rect 33985 36384 34104 36418
rect 34138 36384 34171 36418
rect 33917 36328 34171 36384
rect 33917 36294 33951 36328
rect 33985 36294 34104 36328
rect 34138 36294 34171 36328
rect 32577 36204 32611 36238
rect 32645 36204 32764 36238
rect 32798 36204 32831 36238
rect 32577 36189 32831 36204
rect 33917 36238 34171 36294
rect 35257 37194 35291 37228
rect 35325 37194 35444 37228
rect 35478 37194 35511 37228
rect 36597 37228 36851 37275
rect 35257 37138 35511 37194
rect 35257 37104 35291 37138
rect 35325 37104 35444 37138
rect 35478 37104 35511 37138
rect 35257 37048 35511 37104
rect 35257 37014 35291 37048
rect 35325 37014 35444 37048
rect 35478 37014 35511 37048
rect 35257 36958 35511 37014
rect 35257 36924 35291 36958
rect 35325 36924 35444 36958
rect 35478 36924 35511 36958
rect 35257 36868 35511 36924
rect 35257 36834 35291 36868
rect 35325 36834 35444 36868
rect 35478 36834 35511 36868
rect 35257 36778 35511 36834
rect 35257 36744 35291 36778
rect 35325 36744 35444 36778
rect 35478 36744 35511 36778
rect 35257 36688 35511 36744
rect 35257 36654 35291 36688
rect 35325 36654 35444 36688
rect 35478 36654 35511 36688
rect 35257 36598 35511 36654
rect 35257 36564 35291 36598
rect 35325 36564 35444 36598
rect 35478 36564 35511 36598
rect 35257 36508 35511 36564
rect 35257 36474 35291 36508
rect 35325 36474 35444 36508
rect 35478 36474 35511 36508
rect 35257 36418 35511 36474
rect 35257 36384 35291 36418
rect 35325 36384 35444 36418
rect 35478 36384 35511 36418
rect 35257 36328 35511 36384
rect 35257 36294 35291 36328
rect 35325 36294 35444 36328
rect 35478 36294 35511 36328
rect 33917 36204 33951 36238
rect 33985 36204 34104 36238
rect 34138 36204 34171 36238
rect 33917 36189 34171 36204
rect 35257 36238 35511 36294
rect 36597 37194 36631 37228
rect 36665 37194 36784 37228
rect 36818 37194 36851 37228
rect 37937 37228 38191 37275
rect 36597 37138 36851 37194
rect 36597 37104 36631 37138
rect 36665 37104 36784 37138
rect 36818 37104 36851 37138
rect 36597 37048 36851 37104
rect 36597 37014 36631 37048
rect 36665 37014 36784 37048
rect 36818 37014 36851 37048
rect 36597 36958 36851 37014
rect 36597 36924 36631 36958
rect 36665 36924 36784 36958
rect 36818 36924 36851 36958
rect 36597 36868 36851 36924
rect 36597 36834 36631 36868
rect 36665 36834 36784 36868
rect 36818 36834 36851 36868
rect 36597 36778 36851 36834
rect 36597 36744 36631 36778
rect 36665 36744 36784 36778
rect 36818 36744 36851 36778
rect 36597 36688 36851 36744
rect 36597 36654 36631 36688
rect 36665 36654 36784 36688
rect 36818 36654 36851 36688
rect 36597 36598 36851 36654
rect 36597 36564 36631 36598
rect 36665 36564 36784 36598
rect 36818 36564 36851 36598
rect 36597 36508 36851 36564
rect 36597 36474 36631 36508
rect 36665 36474 36784 36508
rect 36818 36474 36851 36508
rect 36597 36418 36851 36474
rect 36597 36384 36631 36418
rect 36665 36384 36784 36418
rect 36818 36384 36851 36418
rect 36597 36328 36851 36384
rect 36597 36294 36631 36328
rect 36665 36294 36784 36328
rect 36818 36294 36851 36328
rect 35257 36204 35291 36238
rect 35325 36204 35444 36238
rect 35478 36204 35511 36238
rect 35257 36189 35511 36204
rect 36597 36238 36851 36294
rect 37937 37194 37971 37228
rect 38005 37194 38124 37228
rect 38158 37194 38191 37228
rect 39277 37228 39378 37275
rect 37937 37138 38191 37194
rect 37937 37104 37971 37138
rect 38005 37104 38124 37138
rect 38158 37104 38191 37138
rect 37937 37048 38191 37104
rect 37937 37014 37971 37048
rect 38005 37014 38124 37048
rect 38158 37014 38191 37048
rect 37937 36958 38191 37014
rect 37937 36924 37971 36958
rect 38005 36924 38124 36958
rect 38158 36924 38191 36958
rect 37937 36868 38191 36924
rect 37937 36834 37971 36868
rect 38005 36834 38124 36868
rect 38158 36834 38191 36868
rect 37937 36778 38191 36834
rect 37937 36744 37971 36778
rect 38005 36744 38124 36778
rect 38158 36744 38191 36778
rect 37937 36688 38191 36744
rect 37937 36654 37971 36688
rect 38005 36654 38124 36688
rect 38158 36654 38191 36688
rect 37937 36598 38191 36654
rect 37937 36564 37971 36598
rect 38005 36564 38124 36598
rect 38158 36564 38191 36598
rect 37937 36508 38191 36564
rect 37937 36474 37971 36508
rect 38005 36474 38124 36508
rect 38158 36474 38191 36508
rect 37937 36418 38191 36474
rect 37937 36384 37971 36418
rect 38005 36384 38124 36418
rect 38158 36384 38191 36418
rect 37937 36328 38191 36384
rect 37937 36294 37971 36328
rect 38005 36294 38124 36328
rect 38158 36294 38191 36328
rect 36597 36204 36631 36238
rect 36665 36204 36784 36238
rect 36818 36204 36851 36238
rect 36597 36189 36851 36204
rect 37937 36238 38191 36294
rect 39277 37194 39311 37228
rect 39345 37194 39378 37228
rect 39277 37138 39378 37194
rect 39277 37104 39311 37138
rect 39345 37104 39378 37138
rect 39277 37048 39378 37104
rect 39277 37014 39311 37048
rect 39345 37014 39378 37048
rect 39277 36958 39378 37014
rect 39277 36924 39311 36958
rect 39345 36924 39378 36958
rect 39277 36868 39378 36924
rect 39277 36834 39311 36868
rect 39345 36834 39378 36868
rect 39277 36778 39378 36834
rect 39277 36744 39311 36778
rect 39345 36744 39378 36778
rect 39277 36688 39378 36744
rect 39277 36654 39311 36688
rect 39345 36654 39378 36688
rect 39277 36598 39378 36654
rect 39277 36564 39311 36598
rect 39345 36564 39378 36598
rect 40658 36723 41274 36762
rect 40658 36621 40745 36723
rect 41187 36621 41274 36723
rect 40658 36582 41274 36621
rect 39277 36508 39378 36564
rect 39277 36474 39311 36508
rect 39345 36474 39378 36508
rect 39277 36418 39378 36474
rect 39277 36384 39311 36418
rect 39345 36384 39378 36418
rect 39277 36328 39378 36384
rect 39277 36294 39311 36328
rect 39345 36294 39378 36328
rect 37937 36204 37971 36238
rect 38005 36204 38124 36238
rect 38158 36204 38191 36238
rect 37937 36189 38191 36204
rect 39277 36238 39378 36294
rect 39277 36204 39311 36238
rect 39345 36204 39378 36238
rect 39277 36189 39378 36204
rect 30050 36154 39378 36189
rect 30050 36120 30180 36154
rect 30214 36120 30270 36154
rect 30304 36120 30360 36154
rect 30394 36120 30450 36154
rect 30484 36120 30540 36154
rect 30574 36120 30630 36154
rect 30664 36120 30720 36154
rect 30754 36120 30810 36154
rect 30844 36120 30900 36154
rect 30934 36120 30990 36154
rect 31024 36120 31080 36154
rect 31114 36120 31170 36154
rect 31204 36120 31520 36154
rect 31554 36120 31610 36154
rect 31644 36120 31700 36154
rect 31734 36120 31790 36154
rect 31824 36120 31880 36154
rect 31914 36120 31970 36154
rect 32004 36120 32060 36154
rect 32094 36120 32150 36154
rect 32184 36120 32240 36154
rect 32274 36120 32330 36154
rect 32364 36120 32420 36154
rect 32454 36120 32510 36154
rect 32544 36120 32860 36154
rect 32894 36120 32950 36154
rect 32984 36120 33040 36154
rect 33074 36120 33130 36154
rect 33164 36120 33220 36154
rect 33254 36120 33310 36154
rect 33344 36120 33400 36154
rect 33434 36120 33490 36154
rect 33524 36120 33580 36154
rect 33614 36120 33670 36154
rect 33704 36120 33760 36154
rect 33794 36120 33850 36154
rect 33884 36120 34200 36154
rect 34234 36120 34290 36154
rect 34324 36120 34380 36154
rect 34414 36120 34470 36154
rect 34504 36120 34560 36154
rect 34594 36120 34650 36154
rect 34684 36120 34740 36154
rect 34774 36120 34830 36154
rect 34864 36120 34920 36154
rect 34954 36120 35010 36154
rect 35044 36120 35100 36154
rect 35134 36120 35190 36154
rect 35224 36120 35540 36154
rect 35574 36120 35630 36154
rect 35664 36120 35720 36154
rect 35754 36120 35810 36154
rect 35844 36120 35900 36154
rect 35934 36120 35990 36154
rect 36024 36120 36080 36154
rect 36114 36120 36170 36154
rect 36204 36120 36260 36154
rect 36294 36120 36350 36154
rect 36384 36120 36440 36154
rect 36474 36120 36530 36154
rect 36564 36120 36880 36154
rect 36914 36120 36970 36154
rect 37004 36120 37060 36154
rect 37094 36120 37150 36154
rect 37184 36120 37240 36154
rect 37274 36120 37330 36154
rect 37364 36120 37420 36154
rect 37454 36120 37510 36154
rect 37544 36120 37600 36154
rect 37634 36120 37690 36154
rect 37724 36120 37780 36154
rect 37814 36120 37870 36154
rect 37904 36120 38220 36154
rect 38254 36120 38310 36154
rect 38344 36120 38400 36154
rect 38434 36120 38490 36154
rect 38524 36120 38580 36154
rect 38614 36120 38670 36154
rect 38704 36120 38760 36154
rect 38794 36120 38850 36154
rect 38884 36120 38940 36154
rect 38974 36120 39030 36154
rect 39064 36120 39120 36154
rect 39154 36120 39210 36154
rect 39244 36120 39378 36154
rect 30050 36088 39378 36120
rect 28268 35949 28308 35992
rect 28268 35915 28271 35949
rect 28305 35915 28308 35949
rect 28268 35872 28308 35915
rect 38306 29203 38922 29242
rect 38306 29101 38393 29203
rect 38835 29101 38922 29203
rect 38306 29062 38922 29101
rect 41050 29203 41666 29242
rect 41050 29101 41137 29203
rect 41579 29101 41666 29203
rect 41050 29062 41666 29101
rect 7632 25443 8248 25482
rect 7632 25341 7719 25443
rect 8161 25341 8248 25443
rect 7632 25302 8248 25341
rect 28286 26061 38954 26096
rect 28286 26038 28416 26061
rect 28286 26004 28320 26038
rect 28354 26027 28416 26038
rect 28450 26027 28506 26061
rect 28540 26027 28596 26061
rect 28630 26027 28686 26061
rect 28720 26027 28776 26061
rect 28810 26027 28866 26061
rect 28900 26027 28956 26061
rect 28990 26027 29046 26061
rect 29080 26027 29136 26061
rect 29170 26027 29226 26061
rect 29260 26027 29316 26061
rect 29350 26027 29406 26061
rect 29440 26038 29756 26061
rect 29440 26027 29507 26038
rect 28354 26004 29507 26027
rect 29541 26004 29660 26038
rect 29694 26027 29756 26038
rect 29790 26027 29846 26061
rect 29880 26027 29936 26061
rect 29970 26027 30026 26061
rect 30060 26027 30116 26061
rect 30150 26027 30206 26061
rect 30240 26027 30296 26061
rect 30330 26027 30386 26061
rect 30420 26027 30476 26061
rect 30510 26027 30566 26061
rect 30600 26027 30656 26061
rect 30690 26027 30746 26061
rect 30780 26038 31096 26061
rect 30780 26027 30847 26038
rect 29694 26004 30847 26027
rect 30881 26004 31000 26038
rect 31034 26027 31096 26038
rect 31130 26027 31186 26061
rect 31220 26027 31276 26061
rect 31310 26027 31366 26061
rect 31400 26027 31456 26061
rect 31490 26027 31546 26061
rect 31580 26027 31636 26061
rect 31670 26027 31726 26061
rect 31760 26027 31816 26061
rect 31850 26027 31906 26061
rect 31940 26027 31996 26061
rect 32030 26027 32086 26061
rect 32120 26038 32436 26061
rect 32120 26027 32187 26038
rect 31034 26004 32187 26027
rect 32221 26004 32340 26038
rect 32374 26027 32436 26038
rect 32470 26027 32526 26061
rect 32560 26027 32616 26061
rect 32650 26027 32706 26061
rect 32740 26027 32796 26061
rect 32830 26027 32886 26061
rect 32920 26027 32976 26061
rect 33010 26027 33066 26061
rect 33100 26027 33156 26061
rect 33190 26027 33246 26061
rect 33280 26027 33336 26061
rect 33370 26027 33426 26061
rect 33460 26038 33776 26061
rect 33460 26027 33527 26038
rect 32374 26004 33527 26027
rect 33561 26004 33680 26038
rect 33714 26027 33776 26038
rect 33810 26027 33866 26061
rect 33900 26027 33956 26061
rect 33990 26027 34046 26061
rect 34080 26027 34136 26061
rect 34170 26027 34226 26061
rect 34260 26027 34316 26061
rect 34350 26027 34406 26061
rect 34440 26027 34496 26061
rect 34530 26027 34586 26061
rect 34620 26027 34676 26061
rect 34710 26027 34766 26061
rect 34800 26038 35116 26061
rect 34800 26027 34867 26038
rect 33714 26004 34867 26027
rect 34901 26004 35020 26038
rect 35054 26027 35116 26038
rect 35150 26027 35206 26061
rect 35240 26027 35296 26061
rect 35330 26027 35386 26061
rect 35420 26027 35476 26061
rect 35510 26027 35566 26061
rect 35600 26027 35656 26061
rect 35690 26027 35746 26061
rect 35780 26027 35836 26061
rect 35870 26027 35926 26061
rect 35960 26027 36016 26061
rect 36050 26027 36106 26061
rect 36140 26038 36456 26061
rect 36140 26027 36207 26038
rect 35054 26004 36207 26027
rect 36241 26004 36360 26038
rect 36394 26027 36456 26038
rect 36490 26027 36546 26061
rect 36580 26027 36636 26061
rect 36670 26027 36726 26061
rect 36760 26027 36816 26061
rect 36850 26027 36906 26061
rect 36940 26027 36996 26061
rect 37030 26027 37086 26061
rect 37120 26027 37176 26061
rect 37210 26027 37266 26061
rect 37300 26027 37356 26061
rect 37390 26027 37446 26061
rect 37480 26038 37796 26061
rect 37480 26027 37547 26038
rect 36394 26004 37547 26027
rect 37581 26004 37700 26038
rect 37734 26027 37796 26038
rect 37830 26027 37886 26061
rect 37920 26027 37976 26061
rect 38010 26027 38066 26061
rect 38100 26027 38156 26061
rect 38190 26027 38246 26061
rect 38280 26027 38336 26061
rect 38370 26027 38426 26061
rect 38460 26027 38516 26061
rect 38550 26027 38606 26061
rect 38640 26027 38696 26061
rect 38730 26027 38786 26061
rect 38820 26038 38954 26061
rect 38820 26027 38887 26038
rect 37734 26004 38887 26027
rect 38921 26004 38954 26038
rect 28286 25995 38954 26004
rect 28286 25948 28387 25995
rect 28286 25914 28320 25948
rect 28354 25914 28387 25948
rect 29473 25948 29727 25995
rect 28286 25858 28387 25914
rect 28286 25824 28320 25858
rect 28354 25824 28387 25858
rect 28286 25768 28387 25824
rect 28286 25734 28320 25768
rect 28354 25734 28387 25768
rect 28286 25678 28387 25734
rect 28286 25644 28320 25678
rect 28354 25644 28387 25678
rect 28286 25588 28387 25644
rect 28286 25554 28320 25588
rect 28354 25554 28387 25588
rect 28286 25498 28387 25554
rect 28286 25464 28320 25498
rect 28354 25464 28387 25498
rect 28286 25408 28387 25464
rect 28286 25374 28320 25408
rect 28354 25374 28387 25408
rect 28286 25318 28387 25374
rect 28286 25284 28320 25318
rect 28354 25284 28387 25318
rect 28286 25228 28387 25284
rect 28286 25194 28320 25228
rect 28354 25194 28387 25228
rect 28286 25138 28387 25194
rect 28286 25104 28320 25138
rect 28354 25104 28387 25138
rect 28286 25048 28387 25104
rect 28286 25014 28320 25048
rect 28354 25014 28387 25048
rect 28286 24958 28387 25014
rect 29473 25914 29507 25948
rect 29541 25914 29660 25948
rect 29694 25914 29727 25948
rect 30813 25948 31067 25995
rect 29473 25858 29727 25914
rect 29473 25824 29507 25858
rect 29541 25824 29660 25858
rect 29694 25824 29727 25858
rect 29473 25768 29727 25824
rect 29473 25734 29507 25768
rect 29541 25734 29660 25768
rect 29694 25734 29727 25768
rect 29473 25678 29727 25734
rect 29473 25644 29507 25678
rect 29541 25644 29660 25678
rect 29694 25644 29727 25678
rect 29473 25588 29727 25644
rect 29473 25554 29507 25588
rect 29541 25554 29660 25588
rect 29694 25554 29727 25588
rect 29473 25498 29727 25554
rect 29473 25464 29507 25498
rect 29541 25464 29660 25498
rect 29694 25464 29727 25498
rect 29473 25408 29727 25464
rect 29473 25374 29507 25408
rect 29541 25374 29660 25408
rect 29694 25374 29727 25408
rect 29473 25318 29727 25374
rect 29473 25284 29507 25318
rect 29541 25284 29660 25318
rect 29694 25284 29727 25318
rect 29473 25228 29727 25284
rect 29473 25194 29507 25228
rect 29541 25194 29660 25228
rect 29694 25194 29727 25228
rect 29473 25138 29727 25194
rect 29473 25104 29507 25138
rect 29541 25104 29660 25138
rect 29694 25104 29727 25138
rect 29473 25048 29727 25104
rect 29473 25014 29507 25048
rect 29541 25014 29660 25048
rect 29694 25014 29727 25048
rect 28286 24924 28320 24958
rect 28354 24924 28387 24958
rect 28286 24909 28387 24924
rect 29473 24958 29727 25014
rect 30813 25914 30847 25948
rect 30881 25914 31000 25948
rect 31034 25914 31067 25948
rect 32153 25948 32407 25995
rect 30813 25858 31067 25914
rect 30813 25824 30847 25858
rect 30881 25824 31000 25858
rect 31034 25824 31067 25858
rect 30813 25768 31067 25824
rect 30813 25734 30847 25768
rect 30881 25734 31000 25768
rect 31034 25734 31067 25768
rect 30813 25678 31067 25734
rect 30813 25644 30847 25678
rect 30881 25644 31000 25678
rect 31034 25644 31067 25678
rect 30813 25588 31067 25644
rect 30813 25554 30847 25588
rect 30881 25554 31000 25588
rect 31034 25554 31067 25588
rect 30813 25498 31067 25554
rect 30813 25464 30847 25498
rect 30881 25464 31000 25498
rect 31034 25464 31067 25498
rect 30813 25408 31067 25464
rect 30813 25374 30847 25408
rect 30881 25374 31000 25408
rect 31034 25374 31067 25408
rect 30813 25318 31067 25374
rect 30813 25284 30847 25318
rect 30881 25284 31000 25318
rect 31034 25284 31067 25318
rect 30813 25228 31067 25284
rect 30813 25194 30847 25228
rect 30881 25194 31000 25228
rect 31034 25194 31067 25228
rect 30813 25138 31067 25194
rect 30813 25104 30847 25138
rect 30881 25104 31000 25138
rect 31034 25104 31067 25138
rect 30813 25048 31067 25104
rect 30813 25014 30847 25048
rect 30881 25014 31000 25048
rect 31034 25014 31067 25048
rect 29473 24924 29507 24958
rect 29541 24924 29660 24958
rect 29694 24924 29727 24958
rect 29473 24909 29727 24924
rect 30813 24958 31067 25014
rect 32153 25914 32187 25948
rect 32221 25914 32340 25948
rect 32374 25914 32407 25948
rect 33493 25948 33747 25995
rect 32153 25858 32407 25914
rect 32153 25824 32187 25858
rect 32221 25824 32340 25858
rect 32374 25824 32407 25858
rect 32153 25768 32407 25824
rect 32153 25734 32187 25768
rect 32221 25734 32340 25768
rect 32374 25734 32407 25768
rect 32153 25678 32407 25734
rect 32153 25644 32187 25678
rect 32221 25644 32340 25678
rect 32374 25644 32407 25678
rect 32153 25588 32407 25644
rect 32153 25554 32187 25588
rect 32221 25554 32340 25588
rect 32374 25554 32407 25588
rect 32153 25498 32407 25554
rect 32153 25464 32187 25498
rect 32221 25464 32340 25498
rect 32374 25464 32407 25498
rect 32153 25408 32407 25464
rect 32153 25374 32187 25408
rect 32221 25374 32340 25408
rect 32374 25374 32407 25408
rect 32153 25318 32407 25374
rect 32153 25284 32187 25318
rect 32221 25284 32340 25318
rect 32374 25284 32407 25318
rect 32153 25228 32407 25284
rect 32153 25194 32187 25228
rect 32221 25194 32340 25228
rect 32374 25194 32407 25228
rect 32153 25138 32407 25194
rect 32153 25104 32187 25138
rect 32221 25104 32340 25138
rect 32374 25104 32407 25138
rect 32153 25048 32407 25104
rect 32153 25014 32187 25048
rect 32221 25014 32340 25048
rect 32374 25014 32407 25048
rect 30813 24924 30847 24958
rect 30881 24924 31000 24958
rect 31034 24924 31067 24958
rect 30813 24909 31067 24924
rect 32153 24958 32407 25014
rect 33493 25914 33527 25948
rect 33561 25914 33680 25948
rect 33714 25914 33747 25948
rect 34833 25948 35087 25995
rect 33493 25858 33747 25914
rect 33493 25824 33527 25858
rect 33561 25824 33680 25858
rect 33714 25824 33747 25858
rect 33493 25768 33747 25824
rect 33493 25734 33527 25768
rect 33561 25734 33680 25768
rect 33714 25734 33747 25768
rect 33493 25678 33747 25734
rect 33493 25644 33527 25678
rect 33561 25644 33680 25678
rect 33714 25644 33747 25678
rect 33493 25588 33747 25644
rect 33493 25554 33527 25588
rect 33561 25554 33680 25588
rect 33714 25554 33747 25588
rect 33493 25498 33747 25554
rect 33493 25464 33527 25498
rect 33561 25464 33680 25498
rect 33714 25464 33747 25498
rect 33493 25408 33747 25464
rect 33493 25374 33527 25408
rect 33561 25374 33680 25408
rect 33714 25374 33747 25408
rect 33493 25318 33747 25374
rect 33493 25284 33527 25318
rect 33561 25284 33680 25318
rect 33714 25284 33747 25318
rect 33493 25228 33747 25284
rect 33493 25194 33527 25228
rect 33561 25194 33680 25228
rect 33714 25194 33747 25228
rect 33493 25138 33747 25194
rect 33493 25104 33527 25138
rect 33561 25104 33680 25138
rect 33714 25104 33747 25138
rect 33493 25048 33747 25104
rect 33493 25014 33527 25048
rect 33561 25014 33680 25048
rect 33714 25014 33747 25048
rect 32153 24924 32187 24958
rect 32221 24924 32340 24958
rect 32374 24924 32407 24958
rect 32153 24909 32407 24924
rect 33493 24958 33747 25014
rect 34833 25914 34867 25948
rect 34901 25914 35020 25948
rect 35054 25914 35087 25948
rect 36173 25948 36427 25995
rect 34833 25858 35087 25914
rect 34833 25824 34867 25858
rect 34901 25824 35020 25858
rect 35054 25824 35087 25858
rect 34833 25768 35087 25824
rect 34833 25734 34867 25768
rect 34901 25734 35020 25768
rect 35054 25734 35087 25768
rect 34833 25678 35087 25734
rect 34833 25644 34867 25678
rect 34901 25644 35020 25678
rect 35054 25644 35087 25678
rect 34833 25588 35087 25644
rect 34833 25554 34867 25588
rect 34901 25554 35020 25588
rect 35054 25554 35087 25588
rect 34833 25498 35087 25554
rect 34833 25464 34867 25498
rect 34901 25464 35020 25498
rect 35054 25464 35087 25498
rect 34833 25408 35087 25464
rect 34833 25374 34867 25408
rect 34901 25374 35020 25408
rect 35054 25374 35087 25408
rect 34833 25318 35087 25374
rect 34833 25284 34867 25318
rect 34901 25284 35020 25318
rect 35054 25284 35087 25318
rect 34833 25228 35087 25284
rect 34833 25194 34867 25228
rect 34901 25194 35020 25228
rect 35054 25194 35087 25228
rect 34833 25138 35087 25194
rect 34833 25104 34867 25138
rect 34901 25104 35020 25138
rect 35054 25104 35087 25138
rect 34833 25048 35087 25104
rect 34833 25014 34867 25048
rect 34901 25014 35020 25048
rect 35054 25014 35087 25048
rect 33493 24924 33527 24958
rect 33561 24924 33680 24958
rect 33714 24924 33747 24958
rect 33493 24909 33747 24924
rect 34833 24958 35087 25014
rect 36173 25914 36207 25948
rect 36241 25914 36360 25948
rect 36394 25914 36427 25948
rect 37513 25948 37767 25995
rect 36173 25858 36427 25914
rect 36173 25824 36207 25858
rect 36241 25824 36360 25858
rect 36394 25824 36427 25858
rect 36173 25768 36427 25824
rect 36173 25734 36207 25768
rect 36241 25734 36360 25768
rect 36394 25734 36427 25768
rect 36173 25678 36427 25734
rect 36173 25644 36207 25678
rect 36241 25644 36360 25678
rect 36394 25644 36427 25678
rect 36173 25588 36427 25644
rect 36173 25554 36207 25588
rect 36241 25554 36360 25588
rect 36394 25554 36427 25588
rect 36173 25498 36427 25554
rect 36173 25464 36207 25498
rect 36241 25464 36360 25498
rect 36394 25464 36427 25498
rect 36173 25408 36427 25464
rect 36173 25374 36207 25408
rect 36241 25374 36360 25408
rect 36394 25374 36427 25408
rect 36173 25318 36427 25374
rect 36173 25284 36207 25318
rect 36241 25284 36360 25318
rect 36394 25284 36427 25318
rect 36173 25228 36427 25284
rect 36173 25194 36207 25228
rect 36241 25194 36360 25228
rect 36394 25194 36427 25228
rect 36173 25138 36427 25194
rect 36173 25104 36207 25138
rect 36241 25104 36360 25138
rect 36394 25104 36427 25138
rect 36173 25048 36427 25104
rect 36173 25014 36207 25048
rect 36241 25014 36360 25048
rect 36394 25014 36427 25048
rect 34833 24924 34867 24958
rect 34901 24924 35020 24958
rect 35054 24924 35087 24958
rect 34833 24909 35087 24924
rect 36173 24958 36427 25014
rect 37513 25914 37547 25948
rect 37581 25914 37700 25948
rect 37734 25914 37767 25948
rect 38853 25948 38954 25995
rect 37513 25858 37767 25914
rect 37513 25824 37547 25858
rect 37581 25824 37700 25858
rect 37734 25824 37767 25858
rect 37513 25768 37767 25824
rect 37513 25734 37547 25768
rect 37581 25734 37700 25768
rect 37734 25734 37767 25768
rect 37513 25678 37767 25734
rect 37513 25644 37547 25678
rect 37581 25644 37700 25678
rect 37734 25644 37767 25678
rect 37513 25588 37767 25644
rect 37513 25554 37547 25588
rect 37581 25554 37700 25588
rect 37734 25554 37767 25588
rect 37513 25498 37767 25554
rect 37513 25464 37547 25498
rect 37581 25464 37700 25498
rect 37734 25464 37767 25498
rect 37513 25408 37767 25464
rect 37513 25374 37547 25408
rect 37581 25374 37700 25408
rect 37734 25374 37767 25408
rect 37513 25318 37767 25374
rect 37513 25284 37547 25318
rect 37581 25284 37700 25318
rect 37734 25284 37767 25318
rect 37513 25228 37767 25284
rect 37513 25194 37547 25228
rect 37581 25194 37700 25228
rect 37734 25194 37767 25228
rect 37513 25138 37767 25194
rect 37513 25104 37547 25138
rect 37581 25104 37700 25138
rect 37734 25104 37767 25138
rect 37513 25048 37767 25104
rect 37513 25014 37547 25048
rect 37581 25014 37700 25048
rect 37734 25014 37767 25048
rect 36173 24924 36207 24958
rect 36241 24924 36360 24958
rect 36394 24924 36427 24958
rect 36173 24909 36427 24924
rect 37513 24958 37767 25014
rect 38853 25914 38887 25948
rect 38921 25914 38954 25948
rect 38853 25858 38954 25914
rect 38853 25824 38887 25858
rect 38921 25824 38954 25858
rect 38853 25768 38954 25824
rect 38853 25734 38887 25768
rect 38921 25734 38954 25768
rect 38853 25678 38954 25734
rect 38853 25644 38887 25678
rect 38921 25644 38954 25678
rect 38853 25588 38954 25644
rect 38853 25554 38887 25588
rect 38921 25554 38954 25588
rect 38853 25498 38954 25554
rect 38853 25464 38887 25498
rect 38921 25464 38954 25498
rect 38853 25408 38954 25464
rect 38853 25374 38887 25408
rect 38921 25374 38954 25408
rect 38853 25318 38954 25374
rect 38853 25284 38887 25318
rect 38921 25284 38954 25318
rect 40658 25443 41274 25482
rect 40658 25341 40745 25443
rect 41187 25341 41274 25443
rect 40658 25302 41274 25341
rect 38853 25228 38954 25284
rect 38853 25194 38887 25228
rect 38921 25194 38954 25228
rect 38853 25138 38954 25194
rect 38853 25104 38887 25138
rect 38921 25104 38954 25138
rect 38853 25048 38954 25104
rect 38853 25014 38887 25048
rect 38921 25014 38954 25048
rect 37513 24924 37547 24958
rect 37581 24924 37700 24958
rect 37734 24924 37767 24958
rect 37513 24909 37767 24924
rect 38853 24958 38954 25014
rect 38853 24924 38887 24958
rect 38921 24924 38954 24958
rect 38853 24909 38954 24924
rect 28286 24874 38954 24909
rect 28286 24840 28416 24874
rect 28450 24840 28506 24874
rect 28540 24840 28596 24874
rect 28630 24840 28686 24874
rect 28720 24840 28776 24874
rect 28810 24840 28866 24874
rect 28900 24840 28956 24874
rect 28990 24840 29046 24874
rect 29080 24840 29136 24874
rect 29170 24840 29226 24874
rect 29260 24840 29316 24874
rect 29350 24840 29406 24874
rect 29440 24840 29756 24874
rect 29790 24840 29846 24874
rect 29880 24840 29936 24874
rect 29970 24840 30026 24874
rect 30060 24840 30116 24874
rect 30150 24840 30206 24874
rect 30240 24840 30296 24874
rect 30330 24840 30386 24874
rect 30420 24840 30476 24874
rect 30510 24840 30566 24874
rect 30600 24840 30656 24874
rect 30690 24840 30746 24874
rect 30780 24840 31096 24874
rect 31130 24840 31186 24874
rect 31220 24840 31276 24874
rect 31310 24840 31366 24874
rect 31400 24840 31456 24874
rect 31490 24840 31546 24874
rect 31580 24840 31636 24874
rect 31670 24840 31726 24874
rect 31760 24840 31816 24874
rect 31850 24840 31906 24874
rect 31940 24840 31996 24874
rect 32030 24840 32086 24874
rect 32120 24840 32436 24874
rect 32470 24840 32526 24874
rect 32560 24840 32616 24874
rect 32650 24840 32706 24874
rect 32740 24840 32796 24874
rect 32830 24840 32886 24874
rect 32920 24840 32976 24874
rect 33010 24840 33066 24874
rect 33100 24840 33156 24874
rect 33190 24840 33246 24874
rect 33280 24840 33336 24874
rect 33370 24840 33426 24874
rect 33460 24840 33776 24874
rect 33810 24840 33866 24874
rect 33900 24840 33956 24874
rect 33990 24840 34046 24874
rect 34080 24840 34136 24874
rect 34170 24840 34226 24874
rect 34260 24840 34316 24874
rect 34350 24840 34406 24874
rect 34440 24840 34496 24874
rect 34530 24840 34586 24874
rect 34620 24840 34676 24874
rect 34710 24840 34766 24874
rect 34800 24840 35116 24874
rect 35150 24840 35206 24874
rect 35240 24840 35296 24874
rect 35330 24840 35386 24874
rect 35420 24840 35476 24874
rect 35510 24840 35566 24874
rect 35600 24840 35656 24874
rect 35690 24840 35746 24874
rect 35780 24840 35836 24874
rect 35870 24840 35926 24874
rect 35960 24840 36016 24874
rect 36050 24840 36106 24874
rect 36140 24840 36456 24874
rect 36490 24840 36546 24874
rect 36580 24840 36636 24874
rect 36670 24840 36726 24874
rect 36760 24840 36816 24874
rect 36850 24840 36906 24874
rect 36940 24840 36996 24874
rect 37030 24840 37086 24874
rect 37120 24840 37176 24874
rect 37210 24840 37266 24874
rect 37300 24840 37356 24874
rect 37390 24840 37446 24874
rect 37480 24840 37796 24874
rect 37830 24840 37886 24874
rect 37920 24840 37976 24874
rect 38010 24840 38066 24874
rect 38100 24840 38156 24874
rect 38190 24840 38246 24874
rect 38280 24840 38336 24874
rect 38370 24840 38426 24874
rect 38460 24840 38516 24874
rect 38550 24840 38606 24874
rect 38640 24840 38696 24874
rect 38730 24840 38786 24874
rect 38820 24840 38954 24874
rect 28286 24808 38954 24840
rect 22908 24669 22948 24712
rect 22908 24635 22911 24669
rect 22945 24635 22948 24669
rect 22908 24592 22948 24635
rect 23968 24639 24088 24642
rect 23968 24605 24013 24639
rect 24047 24605 24088 24639
rect 23968 24592 24088 24605
rect 25268 24639 25388 24642
rect 25268 24605 25313 24639
rect 25347 24605 25388 24639
rect 25268 24592 25388 24605
rect 21034 22301 22322 22336
rect 21034 22278 21164 22301
rect 21034 22244 21068 22278
rect 21102 22267 21164 22278
rect 21198 22267 21254 22301
rect 21288 22267 21344 22301
rect 21378 22267 21434 22301
rect 21468 22267 21524 22301
rect 21558 22267 21614 22301
rect 21648 22267 21704 22301
rect 21738 22267 21794 22301
rect 21828 22267 21884 22301
rect 21918 22267 21974 22301
rect 22008 22267 22064 22301
rect 22098 22267 22154 22301
rect 22188 22278 22322 22301
rect 22188 22267 22255 22278
rect 21102 22244 22255 22267
rect 22289 22244 22322 22278
rect 21034 22235 22322 22244
rect 21034 22188 21135 22235
rect 21034 22154 21068 22188
rect 21102 22154 21135 22188
rect 22221 22188 22322 22235
rect 21034 22098 21135 22154
rect 21034 22064 21068 22098
rect 21102 22064 21135 22098
rect 21034 22008 21135 22064
rect 21034 21974 21068 22008
rect 21102 21974 21135 22008
rect 21034 21918 21135 21974
rect 21034 21884 21068 21918
rect 21102 21884 21135 21918
rect 21034 21828 21135 21884
rect 21034 21794 21068 21828
rect 21102 21794 21135 21828
rect 21034 21738 21135 21794
rect 21034 21704 21068 21738
rect 21102 21704 21135 21738
rect 21034 21648 21135 21704
rect 21034 21614 21068 21648
rect 21102 21614 21135 21648
rect 21034 21558 21135 21614
rect 21034 21524 21068 21558
rect 21102 21524 21135 21558
rect 21034 21468 21135 21524
rect 21034 21434 21068 21468
rect 21102 21434 21135 21468
rect 21034 21378 21135 21434
rect 21034 21344 21068 21378
rect 21102 21344 21135 21378
rect 21034 21288 21135 21344
rect 21034 21254 21068 21288
rect 21102 21254 21135 21288
rect 21034 21198 21135 21254
rect 22221 22154 22255 22188
rect 22289 22154 22322 22188
rect 28286 22301 38954 22336
rect 28286 22278 28416 22301
rect 28286 22244 28320 22278
rect 28354 22267 28416 22278
rect 28450 22267 28506 22301
rect 28540 22267 28596 22301
rect 28630 22267 28686 22301
rect 28720 22267 28776 22301
rect 28810 22267 28866 22301
rect 28900 22267 28956 22301
rect 28990 22267 29046 22301
rect 29080 22267 29136 22301
rect 29170 22267 29226 22301
rect 29260 22267 29316 22301
rect 29350 22267 29406 22301
rect 29440 22278 29756 22301
rect 29440 22267 29507 22278
rect 28354 22244 29507 22267
rect 29541 22244 29660 22278
rect 29694 22267 29756 22278
rect 29790 22267 29846 22301
rect 29880 22267 29936 22301
rect 29970 22267 30026 22301
rect 30060 22267 30116 22301
rect 30150 22267 30206 22301
rect 30240 22267 30296 22301
rect 30330 22267 30386 22301
rect 30420 22267 30476 22301
rect 30510 22267 30566 22301
rect 30600 22267 30656 22301
rect 30690 22267 30746 22301
rect 30780 22278 31096 22301
rect 30780 22267 30847 22278
rect 29694 22244 30847 22267
rect 30881 22244 31000 22278
rect 31034 22267 31096 22278
rect 31130 22267 31186 22301
rect 31220 22267 31276 22301
rect 31310 22267 31366 22301
rect 31400 22267 31456 22301
rect 31490 22267 31546 22301
rect 31580 22267 31636 22301
rect 31670 22267 31726 22301
rect 31760 22267 31816 22301
rect 31850 22267 31906 22301
rect 31940 22267 31996 22301
rect 32030 22267 32086 22301
rect 32120 22278 32436 22301
rect 32120 22267 32187 22278
rect 31034 22244 32187 22267
rect 32221 22244 32340 22278
rect 32374 22267 32436 22278
rect 32470 22267 32526 22301
rect 32560 22267 32616 22301
rect 32650 22267 32706 22301
rect 32740 22267 32796 22301
rect 32830 22267 32886 22301
rect 32920 22267 32976 22301
rect 33010 22267 33066 22301
rect 33100 22267 33156 22301
rect 33190 22267 33246 22301
rect 33280 22267 33336 22301
rect 33370 22267 33426 22301
rect 33460 22278 33776 22301
rect 33460 22267 33527 22278
rect 32374 22244 33527 22267
rect 33561 22244 33680 22278
rect 33714 22267 33776 22278
rect 33810 22267 33866 22301
rect 33900 22267 33956 22301
rect 33990 22267 34046 22301
rect 34080 22267 34136 22301
rect 34170 22267 34226 22301
rect 34260 22267 34316 22301
rect 34350 22267 34406 22301
rect 34440 22267 34496 22301
rect 34530 22267 34586 22301
rect 34620 22267 34676 22301
rect 34710 22267 34766 22301
rect 34800 22278 35116 22301
rect 34800 22267 34867 22278
rect 33714 22244 34867 22267
rect 34901 22244 35020 22278
rect 35054 22267 35116 22278
rect 35150 22267 35206 22301
rect 35240 22267 35296 22301
rect 35330 22267 35386 22301
rect 35420 22267 35476 22301
rect 35510 22267 35566 22301
rect 35600 22267 35656 22301
rect 35690 22267 35746 22301
rect 35780 22267 35836 22301
rect 35870 22267 35926 22301
rect 35960 22267 36016 22301
rect 36050 22267 36106 22301
rect 36140 22278 36456 22301
rect 36140 22267 36207 22278
rect 35054 22244 36207 22267
rect 36241 22244 36360 22278
rect 36394 22267 36456 22278
rect 36490 22267 36546 22301
rect 36580 22267 36636 22301
rect 36670 22267 36726 22301
rect 36760 22267 36816 22301
rect 36850 22267 36906 22301
rect 36940 22267 36996 22301
rect 37030 22267 37086 22301
rect 37120 22267 37176 22301
rect 37210 22267 37266 22301
rect 37300 22267 37356 22301
rect 37390 22267 37446 22301
rect 37480 22278 37796 22301
rect 37480 22267 37547 22278
rect 36394 22244 37547 22267
rect 37581 22244 37700 22278
rect 37734 22267 37796 22278
rect 37830 22267 37886 22301
rect 37920 22267 37976 22301
rect 38010 22267 38066 22301
rect 38100 22267 38156 22301
rect 38190 22267 38246 22301
rect 38280 22267 38336 22301
rect 38370 22267 38426 22301
rect 38460 22267 38516 22301
rect 38550 22267 38606 22301
rect 38640 22267 38696 22301
rect 38730 22267 38786 22301
rect 38820 22278 38954 22301
rect 38820 22267 38887 22278
rect 37734 22244 38887 22267
rect 38921 22244 38954 22278
rect 28286 22235 38954 22244
rect 28286 22188 28387 22235
rect 22221 22098 22322 22154
rect 28286 22154 28320 22188
rect 28354 22154 28387 22188
rect 29473 22188 29727 22235
rect 22221 22064 22255 22098
rect 22289 22064 22322 22098
rect 22221 22008 22322 22064
rect 22221 21974 22255 22008
rect 22289 21974 22322 22008
rect 22221 21918 22322 21974
rect 22221 21884 22255 21918
rect 22289 21884 22322 21918
rect 22221 21828 22322 21884
rect 22221 21794 22255 21828
rect 22289 21794 22322 21828
rect 22221 21738 22322 21794
rect 22221 21704 22255 21738
rect 22289 21704 22322 21738
rect 22221 21648 22322 21704
rect 22221 21614 22255 21648
rect 22289 21614 22322 21648
rect 22221 21558 22322 21614
rect 22221 21524 22255 21558
rect 22289 21524 22322 21558
rect 22221 21468 22322 21524
rect 22221 21434 22255 21468
rect 22289 21434 22322 21468
rect 22221 21378 22322 21434
rect 22221 21344 22255 21378
rect 22289 21344 22322 21378
rect 28286 22098 28387 22154
rect 28286 22064 28320 22098
rect 28354 22064 28387 22098
rect 28286 22008 28387 22064
rect 28286 21974 28320 22008
rect 28354 21974 28387 22008
rect 28286 21918 28387 21974
rect 28286 21884 28320 21918
rect 28354 21884 28387 21918
rect 28286 21828 28387 21884
rect 28286 21794 28320 21828
rect 28354 21794 28387 21828
rect 28286 21738 28387 21794
rect 28286 21704 28320 21738
rect 28354 21704 28387 21738
rect 28286 21648 28387 21704
rect 28286 21614 28320 21648
rect 28354 21614 28387 21648
rect 28286 21558 28387 21614
rect 28286 21524 28320 21558
rect 28354 21524 28387 21558
rect 28286 21468 28387 21524
rect 28286 21434 28320 21468
rect 28354 21434 28387 21468
rect 28286 21378 28387 21434
rect 22221 21288 22322 21344
rect 28286 21344 28320 21378
rect 28354 21344 28387 21378
rect 22221 21254 22255 21288
rect 22289 21254 22322 21288
rect 21034 21164 21068 21198
rect 21102 21164 21135 21198
rect 21034 21149 21135 21164
rect 22221 21198 22322 21254
rect 22221 21164 22255 21198
rect 22289 21164 22322 21198
rect 22221 21149 22322 21164
rect 21034 21114 22322 21149
rect 28286 21288 28387 21344
rect 28286 21254 28320 21288
rect 28354 21254 28387 21288
rect 28286 21198 28387 21254
rect 29473 22154 29507 22188
rect 29541 22154 29660 22188
rect 29694 22154 29727 22188
rect 30813 22188 31067 22235
rect 29473 22098 29727 22154
rect 29473 22064 29507 22098
rect 29541 22064 29660 22098
rect 29694 22064 29727 22098
rect 29473 22008 29727 22064
rect 29473 21974 29507 22008
rect 29541 21974 29660 22008
rect 29694 21974 29727 22008
rect 29473 21918 29727 21974
rect 29473 21884 29507 21918
rect 29541 21884 29660 21918
rect 29694 21884 29727 21918
rect 29473 21828 29727 21884
rect 29473 21794 29507 21828
rect 29541 21794 29660 21828
rect 29694 21794 29727 21828
rect 29473 21738 29727 21794
rect 29473 21704 29507 21738
rect 29541 21704 29660 21738
rect 29694 21704 29727 21738
rect 29473 21648 29727 21704
rect 29473 21614 29507 21648
rect 29541 21614 29660 21648
rect 29694 21614 29727 21648
rect 29473 21558 29727 21614
rect 29473 21524 29507 21558
rect 29541 21524 29660 21558
rect 29694 21524 29727 21558
rect 29473 21468 29727 21524
rect 29473 21434 29507 21468
rect 29541 21434 29660 21468
rect 29694 21434 29727 21468
rect 29473 21378 29727 21434
rect 29473 21344 29507 21378
rect 29541 21344 29660 21378
rect 29694 21344 29727 21378
rect 29473 21288 29727 21344
rect 29473 21254 29507 21288
rect 29541 21254 29660 21288
rect 29694 21254 29727 21288
rect 28286 21164 28320 21198
rect 28354 21164 28387 21198
rect 28286 21149 28387 21164
rect 29473 21198 29727 21254
rect 30813 22154 30847 22188
rect 30881 22154 31000 22188
rect 31034 22154 31067 22188
rect 32153 22188 32407 22235
rect 30813 22098 31067 22154
rect 30813 22064 30847 22098
rect 30881 22064 31000 22098
rect 31034 22064 31067 22098
rect 30813 22008 31067 22064
rect 30813 21974 30847 22008
rect 30881 21974 31000 22008
rect 31034 21974 31067 22008
rect 30813 21918 31067 21974
rect 30813 21884 30847 21918
rect 30881 21884 31000 21918
rect 31034 21884 31067 21918
rect 30813 21828 31067 21884
rect 30813 21794 30847 21828
rect 30881 21794 31000 21828
rect 31034 21794 31067 21828
rect 30813 21738 31067 21794
rect 30813 21704 30847 21738
rect 30881 21704 31000 21738
rect 31034 21704 31067 21738
rect 30813 21648 31067 21704
rect 30813 21614 30847 21648
rect 30881 21614 31000 21648
rect 31034 21614 31067 21648
rect 30813 21558 31067 21614
rect 30813 21524 30847 21558
rect 30881 21524 31000 21558
rect 31034 21524 31067 21558
rect 30813 21468 31067 21524
rect 30813 21434 30847 21468
rect 30881 21434 31000 21468
rect 31034 21434 31067 21468
rect 30813 21378 31067 21434
rect 30813 21344 30847 21378
rect 30881 21344 31000 21378
rect 31034 21344 31067 21378
rect 30813 21288 31067 21344
rect 30813 21254 30847 21288
rect 30881 21254 31000 21288
rect 31034 21254 31067 21288
rect 29473 21164 29507 21198
rect 29541 21164 29660 21198
rect 29694 21164 29727 21198
rect 29473 21149 29727 21164
rect 30813 21198 31067 21254
rect 32153 22154 32187 22188
rect 32221 22154 32340 22188
rect 32374 22154 32407 22188
rect 33493 22188 33747 22235
rect 32153 22098 32407 22154
rect 32153 22064 32187 22098
rect 32221 22064 32340 22098
rect 32374 22064 32407 22098
rect 32153 22008 32407 22064
rect 32153 21974 32187 22008
rect 32221 21974 32340 22008
rect 32374 21974 32407 22008
rect 32153 21918 32407 21974
rect 32153 21884 32187 21918
rect 32221 21884 32340 21918
rect 32374 21884 32407 21918
rect 32153 21828 32407 21884
rect 32153 21794 32187 21828
rect 32221 21794 32340 21828
rect 32374 21794 32407 21828
rect 32153 21738 32407 21794
rect 32153 21704 32187 21738
rect 32221 21704 32340 21738
rect 32374 21704 32407 21738
rect 32153 21648 32407 21704
rect 32153 21614 32187 21648
rect 32221 21614 32340 21648
rect 32374 21614 32407 21648
rect 32153 21558 32407 21614
rect 32153 21524 32187 21558
rect 32221 21524 32340 21558
rect 32374 21524 32407 21558
rect 32153 21468 32407 21524
rect 32153 21434 32187 21468
rect 32221 21434 32340 21468
rect 32374 21434 32407 21468
rect 32153 21378 32407 21434
rect 32153 21344 32187 21378
rect 32221 21344 32340 21378
rect 32374 21344 32407 21378
rect 32153 21288 32407 21344
rect 32153 21254 32187 21288
rect 32221 21254 32340 21288
rect 32374 21254 32407 21288
rect 30813 21164 30847 21198
rect 30881 21164 31000 21198
rect 31034 21164 31067 21198
rect 30813 21149 31067 21164
rect 32153 21198 32407 21254
rect 33493 22154 33527 22188
rect 33561 22154 33680 22188
rect 33714 22154 33747 22188
rect 34833 22188 35087 22235
rect 33493 22098 33747 22154
rect 33493 22064 33527 22098
rect 33561 22064 33680 22098
rect 33714 22064 33747 22098
rect 33493 22008 33747 22064
rect 33493 21974 33527 22008
rect 33561 21974 33680 22008
rect 33714 21974 33747 22008
rect 33493 21918 33747 21974
rect 33493 21884 33527 21918
rect 33561 21884 33680 21918
rect 33714 21884 33747 21918
rect 33493 21828 33747 21884
rect 33493 21794 33527 21828
rect 33561 21794 33680 21828
rect 33714 21794 33747 21828
rect 33493 21738 33747 21794
rect 33493 21704 33527 21738
rect 33561 21704 33680 21738
rect 33714 21704 33747 21738
rect 33493 21648 33747 21704
rect 33493 21614 33527 21648
rect 33561 21614 33680 21648
rect 33714 21614 33747 21648
rect 33493 21558 33747 21614
rect 33493 21524 33527 21558
rect 33561 21524 33680 21558
rect 33714 21524 33747 21558
rect 33493 21468 33747 21524
rect 33493 21434 33527 21468
rect 33561 21434 33680 21468
rect 33714 21434 33747 21468
rect 33493 21378 33747 21434
rect 33493 21344 33527 21378
rect 33561 21344 33680 21378
rect 33714 21344 33747 21378
rect 33493 21288 33747 21344
rect 33493 21254 33527 21288
rect 33561 21254 33680 21288
rect 33714 21254 33747 21288
rect 32153 21164 32187 21198
rect 32221 21164 32340 21198
rect 32374 21164 32407 21198
rect 32153 21149 32407 21164
rect 33493 21198 33747 21254
rect 34833 22154 34867 22188
rect 34901 22154 35020 22188
rect 35054 22154 35087 22188
rect 36173 22188 36427 22235
rect 34833 22098 35087 22154
rect 34833 22064 34867 22098
rect 34901 22064 35020 22098
rect 35054 22064 35087 22098
rect 34833 22008 35087 22064
rect 34833 21974 34867 22008
rect 34901 21974 35020 22008
rect 35054 21974 35087 22008
rect 34833 21918 35087 21974
rect 34833 21884 34867 21918
rect 34901 21884 35020 21918
rect 35054 21884 35087 21918
rect 34833 21828 35087 21884
rect 34833 21794 34867 21828
rect 34901 21794 35020 21828
rect 35054 21794 35087 21828
rect 34833 21738 35087 21794
rect 34833 21704 34867 21738
rect 34901 21704 35020 21738
rect 35054 21704 35087 21738
rect 34833 21648 35087 21704
rect 34833 21614 34867 21648
rect 34901 21614 35020 21648
rect 35054 21614 35087 21648
rect 34833 21558 35087 21614
rect 34833 21524 34867 21558
rect 34901 21524 35020 21558
rect 35054 21524 35087 21558
rect 34833 21468 35087 21524
rect 34833 21434 34867 21468
rect 34901 21434 35020 21468
rect 35054 21434 35087 21468
rect 34833 21378 35087 21434
rect 34833 21344 34867 21378
rect 34901 21344 35020 21378
rect 35054 21344 35087 21378
rect 34833 21288 35087 21344
rect 34833 21254 34867 21288
rect 34901 21254 35020 21288
rect 35054 21254 35087 21288
rect 33493 21164 33527 21198
rect 33561 21164 33680 21198
rect 33714 21164 33747 21198
rect 33493 21149 33747 21164
rect 34833 21198 35087 21254
rect 36173 22154 36207 22188
rect 36241 22154 36360 22188
rect 36394 22154 36427 22188
rect 37513 22188 37767 22235
rect 36173 22098 36427 22154
rect 36173 22064 36207 22098
rect 36241 22064 36360 22098
rect 36394 22064 36427 22098
rect 36173 22008 36427 22064
rect 36173 21974 36207 22008
rect 36241 21974 36360 22008
rect 36394 21974 36427 22008
rect 36173 21918 36427 21974
rect 36173 21884 36207 21918
rect 36241 21884 36360 21918
rect 36394 21884 36427 21918
rect 36173 21828 36427 21884
rect 36173 21794 36207 21828
rect 36241 21794 36360 21828
rect 36394 21794 36427 21828
rect 36173 21738 36427 21794
rect 36173 21704 36207 21738
rect 36241 21704 36360 21738
rect 36394 21704 36427 21738
rect 36173 21648 36427 21704
rect 36173 21614 36207 21648
rect 36241 21614 36360 21648
rect 36394 21614 36427 21648
rect 36173 21558 36427 21614
rect 36173 21524 36207 21558
rect 36241 21524 36360 21558
rect 36394 21524 36427 21558
rect 36173 21468 36427 21524
rect 36173 21434 36207 21468
rect 36241 21434 36360 21468
rect 36394 21434 36427 21468
rect 36173 21378 36427 21434
rect 36173 21344 36207 21378
rect 36241 21344 36360 21378
rect 36394 21344 36427 21378
rect 36173 21288 36427 21344
rect 36173 21254 36207 21288
rect 36241 21254 36360 21288
rect 36394 21254 36427 21288
rect 34833 21164 34867 21198
rect 34901 21164 35020 21198
rect 35054 21164 35087 21198
rect 34833 21149 35087 21164
rect 36173 21198 36427 21254
rect 37513 22154 37547 22188
rect 37581 22154 37700 22188
rect 37734 22154 37767 22188
rect 38853 22188 38954 22235
rect 37513 22098 37767 22154
rect 37513 22064 37547 22098
rect 37581 22064 37700 22098
rect 37734 22064 37767 22098
rect 37513 22008 37767 22064
rect 37513 21974 37547 22008
rect 37581 21974 37700 22008
rect 37734 21974 37767 22008
rect 37513 21918 37767 21974
rect 37513 21884 37547 21918
rect 37581 21884 37700 21918
rect 37734 21884 37767 21918
rect 37513 21828 37767 21884
rect 37513 21794 37547 21828
rect 37581 21794 37700 21828
rect 37734 21794 37767 21828
rect 37513 21738 37767 21794
rect 37513 21704 37547 21738
rect 37581 21704 37700 21738
rect 37734 21704 37767 21738
rect 37513 21648 37767 21704
rect 37513 21614 37547 21648
rect 37581 21614 37700 21648
rect 37734 21614 37767 21648
rect 37513 21558 37767 21614
rect 37513 21524 37547 21558
rect 37581 21524 37700 21558
rect 37734 21524 37767 21558
rect 37513 21468 37767 21524
rect 37513 21434 37547 21468
rect 37581 21434 37700 21468
rect 37734 21434 37767 21468
rect 37513 21378 37767 21434
rect 37513 21344 37547 21378
rect 37581 21344 37700 21378
rect 37734 21344 37767 21378
rect 37513 21288 37767 21344
rect 37513 21254 37547 21288
rect 37581 21254 37700 21288
rect 37734 21254 37767 21288
rect 36173 21164 36207 21198
rect 36241 21164 36360 21198
rect 36394 21164 36427 21198
rect 36173 21149 36427 21164
rect 37513 21198 37767 21254
rect 38853 22154 38887 22188
rect 38921 22154 38954 22188
rect 38853 22098 38954 22154
rect 38853 22064 38887 22098
rect 38921 22064 38954 22098
rect 38853 22008 38954 22064
rect 38853 21974 38887 22008
rect 38921 21974 38954 22008
rect 38853 21918 38954 21974
rect 38853 21884 38887 21918
rect 38921 21884 38954 21918
rect 38853 21828 38954 21884
rect 38853 21794 38887 21828
rect 38921 21794 38954 21828
rect 38853 21738 38954 21794
rect 38853 21704 38887 21738
rect 38921 21704 38954 21738
rect 38853 21648 38954 21704
rect 38853 21614 38887 21648
rect 38921 21614 38954 21648
rect 38853 21558 38954 21614
rect 38853 21524 38887 21558
rect 38921 21524 38954 21558
rect 40658 21683 41274 21722
rect 40658 21581 40745 21683
rect 41187 21581 41274 21683
rect 40658 21542 41274 21581
rect 38853 21468 38954 21524
rect 38853 21434 38887 21468
rect 38921 21434 38954 21468
rect 38853 21378 38954 21434
rect 38853 21344 38887 21378
rect 38921 21344 38954 21378
rect 38853 21288 38954 21344
rect 38853 21254 38887 21288
rect 38921 21254 38954 21288
rect 37513 21164 37547 21198
rect 37581 21164 37700 21198
rect 37734 21164 37767 21198
rect 37513 21149 37767 21164
rect 38853 21198 38954 21254
rect 38853 21164 38887 21198
rect 38921 21164 38954 21198
rect 38853 21149 38954 21164
rect 21034 21080 21164 21114
rect 21198 21080 21254 21114
rect 21288 21080 21344 21114
rect 21378 21080 21434 21114
rect 21468 21080 21524 21114
rect 21558 21080 21614 21114
rect 21648 21080 21704 21114
rect 21738 21080 21794 21114
rect 21828 21080 21884 21114
rect 21918 21080 21974 21114
rect 22008 21080 22064 21114
rect 22098 21080 22154 21114
rect 22188 21080 22322 21114
rect 21034 21048 22322 21080
rect 28286 21114 38954 21149
rect 28286 21080 28416 21114
rect 28450 21080 28506 21114
rect 28540 21080 28596 21114
rect 28630 21080 28686 21114
rect 28720 21080 28776 21114
rect 28810 21080 28866 21114
rect 28900 21080 28956 21114
rect 28990 21080 29046 21114
rect 29080 21080 29136 21114
rect 29170 21080 29226 21114
rect 29260 21080 29316 21114
rect 29350 21080 29406 21114
rect 29440 21080 29756 21114
rect 29790 21080 29846 21114
rect 29880 21080 29936 21114
rect 29970 21080 30026 21114
rect 30060 21080 30116 21114
rect 30150 21080 30206 21114
rect 30240 21080 30296 21114
rect 30330 21080 30386 21114
rect 30420 21080 30476 21114
rect 30510 21080 30566 21114
rect 30600 21080 30656 21114
rect 30690 21080 30746 21114
rect 30780 21080 31096 21114
rect 31130 21080 31186 21114
rect 31220 21080 31276 21114
rect 31310 21080 31366 21114
rect 31400 21080 31456 21114
rect 31490 21080 31546 21114
rect 31580 21080 31636 21114
rect 31670 21080 31726 21114
rect 31760 21080 31816 21114
rect 31850 21080 31906 21114
rect 31940 21080 31996 21114
rect 32030 21080 32086 21114
rect 32120 21080 32436 21114
rect 32470 21080 32526 21114
rect 32560 21080 32616 21114
rect 32650 21080 32706 21114
rect 32740 21080 32796 21114
rect 32830 21080 32886 21114
rect 32920 21080 32976 21114
rect 33010 21080 33066 21114
rect 33100 21080 33156 21114
rect 33190 21080 33246 21114
rect 33280 21080 33336 21114
rect 33370 21080 33426 21114
rect 33460 21080 33776 21114
rect 33810 21080 33866 21114
rect 33900 21080 33956 21114
rect 33990 21080 34046 21114
rect 34080 21080 34136 21114
rect 34170 21080 34226 21114
rect 34260 21080 34316 21114
rect 34350 21080 34406 21114
rect 34440 21080 34496 21114
rect 34530 21080 34586 21114
rect 34620 21080 34676 21114
rect 34710 21080 34766 21114
rect 34800 21080 35116 21114
rect 35150 21080 35206 21114
rect 35240 21080 35296 21114
rect 35330 21080 35386 21114
rect 35420 21080 35476 21114
rect 35510 21080 35566 21114
rect 35600 21080 35656 21114
rect 35690 21080 35746 21114
rect 35780 21080 35836 21114
rect 35870 21080 35926 21114
rect 35960 21080 36016 21114
rect 36050 21080 36106 21114
rect 36140 21080 36456 21114
rect 36490 21080 36546 21114
rect 36580 21080 36636 21114
rect 36670 21080 36726 21114
rect 36760 21080 36816 21114
rect 36850 21080 36906 21114
rect 36940 21080 36996 21114
rect 37030 21080 37086 21114
rect 37120 21080 37176 21114
rect 37210 21080 37266 21114
rect 37300 21080 37356 21114
rect 37390 21080 37446 21114
rect 37480 21080 37796 21114
rect 37830 21080 37886 21114
rect 37920 21080 37976 21114
rect 38010 21080 38066 21114
rect 38100 21080 38156 21114
rect 38190 21080 38246 21114
rect 38280 21080 38336 21114
rect 38370 21080 38426 21114
rect 38460 21080 38516 21114
rect 38550 21080 38606 21114
rect 38640 21080 38696 21114
rect 38730 21080 38786 21114
rect 38820 21080 38954 21114
rect 28286 21048 38954 21080
rect 22908 20909 22948 20952
rect 22908 20875 22911 20909
rect 22945 20875 22948 20909
rect 22908 20832 22948 20875
rect 23968 20879 24088 20882
rect 23968 20845 24013 20879
rect 24047 20845 24088 20879
rect 23968 20832 24088 20845
rect 25268 20879 25388 20882
rect 25268 20845 25313 20879
rect 25347 20845 25388 20879
rect 25268 20832 25388 20845
rect 11552 17923 12168 17962
rect 11552 17821 11639 17923
rect 12081 17821 12168 17923
rect 11552 17782 12168 17821
rect 14296 17923 14912 17962
rect 14296 17821 14383 17923
rect 14825 17821 14912 17923
rect 14296 17782 14912 17821
rect 5954 17149 5994 17192
rect 5954 17115 5957 17149
rect 5991 17115 5994 17149
rect 5954 17072 5994 17115
rect 7014 17119 7134 17122
rect 7014 17085 7059 17119
rect 7093 17085 7134 17119
rect 7014 17072 7134 17085
rect 8314 17119 8434 17122
rect 8314 17085 8359 17119
rect 8393 17085 8434 17119
rect 28286 18541 38954 18576
rect 28286 18518 28416 18541
rect 28286 18484 28320 18518
rect 28354 18507 28416 18518
rect 28450 18507 28506 18541
rect 28540 18507 28596 18541
rect 28630 18507 28686 18541
rect 28720 18507 28776 18541
rect 28810 18507 28866 18541
rect 28900 18507 28956 18541
rect 28990 18507 29046 18541
rect 29080 18507 29136 18541
rect 29170 18507 29226 18541
rect 29260 18507 29316 18541
rect 29350 18507 29406 18541
rect 29440 18518 29756 18541
rect 29440 18507 29507 18518
rect 28354 18484 29507 18507
rect 29541 18484 29660 18518
rect 29694 18507 29756 18518
rect 29790 18507 29846 18541
rect 29880 18507 29936 18541
rect 29970 18507 30026 18541
rect 30060 18507 30116 18541
rect 30150 18507 30206 18541
rect 30240 18507 30296 18541
rect 30330 18507 30386 18541
rect 30420 18507 30476 18541
rect 30510 18507 30566 18541
rect 30600 18507 30656 18541
rect 30690 18507 30746 18541
rect 30780 18518 31096 18541
rect 30780 18507 30847 18518
rect 29694 18484 30847 18507
rect 30881 18484 31000 18518
rect 31034 18507 31096 18518
rect 31130 18507 31186 18541
rect 31220 18507 31276 18541
rect 31310 18507 31366 18541
rect 31400 18507 31456 18541
rect 31490 18507 31546 18541
rect 31580 18507 31636 18541
rect 31670 18507 31726 18541
rect 31760 18507 31816 18541
rect 31850 18507 31906 18541
rect 31940 18507 31996 18541
rect 32030 18507 32086 18541
rect 32120 18518 32436 18541
rect 32120 18507 32187 18518
rect 31034 18484 32187 18507
rect 32221 18484 32340 18518
rect 32374 18507 32436 18518
rect 32470 18507 32526 18541
rect 32560 18507 32616 18541
rect 32650 18507 32706 18541
rect 32740 18507 32796 18541
rect 32830 18507 32886 18541
rect 32920 18507 32976 18541
rect 33010 18507 33066 18541
rect 33100 18507 33156 18541
rect 33190 18507 33246 18541
rect 33280 18507 33336 18541
rect 33370 18507 33426 18541
rect 33460 18518 33776 18541
rect 33460 18507 33527 18518
rect 32374 18484 33527 18507
rect 33561 18484 33680 18518
rect 33714 18507 33776 18518
rect 33810 18507 33866 18541
rect 33900 18507 33956 18541
rect 33990 18507 34046 18541
rect 34080 18507 34136 18541
rect 34170 18507 34226 18541
rect 34260 18507 34316 18541
rect 34350 18507 34406 18541
rect 34440 18507 34496 18541
rect 34530 18507 34586 18541
rect 34620 18507 34676 18541
rect 34710 18507 34766 18541
rect 34800 18518 35116 18541
rect 34800 18507 34867 18518
rect 33714 18484 34867 18507
rect 34901 18484 35020 18518
rect 35054 18507 35116 18518
rect 35150 18507 35206 18541
rect 35240 18507 35296 18541
rect 35330 18507 35386 18541
rect 35420 18507 35476 18541
rect 35510 18507 35566 18541
rect 35600 18507 35656 18541
rect 35690 18507 35746 18541
rect 35780 18507 35836 18541
rect 35870 18507 35926 18541
rect 35960 18507 36016 18541
rect 36050 18507 36106 18541
rect 36140 18518 36456 18541
rect 36140 18507 36207 18518
rect 35054 18484 36207 18507
rect 36241 18484 36360 18518
rect 36394 18507 36456 18518
rect 36490 18507 36546 18541
rect 36580 18507 36636 18541
rect 36670 18507 36726 18541
rect 36760 18507 36816 18541
rect 36850 18507 36906 18541
rect 36940 18507 36996 18541
rect 37030 18507 37086 18541
rect 37120 18507 37176 18541
rect 37210 18507 37266 18541
rect 37300 18507 37356 18541
rect 37390 18507 37446 18541
rect 37480 18518 37796 18541
rect 37480 18507 37547 18518
rect 36394 18484 37547 18507
rect 37581 18484 37700 18518
rect 37734 18507 37796 18518
rect 37830 18507 37886 18541
rect 37920 18507 37976 18541
rect 38010 18507 38066 18541
rect 38100 18507 38156 18541
rect 38190 18507 38246 18541
rect 38280 18507 38336 18541
rect 38370 18507 38426 18541
rect 38460 18507 38516 18541
rect 38550 18507 38606 18541
rect 38640 18507 38696 18541
rect 38730 18507 38786 18541
rect 38820 18518 38954 18541
rect 38820 18507 38887 18518
rect 37734 18484 38887 18507
rect 38921 18484 38954 18518
rect 28286 18475 38954 18484
rect 28286 18428 28387 18475
rect 28286 18394 28320 18428
rect 28354 18394 28387 18428
rect 29473 18428 29727 18475
rect 28286 18338 28387 18394
rect 28286 18304 28320 18338
rect 28354 18304 28387 18338
rect 28286 18248 28387 18304
rect 28286 18214 28320 18248
rect 28354 18214 28387 18248
rect 28286 18158 28387 18214
rect 28286 18124 28320 18158
rect 28354 18124 28387 18158
rect 28286 18068 28387 18124
rect 28286 18034 28320 18068
rect 28354 18034 28387 18068
rect 28286 17978 28387 18034
rect 28286 17944 28320 17978
rect 28354 17944 28387 17978
rect 28286 17888 28387 17944
rect 28286 17854 28320 17888
rect 28354 17854 28387 17888
rect 28286 17798 28387 17854
rect 28286 17764 28320 17798
rect 28354 17764 28387 17798
rect 28286 17708 28387 17764
rect 28286 17674 28320 17708
rect 28354 17674 28387 17708
rect 28286 17618 28387 17674
rect 28286 17584 28320 17618
rect 28354 17584 28387 17618
rect 28286 17528 28387 17584
rect 28286 17494 28320 17528
rect 28354 17494 28387 17528
rect 28286 17438 28387 17494
rect 29473 18394 29507 18428
rect 29541 18394 29660 18428
rect 29694 18394 29727 18428
rect 30813 18428 31067 18475
rect 29473 18338 29727 18394
rect 29473 18304 29507 18338
rect 29541 18304 29660 18338
rect 29694 18304 29727 18338
rect 29473 18248 29727 18304
rect 29473 18214 29507 18248
rect 29541 18214 29660 18248
rect 29694 18214 29727 18248
rect 29473 18158 29727 18214
rect 29473 18124 29507 18158
rect 29541 18124 29660 18158
rect 29694 18124 29727 18158
rect 29473 18068 29727 18124
rect 29473 18034 29507 18068
rect 29541 18034 29660 18068
rect 29694 18034 29727 18068
rect 29473 17978 29727 18034
rect 29473 17944 29507 17978
rect 29541 17944 29660 17978
rect 29694 17944 29727 17978
rect 29473 17888 29727 17944
rect 29473 17854 29507 17888
rect 29541 17854 29660 17888
rect 29694 17854 29727 17888
rect 29473 17798 29727 17854
rect 29473 17764 29507 17798
rect 29541 17764 29660 17798
rect 29694 17764 29727 17798
rect 29473 17708 29727 17764
rect 29473 17674 29507 17708
rect 29541 17674 29660 17708
rect 29694 17674 29727 17708
rect 29473 17618 29727 17674
rect 29473 17584 29507 17618
rect 29541 17584 29660 17618
rect 29694 17584 29727 17618
rect 29473 17528 29727 17584
rect 29473 17494 29507 17528
rect 29541 17494 29660 17528
rect 29694 17494 29727 17528
rect 28286 17404 28320 17438
rect 28354 17404 28387 17438
rect 28286 17389 28387 17404
rect 29473 17438 29727 17494
rect 30813 18394 30847 18428
rect 30881 18394 31000 18428
rect 31034 18394 31067 18428
rect 32153 18428 32407 18475
rect 30813 18338 31067 18394
rect 30813 18304 30847 18338
rect 30881 18304 31000 18338
rect 31034 18304 31067 18338
rect 30813 18248 31067 18304
rect 30813 18214 30847 18248
rect 30881 18214 31000 18248
rect 31034 18214 31067 18248
rect 30813 18158 31067 18214
rect 30813 18124 30847 18158
rect 30881 18124 31000 18158
rect 31034 18124 31067 18158
rect 30813 18068 31067 18124
rect 30813 18034 30847 18068
rect 30881 18034 31000 18068
rect 31034 18034 31067 18068
rect 30813 17978 31067 18034
rect 30813 17944 30847 17978
rect 30881 17944 31000 17978
rect 31034 17944 31067 17978
rect 30813 17888 31067 17944
rect 30813 17854 30847 17888
rect 30881 17854 31000 17888
rect 31034 17854 31067 17888
rect 30813 17798 31067 17854
rect 30813 17764 30847 17798
rect 30881 17764 31000 17798
rect 31034 17764 31067 17798
rect 30813 17708 31067 17764
rect 30813 17674 30847 17708
rect 30881 17674 31000 17708
rect 31034 17674 31067 17708
rect 30813 17618 31067 17674
rect 30813 17584 30847 17618
rect 30881 17584 31000 17618
rect 31034 17584 31067 17618
rect 30813 17528 31067 17584
rect 30813 17494 30847 17528
rect 30881 17494 31000 17528
rect 31034 17494 31067 17528
rect 29473 17404 29507 17438
rect 29541 17404 29660 17438
rect 29694 17404 29727 17438
rect 29473 17389 29727 17404
rect 30813 17438 31067 17494
rect 32153 18394 32187 18428
rect 32221 18394 32340 18428
rect 32374 18394 32407 18428
rect 33493 18428 33747 18475
rect 32153 18338 32407 18394
rect 32153 18304 32187 18338
rect 32221 18304 32340 18338
rect 32374 18304 32407 18338
rect 32153 18248 32407 18304
rect 32153 18214 32187 18248
rect 32221 18214 32340 18248
rect 32374 18214 32407 18248
rect 32153 18158 32407 18214
rect 32153 18124 32187 18158
rect 32221 18124 32340 18158
rect 32374 18124 32407 18158
rect 32153 18068 32407 18124
rect 32153 18034 32187 18068
rect 32221 18034 32340 18068
rect 32374 18034 32407 18068
rect 32153 17978 32407 18034
rect 32153 17944 32187 17978
rect 32221 17944 32340 17978
rect 32374 17944 32407 17978
rect 32153 17888 32407 17944
rect 32153 17854 32187 17888
rect 32221 17854 32340 17888
rect 32374 17854 32407 17888
rect 32153 17798 32407 17854
rect 32153 17764 32187 17798
rect 32221 17764 32340 17798
rect 32374 17764 32407 17798
rect 32153 17708 32407 17764
rect 32153 17674 32187 17708
rect 32221 17674 32340 17708
rect 32374 17674 32407 17708
rect 32153 17618 32407 17674
rect 32153 17584 32187 17618
rect 32221 17584 32340 17618
rect 32374 17584 32407 17618
rect 32153 17528 32407 17584
rect 32153 17494 32187 17528
rect 32221 17494 32340 17528
rect 32374 17494 32407 17528
rect 30813 17404 30847 17438
rect 30881 17404 31000 17438
rect 31034 17404 31067 17438
rect 30813 17389 31067 17404
rect 32153 17438 32407 17494
rect 33493 18394 33527 18428
rect 33561 18394 33680 18428
rect 33714 18394 33747 18428
rect 34833 18428 35087 18475
rect 33493 18338 33747 18394
rect 33493 18304 33527 18338
rect 33561 18304 33680 18338
rect 33714 18304 33747 18338
rect 33493 18248 33747 18304
rect 33493 18214 33527 18248
rect 33561 18214 33680 18248
rect 33714 18214 33747 18248
rect 33493 18158 33747 18214
rect 33493 18124 33527 18158
rect 33561 18124 33680 18158
rect 33714 18124 33747 18158
rect 33493 18068 33747 18124
rect 33493 18034 33527 18068
rect 33561 18034 33680 18068
rect 33714 18034 33747 18068
rect 33493 17978 33747 18034
rect 33493 17944 33527 17978
rect 33561 17944 33680 17978
rect 33714 17944 33747 17978
rect 33493 17888 33747 17944
rect 33493 17854 33527 17888
rect 33561 17854 33680 17888
rect 33714 17854 33747 17888
rect 33493 17798 33747 17854
rect 33493 17764 33527 17798
rect 33561 17764 33680 17798
rect 33714 17764 33747 17798
rect 33493 17708 33747 17764
rect 33493 17674 33527 17708
rect 33561 17674 33680 17708
rect 33714 17674 33747 17708
rect 33493 17618 33747 17674
rect 33493 17584 33527 17618
rect 33561 17584 33680 17618
rect 33714 17584 33747 17618
rect 33493 17528 33747 17584
rect 33493 17494 33527 17528
rect 33561 17494 33680 17528
rect 33714 17494 33747 17528
rect 32153 17404 32187 17438
rect 32221 17404 32340 17438
rect 32374 17404 32407 17438
rect 32153 17389 32407 17404
rect 33493 17438 33747 17494
rect 34833 18394 34867 18428
rect 34901 18394 35020 18428
rect 35054 18394 35087 18428
rect 36173 18428 36427 18475
rect 34833 18338 35087 18394
rect 34833 18304 34867 18338
rect 34901 18304 35020 18338
rect 35054 18304 35087 18338
rect 34833 18248 35087 18304
rect 34833 18214 34867 18248
rect 34901 18214 35020 18248
rect 35054 18214 35087 18248
rect 34833 18158 35087 18214
rect 34833 18124 34867 18158
rect 34901 18124 35020 18158
rect 35054 18124 35087 18158
rect 34833 18068 35087 18124
rect 34833 18034 34867 18068
rect 34901 18034 35020 18068
rect 35054 18034 35087 18068
rect 34833 17978 35087 18034
rect 34833 17944 34867 17978
rect 34901 17944 35020 17978
rect 35054 17944 35087 17978
rect 34833 17888 35087 17944
rect 34833 17854 34867 17888
rect 34901 17854 35020 17888
rect 35054 17854 35087 17888
rect 34833 17798 35087 17854
rect 34833 17764 34867 17798
rect 34901 17764 35020 17798
rect 35054 17764 35087 17798
rect 34833 17708 35087 17764
rect 34833 17674 34867 17708
rect 34901 17674 35020 17708
rect 35054 17674 35087 17708
rect 34833 17618 35087 17674
rect 34833 17584 34867 17618
rect 34901 17584 35020 17618
rect 35054 17584 35087 17618
rect 34833 17528 35087 17584
rect 34833 17494 34867 17528
rect 34901 17494 35020 17528
rect 35054 17494 35087 17528
rect 33493 17404 33527 17438
rect 33561 17404 33680 17438
rect 33714 17404 33747 17438
rect 33493 17389 33747 17404
rect 34833 17438 35087 17494
rect 36173 18394 36207 18428
rect 36241 18394 36360 18428
rect 36394 18394 36427 18428
rect 37513 18428 37767 18475
rect 36173 18338 36427 18394
rect 36173 18304 36207 18338
rect 36241 18304 36360 18338
rect 36394 18304 36427 18338
rect 36173 18248 36427 18304
rect 36173 18214 36207 18248
rect 36241 18214 36360 18248
rect 36394 18214 36427 18248
rect 36173 18158 36427 18214
rect 36173 18124 36207 18158
rect 36241 18124 36360 18158
rect 36394 18124 36427 18158
rect 36173 18068 36427 18124
rect 36173 18034 36207 18068
rect 36241 18034 36360 18068
rect 36394 18034 36427 18068
rect 36173 17978 36427 18034
rect 36173 17944 36207 17978
rect 36241 17944 36360 17978
rect 36394 17944 36427 17978
rect 36173 17888 36427 17944
rect 36173 17854 36207 17888
rect 36241 17854 36360 17888
rect 36394 17854 36427 17888
rect 36173 17798 36427 17854
rect 36173 17764 36207 17798
rect 36241 17764 36360 17798
rect 36394 17764 36427 17798
rect 36173 17708 36427 17764
rect 36173 17674 36207 17708
rect 36241 17674 36360 17708
rect 36394 17674 36427 17708
rect 36173 17618 36427 17674
rect 36173 17584 36207 17618
rect 36241 17584 36360 17618
rect 36394 17584 36427 17618
rect 36173 17528 36427 17584
rect 36173 17494 36207 17528
rect 36241 17494 36360 17528
rect 36394 17494 36427 17528
rect 34833 17404 34867 17438
rect 34901 17404 35020 17438
rect 35054 17404 35087 17438
rect 34833 17389 35087 17404
rect 36173 17438 36427 17494
rect 37513 18394 37547 18428
rect 37581 18394 37700 18428
rect 37734 18394 37767 18428
rect 38853 18428 38954 18475
rect 37513 18338 37767 18394
rect 37513 18304 37547 18338
rect 37581 18304 37700 18338
rect 37734 18304 37767 18338
rect 37513 18248 37767 18304
rect 37513 18214 37547 18248
rect 37581 18214 37700 18248
rect 37734 18214 37767 18248
rect 37513 18158 37767 18214
rect 37513 18124 37547 18158
rect 37581 18124 37700 18158
rect 37734 18124 37767 18158
rect 37513 18068 37767 18124
rect 37513 18034 37547 18068
rect 37581 18034 37700 18068
rect 37734 18034 37767 18068
rect 37513 17978 37767 18034
rect 37513 17944 37547 17978
rect 37581 17944 37700 17978
rect 37734 17944 37767 17978
rect 37513 17888 37767 17944
rect 37513 17854 37547 17888
rect 37581 17854 37700 17888
rect 37734 17854 37767 17888
rect 37513 17798 37767 17854
rect 37513 17764 37547 17798
rect 37581 17764 37700 17798
rect 37734 17764 37767 17798
rect 37513 17708 37767 17764
rect 37513 17674 37547 17708
rect 37581 17674 37700 17708
rect 37734 17674 37767 17708
rect 37513 17618 37767 17674
rect 37513 17584 37547 17618
rect 37581 17584 37700 17618
rect 37734 17584 37767 17618
rect 37513 17528 37767 17584
rect 37513 17494 37547 17528
rect 37581 17494 37700 17528
rect 37734 17494 37767 17528
rect 36173 17404 36207 17438
rect 36241 17404 36360 17438
rect 36394 17404 36427 17438
rect 36173 17389 36427 17404
rect 37513 17438 37767 17494
rect 38853 18394 38887 18428
rect 38921 18394 38954 18428
rect 38853 18338 38954 18394
rect 38853 18304 38887 18338
rect 38921 18304 38954 18338
rect 38853 18248 38954 18304
rect 38853 18214 38887 18248
rect 38921 18214 38954 18248
rect 38853 18158 38954 18214
rect 38853 18124 38887 18158
rect 38921 18124 38954 18158
rect 38853 18068 38954 18124
rect 38853 18034 38887 18068
rect 38921 18034 38954 18068
rect 38853 17978 38954 18034
rect 38853 17944 38887 17978
rect 38921 17944 38954 17978
rect 38853 17888 38954 17944
rect 38853 17854 38887 17888
rect 38921 17854 38954 17888
rect 38853 17798 38954 17854
rect 38853 17764 38887 17798
rect 38921 17764 38954 17798
rect 40168 17923 40784 17962
rect 40168 17821 40255 17923
rect 40697 17821 40784 17923
rect 40168 17782 40784 17821
rect 38853 17708 38954 17764
rect 38853 17674 38887 17708
rect 38921 17674 38954 17708
rect 38853 17618 38954 17674
rect 38853 17584 38887 17618
rect 38921 17584 38954 17618
rect 38853 17528 38954 17584
rect 38853 17494 38887 17528
rect 38921 17494 38954 17528
rect 37513 17404 37547 17438
rect 37581 17404 37700 17438
rect 37734 17404 37767 17438
rect 37513 17389 37767 17404
rect 38853 17438 38954 17494
rect 38853 17404 38887 17438
rect 38921 17404 38954 17438
rect 38853 17389 38954 17404
rect 28286 17354 38954 17389
rect 28286 17320 28416 17354
rect 28450 17320 28506 17354
rect 28540 17320 28596 17354
rect 28630 17320 28686 17354
rect 28720 17320 28776 17354
rect 28810 17320 28866 17354
rect 28900 17320 28956 17354
rect 28990 17320 29046 17354
rect 29080 17320 29136 17354
rect 29170 17320 29226 17354
rect 29260 17320 29316 17354
rect 29350 17320 29406 17354
rect 29440 17320 29756 17354
rect 29790 17320 29846 17354
rect 29880 17320 29936 17354
rect 29970 17320 30026 17354
rect 30060 17320 30116 17354
rect 30150 17320 30206 17354
rect 30240 17320 30296 17354
rect 30330 17320 30386 17354
rect 30420 17320 30476 17354
rect 30510 17320 30566 17354
rect 30600 17320 30656 17354
rect 30690 17320 30746 17354
rect 30780 17320 31096 17354
rect 31130 17320 31186 17354
rect 31220 17320 31276 17354
rect 31310 17320 31366 17354
rect 31400 17320 31456 17354
rect 31490 17320 31546 17354
rect 31580 17320 31636 17354
rect 31670 17320 31726 17354
rect 31760 17320 31816 17354
rect 31850 17320 31906 17354
rect 31940 17320 31996 17354
rect 32030 17320 32086 17354
rect 32120 17320 32436 17354
rect 32470 17320 32526 17354
rect 32560 17320 32616 17354
rect 32650 17320 32706 17354
rect 32740 17320 32796 17354
rect 32830 17320 32886 17354
rect 32920 17320 32976 17354
rect 33010 17320 33066 17354
rect 33100 17320 33156 17354
rect 33190 17320 33246 17354
rect 33280 17320 33336 17354
rect 33370 17320 33426 17354
rect 33460 17320 33776 17354
rect 33810 17320 33866 17354
rect 33900 17320 33956 17354
rect 33990 17320 34046 17354
rect 34080 17320 34136 17354
rect 34170 17320 34226 17354
rect 34260 17320 34316 17354
rect 34350 17320 34406 17354
rect 34440 17320 34496 17354
rect 34530 17320 34586 17354
rect 34620 17320 34676 17354
rect 34710 17320 34766 17354
rect 34800 17320 35116 17354
rect 35150 17320 35206 17354
rect 35240 17320 35296 17354
rect 35330 17320 35386 17354
rect 35420 17320 35476 17354
rect 35510 17320 35566 17354
rect 35600 17320 35656 17354
rect 35690 17320 35746 17354
rect 35780 17320 35836 17354
rect 35870 17320 35926 17354
rect 35960 17320 36016 17354
rect 36050 17320 36106 17354
rect 36140 17320 36456 17354
rect 36490 17320 36546 17354
rect 36580 17320 36636 17354
rect 36670 17320 36726 17354
rect 36760 17320 36816 17354
rect 36850 17320 36906 17354
rect 36940 17320 36996 17354
rect 37030 17320 37086 17354
rect 37120 17320 37176 17354
rect 37210 17320 37266 17354
rect 37300 17320 37356 17354
rect 37390 17320 37446 17354
rect 37480 17320 37796 17354
rect 37830 17320 37886 17354
rect 37920 17320 37976 17354
rect 38010 17320 38066 17354
rect 38100 17320 38156 17354
rect 38190 17320 38246 17354
rect 38280 17320 38336 17354
rect 38370 17320 38426 17354
rect 38460 17320 38516 17354
rect 38550 17320 38606 17354
rect 38640 17320 38696 17354
rect 38730 17320 38786 17354
rect 38820 17320 38954 17354
rect 28286 17288 38954 17320
rect 8314 17072 8434 17085
rect 28286 14781 38954 14816
rect 28286 14758 28416 14781
rect 28286 14724 28320 14758
rect 28354 14747 28416 14758
rect 28450 14747 28506 14781
rect 28540 14747 28596 14781
rect 28630 14747 28686 14781
rect 28720 14747 28776 14781
rect 28810 14747 28866 14781
rect 28900 14747 28956 14781
rect 28990 14747 29046 14781
rect 29080 14747 29136 14781
rect 29170 14747 29226 14781
rect 29260 14747 29316 14781
rect 29350 14747 29406 14781
rect 29440 14758 29756 14781
rect 29440 14747 29507 14758
rect 28354 14724 29507 14747
rect 29541 14724 29660 14758
rect 29694 14747 29756 14758
rect 29790 14747 29846 14781
rect 29880 14747 29936 14781
rect 29970 14747 30026 14781
rect 30060 14747 30116 14781
rect 30150 14747 30206 14781
rect 30240 14747 30296 14781
rect 30330 14747 30386 14781
rect 30420 14747 30476 14781
rect 30510 14747 30566 14781
rect 30600 14747 30656 14781
rect 30690 14747 30746 14781
rect 30780 14758 31096 14781
rect 30780 14747 30847 14758
rect 29694 14724 30847 14747
rect 30881 14724 31000 14758
rect 31034 14747 31096 14758
rect 31130 14747 31186 14781
rect 31220 14747 31276 14781
rect 31310 14747 31366 14781
rect 31400 14747 31456 14781
rect 31490 14747 31546 14781
rect 31580 14747 31636 14781
rect 31670 14747 31726 14781
rect 31760 14747 31816 14781
rect 31850 14747 31906 14781
rect 31940 14747 31996 14781
rect 32030 14747 32086 14781
rect 32120 14758 32436 14781
rect 32120 14747 32187 14758
rect 31034 14724 32187 14747
rect 32221 14724 32340 14758
rect 32374 14747 32436 14758
rect 32470 14747 32526 14781
rect 32560 14747 32616 14781
rect 32650 14747 32706 14781
rect 32740 14747 32796 14781
rect 32830 14747 32886 14781
rect 32920 14747 32976 14781
rect 33010 14747 33066 14781
rect 33100 14747 33156 14781
rect 33190 14747 33246 14781
rect 33280 14747 33336 14781
rect 33370 14747 33426 14781
rect 33460 14758 33776 14781
rect 33460 14747 33527 14758
rect 32374 14724 33527 14747
rect 33561 14724 33680 14758
rect 33714 14747 33776 14758
rect 33810 14747 33866 14781
rect 33900 14747 33956 14781
rect 33990 14747 34046 14781
rect 34080 14747 34136 14781
rect 34170 14747 34226 14781
rect 34260 14747 34316 14781
rect 34350 14747 34406 14781
rect 34440 14747 34496 14781
rect 34530 14747 34586 14781
rect 34620 14747 34676 14781
rect 34710 14747 34766 14781
rect 34800 14758 35116 14781
rect 34800 14747 34867 14758
rect 33714 14724 34867 14747
rect 34901 14724 35020 14758
rect 35054 14747 35116 14758
rect 35150 14747 35206 14781
rect 35240 14747 35296 14781
rect 35330 14747 35386 14781
rect 35420 14747 35476 14781
rect 35510 14747 35566 14781
rect 35600 14747 35656 14781
rect 35690 14747 35746 14781
rect 35780 14747 35836 14781
rect 35870 14747 35926 14781
rect 35960 14747 36016 14781
rect 36050 14747 36106 14781
rect 36140 14758 36456 14781
rect 36140 14747 36207 14758
rect 35054 14724 36207 14747
rect 36241 14724 36360 14758
rect 36394 14747 36456 14758
rect 36490 14747 36546 14781
rect 36580 14747 36636 14781
rect 36670 14747 36726 14781
rect 36760 14747 36816 14781
rect 36850 14747 36906 14781
rect 36940 14747 36996 14781
rect 37030 14747 37086 14781
rect 37120 14747 37176 14781
rect 37210 14747 37266 14781
rect 37300 14747 37356 14781
rect 37390 14747 37446 14781
rect 37480 14758 37796 14781
rect 37480 14747 37547 14758
rect 36394 14724 37547 14747
rect 37581 14724 37700 14758
rect 37734 14747 37796 14758
rect 37830 14747 37886 14781
rect 37920 14747 37976 14781
rect 38010 14747 38066 14781
rect 38100 14747 38156 14781
rect 38190 14747 38246 14781
rect 38280 14747 38336 14781
rect 38370 14747 38426 14781
rect 38460 14747 38516 14781
rect 38550 14747 38606 14781
rect 38640 14747 38696 14781
rect 38730 14747 38786 14781
rect 38820 14758 38954 14781
rect 38820 14747 38887 14758
rect 37734 14724 38887 14747
rect 38921 14724 38954 14758
rect 28286 14715 38954 14724
rect 28286 14668 28387 14715
rect 28286 14634 28320 14668
rect 28354 14634 28387 14668
rect 29473 14668 29727 14715
rect 28286 14578 28387 14634
rect 28286 14544 28320 14578
rect 28354 14544 28387 14578
rect 28286 14488 28387 14544
rect 28286 14454 28320 14488
rect 28354 14454 28387 14488
rect 28286 14398 28387 14454
rect 28286 14364 28320 14398
rect 28354 14364 28387 14398
rect 28286 14308 28387 14364
rect 28286 14274 28320 14308
rect 28354 14274 28387 14308
rect 28286 14218 28387 14274
rect 8808 14163 9424 14202
rect 8808 14061 8895 14163
rect 9337 14061 9424 14163
rect 8808 14022 9424 14061
rect 11552 14163 12168 14202
rect 11552 14061 11639 14163
rect 12081 14061 12168 14163
rect 11552 14022 12168 14061
rect 14296 14163 14912 14202
rect 14296 14061 14383 14163
rect 14825 14061 14912 14163
rect 14296 14022 14912 14061
rect 24488 14163 25104 14202
rect 24488 14061 24575 14163
rect 25017 14061 25104 14163
rect 24488 14022 25104 14061
rect 28286 14184 28320 14218
rect 28354 14184 28387 14218
rect 28286 14128 28387 14184
rect 28286 14094 28320 14128
rect 28354 14094 28387 14128
rect 28286 14038 28387 14094
rect 28286 14004 28320 14038
rect 28354 14004 28387 14038
rect 28286 13948 28387 14004
rect 28286 13914 28320 13948
rect 28354 13914 28387 13948
rect 28286 13858 28387 13914
rect 28286 13824 28320 13858
rect 28354 13824 28387 13858
rect 28286 13768 28387 13824
rect 28286 13734 28320 13768
rect 28354 13734 28387 13768
rect 28286 13678 28387 13734
rect 29473 14634 29507 14668
rect 29541 14634 29660 14668
rect 29694 14634 29727 14668
rect 30813 14668 31067 14715
rect 29473 14578 29727 14634
rect 29473 14544 29507 14578
rect 29541 14544 29660 14578
rect 29694 14544 29727 14578
rect 29473 14488 29727 14544
rect 29473 14454 29507 14488
rect 29541 14454 29660 14488
rect 29694 14454 29727 14488
rect 29473 14398 29727 14454
rect 29473 14364 29507 14398
rect 29541 14364 29660 14398
rect 29694 14364 29727 14398
rect 29473 14308 29727 14364
rect 29473 14274 29507 14308
rect 29541 14274 29660 14308
rect 29694 14274 29727 14308
rect 29473 14218 29727 14274
rect 29473 14184 29507 14218
rect 29541 14184 29660 14218
rect 29694 14184 29727 14218
rect 29473 14128 29727 14184
rect 29473 14094 29507 14128
rect 29541 14094 29660 14128
rect 29694 14094 29727 14128
rect 29473 14038 29727 14094
rect 29473 14004 29507 14038
rect 29541 14004 29660 14038
rect 29694 14004 29727 14038
rect 29473 13948 29727 14004
rect 29473 13914 29507 13948
rect 29541 13914 29660 13948
rect 29694 13914 29727 13948
rect 29473 13858 29727 13914
rect 29473 13824 29507 13858
rect 29541 13824 29660 13858
rect 29694 13824 29727 13858
rect 29473 13768 29727 13824
rect 29473 13734 29507 13768
rect 29541 13734 29660 13768
rect 29694 13734 29727 13768
rect 28286 13644 28320 13678
rect 28354 13644 28387 13678
rect 28286 13629 28387 13644
rect 29473 13678 29727 13734
rect 30813 14634 30847 14668
rect 30881 14634 31000 14668
rect 31034 14634 31067 14668
rect 32153 14668 32407 14715
rect 30813 14578 31067 14634
rect 30813 14544 30847 14578
rect 30881 14544 31000 14578
rect 31034 14544 31067 14578
rect 30813 14488 31067 14544
rect 30813 14454 30847 14488
rect 30881 14454 31000 14488
rect 31034 14454 31067 14488
rect 30813 14398 31067 14454
rect 30813 14364 30847 14398
rect 30881 14364 31000 14398
rect 31034 14364 31067 14398
rect 30813 14308 31067 14364
rect 30813 14274 30847 14308
rect 30881 14274 31000 14308
rect 31034 14274 31067 14308
rect 30813 14218 31067 14274
rect 30813 14184 30847 14218
rect 30881 14184 31000 14218
rect 31034 14184 31067 14218
rect 30813 14128 31067 14184
rect 30813 14094 30847 14128
rect 30881 14094 31000 14128
rect 31034 14094 31067 14128
rect 30813 14038 31067 14094
rect 30813 14004 30847 14038
rect 30881 14004 31000 14038
rect 31034 14004 31067 14038
rect 30813 13948 31067 14004
rect 30813 13914 30847 13948
rect 30881 13914 31000 13948
rect 31034 13914 31067 13948
rect 30813 13858 31067 13914
rect 30813 13824 30847 13858
rect 30881 13824 31000 13858
rect 31034 13824 31067 13858
rect 30813 13768 31067 13824
rect 30813 13734 30847 13768
rect 30881 13734 31000 13768
rect 31034 13734 31067 13768
rect 29473 13644 29507 13678
rect 29541 13644 29660 13678
rect 29694 13644 29727 13678
rect 29473 13629 29727 13644
rect 30813 13678 31067 13734
rect 32153 14634 32187 14668
rect 32221 14634 32340 14668
rect 32374 14634 32407 14668
rect 33493 14668 33747 14715
rect 32153 14578 32407 14634
rect 32153 14544 32187 14578
rect 32221 14544 32340 14578
rect 32374 14544 32407 14578
rect 32153 14488 32407 14544
rect 32153 14454 32187 14488
rect 32221 14454 32340 14488
rect 32374 14454 32407 14488
rect 32153 14398 32407 14454
rect 32153 14364 32187 14398
rect 32221 14364 32340 14398
rect 32374 14364 32407 14398
rect 32153 14308 32407 14364
rect 32153 14274 32187 14308
rect 32221 14274 32340 14308
rect 32374 14274 32407 14308
rect 32153 14218 32407 14274
rect 32153 14184 32187 14218
rect 32221 14184 32340 14218
rect 32374 14184 32407 14218
rect 32153 14128 32407 14184
rect 32153 14094 32187 14128
rect 32221 14094 32340 14128
rect 32374 14094 32407 14128
rect 32153 14038 32407 14094
rect 32153 14004 32187 14038
rect 32221 14004 32340 14038
rect 32374 14004 32407 14038
rect 32153 13948 32407 14004
rect 32153 13914 32187 13948
rect 32221 13914 32340 13948
rect 32374 13914 32407 13948
rect 32153 13858 32407 13914
rect 32153 13824 32187 13858
rect 32221 13824 32340 13858
rect 32374 13824 32407 13858
rect 32153 13768 32407 13824
rect 32153 13734 32187 13768
rect 32221 13734 32340 13768
rect 32374 13734 32407 13768
rect 30813 13644 30847 13678
rect 30881 13644 31000 13678
rect 31034 13644 31067 13678
rect 30813 13629 31067 13644
rect 32153 13678 32407 13734
rect 33493 14634 33527 14668
rect 33561 14634 33680 14668
rect 33714 14634 33747 14668
rect 34833 14668 35087 14715
rect 33493 14578 33747 14634
rect 33493 14544 33527 14578
rect 33561 14544 33680 14578
rect 33714 14544 33747 14578
rect 33493 14488 33747 14544
rect 33493 14454 33527 14488
rect 33561 14454 33680 14488
rect 33714 14454 33747 14488
rect 33493 14398 33747 14454
rect 33493 14364 33527 14398
rect 33561 14364 33680 14398
rect 33714 14364 33747 14398
rect 33493 14308 33747 14364
rect 33493 14274 33527 14308
rect 33561 14274 33680 14308
rect 33714 14274 33747 14308
rect 33493 14218 33747 14274
rect 33493 14184 33527 14218
rect 33561 14184 33680 14218
rect 33714 14184 33747 14218
rect 33493 14128 33747 14184
rect 33493 14094 33527 14128
rect 33561 14094 33680 14128
rect 33714 14094 33747 14128
rect 33493 14038 33747 14094
rect 33493 14004 33527 14038
rect 33561 14004 33680 14038
rect 33714 14004 33747 14038
rect 33493 13948 33747 14004
rect 33493 13914 33527 13948
rect 33561 13914 33680 13948
rect 33714 13914 33747 13948
rect 33493 13858 33747 13914
rect 33493 13824 33527 13858
rect 33561 13824 33680 13858
rect 33714 13824 33747 13858
rect 33493 13768 33747 13824
rect 33493 13734 33527 13768
rect 33561 13734 33680 13768
rect 33714 13734 33747 13768
rect 32153 13644 32187 13678
rect 32221 13644 32340 13678
rect 32374 13644 32407 13678
rect 32153 13629 32407 13644
rect 33493 13678 33747 13734
rect 34833 14634 34867 14668
rect 34901 14634 35020 14668
rect 35054 14634 35087 14668
rect 36173 14668 36427 14715
rect 34833 14578 35087 14634
rect 34833 14544 34867 14578
rect 34901 14544 35020 14578
rect 35054 14544 35087 14578
rect 34833 14488 35087 14544
rect 34833 14454 34867 14488
rect 34901 14454 35020 14488
rect 35054 14454 35087 14488
rect 34833 14398 35087 14454
rect 34833 14364 34867 14398
rect 34901 14364 35020 14398
rect 35054 14364 35087 14398
rect 34833 14308 35087 14364
rect 34833 14274 34867 14308
rect 34901 14274 35020 14308
rect 35054 14274 35087 14308
rect 34833 14218 35087 14274
rect 34833 14184 34867 14218
rect 34901 14184 35020 14218
rect 35054 14184 35087 14218
rect 34833 14128 35087 14184
rect 34833 14094 34867 14128
rect 34901 14094 35020 14128
rect 35054 14094 35087 14128
rect 34833 14038 35087 14094
rect 34833 14004 34867 14038
rect 34901 14004 35020 14038
rect 35054 14004 35087 14038
rect 34833 13948 35087 14004
rect 34833 13914 34867 13948
rect 34901 13914 35020 13948
rect 35054 13914 35087 13948
rect 34833 13858 35087 13914
rect 34833 13824 34867 13858
rect 34901 13824 35020 13858
rect 35054 13824 35087 13858
rect 34833 13768 35087 13824
rect 34833 13734 34867 13768
rect 34901 13734 35020 13768
rect 35054 13734 35087 13768
rect 33493 13644 33527 13678
rect 33561 13644 33680 13678
rect 33714 13644 33747 13678
rect 33493 13629 33747 13644
rect 34833 13678 35087 13734
rect 36173 14634 36207 14668
rect 36241 14634 36360 14668
rect 36394 14634 36427 14668
rect 37513 14668 37767 14715
rect 36173 14578 36427 14634
rect 36173 14544 36207 14578
rect 36241 14544 36360 14578
rect 36394 14544 36427 14578
rect 36173 14488 36427 14544
rect 36173 14454 36207 14488
rect 36241 14454 36360 14488
rect 36394 14454 36427 14488
rect 36173 14398 36427 14454
rect 36173 14364 36207 14398
rect 36241 14364 36360 14398
rect 36394 14364 36427 14398
rect 36173 14308 36427 14364
rect 36173 14274 36207 14308
rect 36241 14274 36360 14308
rect 36394 14274 36427 14308
rect 36173 14218 36427 14274
rect 36173 14184 36207 14218
rect 36241 14184 36360 14218
rect 36394 14184 36427 14218
rect 36173 14128 36427 14184
rect 36173 14094 36207 14128
rect 36241 14094 36360 14128
rect 36394 14094 36427 14128
rect 36173 14038 36427 14094
rect 36173 14004 36207 14038
rect 36241 14004 36360 14038
rect 36394 14004 36427 14038
rect 36173 13948 36427 14004
rect 36173 13914 36207 13948
rect 36241 13914 36360 13948
rect 36394 13914 36427 13948
rect 36173 13858 36427 13914
rect 36173 13824 36207 13858
rect 36241 13824 36360 13858
rect 36394 13824 36427 13858
rect 36173 13768 36427 13824
rect 36173 13734 36207 13768
rect 36241 13734 36360 13768
rect 36394 13734 36427 13768
rect 34833 13644 34867 13678
rect 34901 13644 35020 13678
rect 35054 13644 35087 13678
rect 34833 13629 35087 13644
rect 36173 13678 36427 13734
rect 37513 14634 37547 14668
rect 37581 14634 37700 14668
rect 37734 14634 37767 14668
rect 38853 14668 38954 14715
rect 37513 14578 37767 14634
rect 37513 14544 37547 14578
rect 37581 14544 37700 14578
rect 37734 14544 37767 14578
rect 37513 14488 37767 14544
rect 37513 14454 37547 14488
rect 37581 14454 37700 14488
rect 37734 14454 37767 14488
rect 37513 14398 37767 14454
rect 37513 14364 37547 14398
rect 37581 14364 37700 14398
rect 37734 14364 37767 14398
rect 37513 14308 37767 14364
rect 37513 14274 37547 14308
rect 37581 14274 37700 14308
rect 37734 14274 37767 14308
rect 37513 14218 37767 14274
rect 37513 14184 37547 14218
rect 37581 14184 37700 14218
rect 37734 14184 37767 14218
rect 37513 14128 37767 14184
rect 37513 14094 37547 14128
rect 37581 14094 37700 14128
rect 37734 14094 37767 14128
rect 37513 14038 37767 14094
rect 37513 14004 37547 14038
rect 37581 14004 37700 14038
rect 37734 14004 37767 14038
rect 37513 13948 37767 14004
rect 37513 13914 37547 13948
rect 37581 13914 37700 13948
rect 37734 13914 37767 13948
rect 37513 13858 37767 13914
rect 37513 13824 37547 13858
rect 37581 13824 37700 13858
rect 37734 13824 37767 13858
rect 37513 13768 37767 13824
rect 37513 13734 37547 13768
rect 37581 13734 37700 13768
rect 37734 13734 37767 13768
rect 36173 13644 36207 13678
rect 36241 13644 36360 13678
rect 36394 13644 36427 13678
rect 36173 13629 36427 13644
rect 37513 13678 37767 13734
rect 38853 14634 38887 14668
rect 38921 14634 38954 14668
rect 38853 14578 38954 14634
rect 38853 14544 38887 14578
rect 38921 14544 38954 14578
rect 38853 14488 38954 14544
rect 38853 14454 38887 14488
rect 38921 14454 38954 14488
rect 38853 14398 38954 14454
rect 38853 14364 38887 14398
rect 38921 14364 38954 14398
rect 38853 14308 38954 14364
rect 38853 14274 38887 14308
rect 38921 14274 38954 14308
rect 38853 14218 38954 14274
rect 38853 14184 38887 14218
rect 38921 14184 38954 14218
rect 38853 14128 38954 14184
rect 38853 14094 38887 14128
rect 38921 14094 38954 14128
rect 38853 14038 38954 14094
rect 38853 14004 38887 14038
rect 38921 14004 38954 14038
rect 40168 14163 40784 14202
rect 40168 14061 40255 14163
rect 40697 14061 40784 14163
rect 40168 14022 40784 14061
rect 38853 13948 38954 14004
rect 38853 13914 38887 13948
rect 38921 13914 38954 13948
rect 38853 13858 38954 13914
rect 38853 13824 38887 13858
rect 38921 13824 38954 13858
rect 38853 13768 38954 13824
rect 38853 13734 38887 13768
rect 38921 13734 38954 13768
rect 37513 13644 37547 13678
rect 37581 13644 37700 13678
rect 37734 13644 37767 13678
rect 37513 13629 37767 13644
rect 38853 13678 38954 13734
rect 38853 13644 38887 13678
rect 38921 13644 38954 13678
rect 38853 13629 38954 13644
rect 28286 13594 38954 13629
rect 28286 13560 28416 13594
rect 28450 13560 28506 13594
rect 28540 13560 28596 13594
rect 28630 13560 28686 13594
rect 28720 13560 28776 13594
rect 28810 13560 28866 13594
rect 28900 13560 28956 13594
rect 28990 13560 29046 13594
rect 29080 13560 29136 13594
rect 29170 13560 29226 13594
rect 29260 13560 29316 13594
rect 29350 13560 29406 13594
rect 29440 13560 29756 13594
rect 29790 13560 29846 13594
rect 29880 13560 29936 13594
rect 29970 13560 30026 13594
rect 30060 13560 30116 13594
rect 30150 13560 30206 13594
rect 30240 13560 30296 13594
rect 30330 13560 30386 13594
rect 30420 13560 30476 13594
rect 30510 13560 30566 13594
rect 30600 13560 30656 13594
rect 30690 13560 30746 13594
rect 30780 13560 31096 13594
rect 31130 13560 31186 13594
rect 31220 13560 31276 13594
rect 31310 13560 31366 13594
rect 31400 13560 31456 13594
rect 31490 13560 31546 13594
rect 31580 13560 31636 13594
rect 31670 13560 31726 13594
rect 31760 13560 31816 13594
rect 31850 13560 31906 13594
rect 31940 13560 31996 13594
rect 32030 13560 32086 13594
rect 32120 13560 32436 13594
rect 32470 13560 32526 13594
rect 32560 13560 32616 13594
rect 32650 13560 32706 13594
rect 32740 13560 32796 13594
rect 32830 13560 32886 13594
rect 32920 13560 32976 13594
rect 33010 13560 33066 13594
rect 33100 13560 33156 13594
rect 33190 13560 33246 13594
rect 33280 13560 33336 13594
rect 33370 13560 33426 13594
rect 33460 13560 33776 13594
rect 33810 13560 33866 13594
rect 33900 13560 33956 13594
rect 33990 13560 34046 13594
rect 34080 13560 34136 13594
rect 34170 13560 34226 13594
rect 34260 13560 34316 13594
rect 34350 13560 34406 13594
rect 34440 13560 34496 13594
rect 34530 13560 34586 13594
rect 34620 13560 34676 13594
rect 34710 13560 34766 13594
rect 34800 13560 35116 13594
rect 35150 13560 35206 13594
rect 35240 13560 35296 13594
rect 35330 13560 35386 13594
rect 35420 13560 35476 13594
rect 35510 13560 35566 13594
rect 35600 13560 35656 13594
rect 35690 13560 35746 13594
rect 35780 13560 35836 13594
rect 35870 13560 35926 13594
rect 35960 13560 36016 13594
rect 36050 13560 36106 13594
rect 36140 13560 36456 13594
rect 36490 13560 36546 13594
rect 36580 13560 36636 13594
rect 36670 13560 36726 13594
rect 36760 13560 36816 13594
rect 36850 13560 36906 13594
rect 36940 13560 36996 13594
rect 37030 13560 37086 13594
rect 37120 13560 37176 13594
rect 37210 13560 37266 13594
rect 37300 13560 37356 13594
rect 37390 13560 37446 13594
rect 37480 13560 37796 13594
rect 37830 13560 37886 13594
rect 37920 13560 37976 13594
rect 38010 13560 38066 13594
rect 38100 13560 38156 13594
rect 38190 13560 38246 13594
rect 38280 13560 38336 13594
rect 38370 13560 38426 13594
rect 38460 13560 38516 13594
rect 38550 13560 38606 13594
rect 38640 13560 38696 13594
rect 38730 13560 38786 13594
rect 38820 13560 38954 13594
rect 28286 13528 38954 13560
rect 8808 10403 9424 10442
rect 8808 10301 8895 10403
rect 9337 10301 9424 10403
rect 8808 10262 9424 10301
rect 11552 10403 12168 10442
rect 11552 10301 11639 10403
rect 12081 10301 12168 10403
rect 11552 10262 12168 10301
rect 14296 10403 14912 10442
rect 14296 10301 14383 10403
rect 14825 10301 14912 10403
rect 14296 10262 14912 10301
rect 24776 10403 25392 10442
rect 24776 10301 24863 10403
rect 25305 10301 25392 10403
rect 24776 10262 25392 10301
rect 27820 10403 28436 10442
rect 27820 10301 27907 10403
rect 28349 10301 28436 10403
rect 27820 10262 28436 10301
rect 30564 10403 31180 10442
rect 30564 10301 30651 10403
rect 31093 10301 31180 10403
rect 30564 10262 31180 10301
rect 33308 10403 33924 10442
rect 33308 10301 33395 10403
rect 33837 10301 33924 10403
rect 33308 10262 33924 10301
rect 36052 10403 36668 10442
rect 36052 10301 36139 10403
rect 36581 10301 36668 10403
rect 36052 10262 36668 10301
rect 38796 10403 39412 10442
rect 38796 10301 38883 10403
rect 39325 10301 39412 10403
rect 38796 10262 39412 10301
rect 8808 6643 9424 6682
rect 8808 6541 8895 6643
rect 9337 6541 9424 6643
rect 8808 6502 9424 6541
rect 15466 6643 16082 6682
rect 15466 6541 15553 6643
rect 15995 6541 16082 6643
rect 15466 6502 16082 6541
rect 18510 6643 19126 6682
rect 18510 6541 18597 6643
rect 19039 6541 19126 6643
rect 18510 6502 19126 6541
rect 21254 6643 21870 6682
rect 21254 6541 21341 6643
rect 21783 6541 21870 6643
rect 21254 6502 21870 6541
rect 23998 6643 24614 6682
rect 23998 6541 24085 6643
rect 24527 6541 24614 6643
rect 23998 6502 24614 6541
rect 26742 6643 27358 6682
rect 26742 6541 26829 6643
rect 27271 6541 27358 6643
rect 26742 6502 27358 6541
rect 29486 6643 30102 6682
rect 29486 6541 29573 6643
rect 30015 6541 30102 6643
rect 29486 6502 30102 6541
rect 32230 6643 32846 6682
rect 32230 6541 32317 6643
rect 32759 6541 32846 6643
rect 32230 6502 32846 6541
rect 36052 6643 36668 6682
rect 36052 6541 36139 6643
rect 36581 6541 36668 6643
rect 36052 6502 36668 6541
rect 38796 6643 39412 6682
rect 38796 6541 38883 6643
rect 39325 6541 39412 6643
rect 38796 6502 39412 6541
<< nsubdiff >>
rect 16028 41359 16148 41362
rect 14970 41309 15010 41352
rect 16028 41325 16073 41359
rect 16107 41325 16148 41359
rect 16028 41322 16148 41325
rect 17328 41359 17448 41362
rect 17328 41325 17373 41359
rect 17407 41325 17448 41359
rect 17328 41322 17448 41325
rect 18628 41359 18748 41362
rect 18628 41325 18673 41359
rect 18707 41325 18748 41359
rect 18628 41322 18748 41325
rect 19928 41359 20048 41362
rect 19928 41325 19973 41359
rect 20007 41325 20048 41359
rect 19928 41322 20048 41325
rect 21228 41359 21348 41362
rect 21228 41325 21273 41359
rect 21307 41325 21348 41359
rect 21228 41322 21348 41325
rect 22528 41359 22648 41362
rect 22528 41325 22573 41359
rect 22607 41325 22648 41359
rect 22528 41322 22648 41325
rect 23828 41359 23948 41362
rect 23828 41325 23873 41359
rect 23907 41325 23948 41359
rect 23828 41322 23948 41325
rect 25128 41359 25248 41362
rect 25128 41325 25173 41359
rect 25207 41325 25248 41359
rect 25128 41322 25248 41325
rect 26428 41359 26548 41362
rect 26428 41325 26473 41359
rect 26507 41325 26548 41359
rect 26428 41322 26548 41325
rect 27728 41359 27848 41362
rect 27728 41325 27773 41359
rect 27807 41325 27848 41359
rect 27728 41322 27848 41325
rect 29028 41359 29148 41362
rect 29028 41325 29073 41359
rect 29107 41325 29148 41359
rect 29028 41322 29148 41325
rect 30328 41359 30448 41362
rect 30328 41325 30373 41359
rect 30407 41325 30448 41359
rect 30328 41322 30448 41325
rect 31628 41359 31748 41362
rect 31628 41325 31673 41359
rect 31707 41325 31748 41359
rect 31628 41322 31748 41325
rect 32928 41359 33048 41362
rect 32928 41325 32973 41359
rect 33007 41325 33048 41359
rect 32928 41322 33048 41325
rect 34228 41359 34348 41362
rect 34228 41325 34273 41359
rect 34307 41325 34348 41359
rect 34228 41322 34348 41325
rect 35528 41359 35648 41362
rect 35528 41325 35573 41359
rect 35607 41325 35648 41359
rect 35528 41322 35648 41325
rect 36828 41359 36948 41362
rect 36828 41325 36873 41359
rect 36907 41325 36948 41359
rect 36828 41322 36948 41325
rect 38128 41359 38248 41362
rect 38128 41325 38173 41359
rect 38207 41325 38248 41359
rect 38128 41322 38248 41325
rect 39428 41359 39548 41362
rect 39428 41325 39473 41359
rect 39507 41325 39548 41359
rect 39428 41322 39548 41325
rect 40728 41359 40848 41362
rect 40728 41325 40773 41359
rect 40807 41325 40848 41359
rect 40728 41322 40848 41325
rect 14970 41275 14973 41309
rect 15007 41275 15010 41309
rect 14970 41232 15010 41275
rect 30213 37194 31175 37213
rect 30213 37160 30344 37194
rect 30378 37160 30434 37194
rect 30468 37160 30524 37194
rect 30558 37160 30614 37194
rect 30648 37160 30704 37194
rect 30738 37160 30794 37194
rect 30828 37160 30884 37194
rect 30918 37160 30974 37194
rect 31008 37160 31064 37194
rect 31098 37160 31175 37194
rect 30213 37141 31175 37160
rect 30213 37137 30285 37141
rect 30213 37103 30232 37137
rect 30266 37103 30285 37137
rect 30213 37047 30285 37103
rect 31103 37118 31175 37141
rect 31103 37084 31122 37118
rect 31156 37084 31175 37118
rect 30213 37013 30232 37047
rect 30266 37013 30285 37047
rect 30213 36957 30285 37013
rect 30213 36923 30232 36957
rect 30266 36923 30285 36957
rect 30213 36867 30285 36923
rect 30213 36833 30232 36867
rect 30266 36833 30285 36867
rect 30213 36777 30285 36833
rect 30213 36743 30232 36777
rect 30266 36743 30285 36777
rect 30213 36687 30285 36743
rect 30213 36653 30232 36687
rect 30266 36653 30285 36687
rect 30213 36597 30285 36653
rect 30213 36563 30232 36597
rect 30266 36563 30285 36597
rect 30213 36507 30285 36563
rect 30213 36473 30232 36507
rect 30266 36473 30285 36507
rect 30213 36417 30285 36473
rect 30213 36383 30232 36417
rect 30266 36383 30285 36417
rect 31103 37028 31175 37084
rect 31103 36994 31122 37028
rect 31156 36994 31175 37028
rect 31103 36938 31175 36994
rect 31103 36904 31122 36938
rect 31156 36904 31175 36938
rect 31103 36848 31175 36904
rect 31103 36814 31122 36848
rect 31156 36814 31175 36848
rect 31103 36758 31175 36814
rect 31103 36724 31122 36758
rect 31156 36724 31175 36758
rect 31103 36668 31175 36724
rect 31103 36634 31122 36668
rect 31156 36634 31175 36668
rect 31103 36578 31175 36634
rect 31103 36544 31122 36578
rect 31156 36544 31175 36578
rect 31103 36488 31175 36544
rect 31103 36454 31122 36488
rect 31156 36454 31175 36488
rect 31103 36398 31175 36454
rect 30213 36323 30285 36383
rect 31103 36364 31122 36398
rect 31156 36364 31175 36398
rect 31103 36323 31175 36364
rect 30213 36304 31175 36323
rect 30213 36270 30310 36304
rect 30344 36270 30400 36304
rect 30434 36270 30490 36304
rect 30524 36270 30580 36304
rect 30614 36270 30670 36304
rect 30704 36270 30760 36304
rect 30794 36270 30850 36304
rect 30884 36270 30940 36304
rect 30974 36270 31030 36304
rect 31064 36270 31175 36304
rect 30213 36251 31175 36270
rect 31553 37194 32515 37213
rect 31553 37160 31684 37194
rect 31718 37160 31774 37194
rect 31808 37160 31864 37194
rect 31898 37160 31954 37194
rect 31988 37160 32044 37194
rect 32078 37160 32134 37194
rect 32168 37160 32224 37194
rect 32258 37160 32314 37194
rect 32348 37160 32404 37194
rect 32438 37160 32515 37194
rect 31553 37141 32515 37160
rect 31553 37137 31625 37141
rect 31553 37103 31572 37137
rect 31606 37103 31625 37137
rect 31553 37047 31625 37103
rect 32443 37118 32515 37141
rect 32443 37084 32462 37118
rect 32496 37084 32515 37118
rect 31553 37013 31572 37047
rect 31606 37013 31625 37047
rect 31553 36957 31625 37013
rect 31553 36923 31572 36957
rect 31606 36923 31625 36957
rect 31553 36867 31625 36923
rect 31553 36833 31572 36867
rect 31606 36833 31625 36867
rect 31553 36777 31625 36833
rect 31553 36743 31572 36777
rect 31606 36743 31625 36777
rect 31553 36687 31625 36743
rect 31553 36653 31572 36687
rect 31606 36653 31625 36687
rect 31553 36597 31625 36653
rect 31553 36563 31572 36597
rect 31606 36563 31625 36597
rect 31553 36507 31625 36563
rect 31553 36473 31572 36507
rect 31606 36473 31625 36507
rect 31553 36417 31625 36473
rect 31553 36383 31572 36417
rect 31606 36383 31625 36417
rect 32443 37028 32515 37084
rect 32443 36994 32462 37028
rect 32496 36994 32515 37028
rect 32443 36938 32515 36994
rect 32443 36904 32462 36938
rect 32496 36904 32515 36938
rect 32443 36848 32515 36904
rect 32443 36814 32462 36848
rect 32496 36814 32515 36848
rect 32443 36758 32515 36814
rect 32443 36724 32462 36758
rect 32496 36724 32515 36758
rect 32443 36668 32515 36724
rect 32443 36634 32462 36668
rect 32496 36634 32515 36668
rect 32443 36578 32515 36634
rect 32443 36544 32462 36578
rect 32496 36544 32515 36578
rect 32443 36488 32515 36544
rect 32443 36454 32462 36488
rect 32496 36454 32515 36488
rect 32443 36398 32515 36454
rect 31553 36323 31625 36383
rect 32443 36364 32462 36398
rect 32496 36364 32515 36398
rect 32443 36323 32515 36364
rect 31553 36304 32515 36323
rect 31553 36270 31650 36304
rect 31684 36270 31740 36304
rect 31774 36270 31830 36304
rect 31864 36270 31920 36304
rect 31954 36270 32010 36304
rect 32044 36270 32100 36304
rect 32134 36270 32190 36304
rect 32224 36270 32280 36304
rect 32314 36270 32370 36304
rect 32404 36270 32515 36304
rect 31553 36251 32515 36270
rect 32893 37194 33855 37213
rect 32893 37160 33024 37194
rect 33058 37160 33114 37194
rect 33148 37160 33204 37194
rect 33238 37160 33294 37194
rect 33328 37160 33384 37194
rect 33418 37160 33474 37194
rect 33508 37160 33564 37194
rect 33598 37160 33654 37194
rect 33688 37160 33744 37194
rect 33778 37160 33855 37194
rect 32893 37141 33855 37160
rect 32893 37137 32965 37141
rect 32893 37103 32912 37137
rect 32946 37103 32965 37137
rect 32893 37047 32965 37103
rect 33783 37118 33855 37141
rect 33783 37084 33802 37118
rect 33836 37084 33855 37118
rect 32893 37013 32912 37047
rect 32946 37013 32965 37047
rect 32893 36957 32965 37013
rect 32893 36923 32912 36957
rect 32946 36923 32965 36957
rect 32893 36867 32965 36923
rect 32893 36833 32912 36867
rect 32946 36833 32965 36867
rect 32893 36777 32965 36833
rect 32893 36743 32912 36777
rect 32946 36743 32965 36777
rect 32893 36687 32965 36743
rect 32893 36653 32912 36687
rect 32946 36653 32965 36687
rect 32893 36597 32965 36653
rect 32893 36563 32912 36597
rect 32946 36563 32965 36597
rect 32893 36507 32965 36563
rect 32893 36473 32912 36507
rect 32946 36473 32965 36507
rect 32893 36417 32965 36473
rect 32893 36383 32912 36417
rect 32946 36383 32965 36417
rect 33783 37028 33855 37084
rect 33783 36994 33802 37028
rect 33836 36994 33855 37028
rect 33783 36938 33855 36994
rect 33783 36904 33802 36938
rect 33836 36904 33855 36938
rect 33783 36848 33855 36904
rect 33783 36814 33802 36848
rect 33836 36814 33855 36848
rect 33783 36758 33855 36814
rect 33783 36724 33802 36758
rect 33836 36724 33855 36758
rect 33783 36668 33855 36724
rect 33783 36634 33802 36668
rect 33836 36634 33855 36668
rect 33783 36578 33855 36634
rect 33783 36544 33802 36578
rect 33836 36544 33855 36578
rect 33783 36488 33855 36544
rect 33783 36454 33802 36488
rect 33836 36454 33855 36488
rect 33783 36398 33855 36454
rect 32893 36323 32965 36383
rect 33783 36364 33802 36398
rect 33836 36364 33855 36398
rect 33783 36323 33855 36364
rect 32893 36304 33855 36323
rect 32893 36270 32990 36304
rect 33024 36270 33080 36304
rect 33114 36270 33170 36304
rect 33204 36270 33260 36304
rect 33294 36270 33350 36304
rect 33384 36270 33440 36304
rect 33474 36270 33530 36304
rect 33564 36270 33620 36304
rect 33654 36270 33710 36304
rect 33744 36270 33855 36304
rect 32893 36251 33855 36270
rect 34233 37194 35195 37213
rect 34233 37160 34364 37194
rect 34398 37160 34454 37194
rect 34488 37160 34544 37194
rect 34578 37160 34634 37194
rect 34668 37160 34724 37194
rect 34758 37160 34814 37194
rect 34848 37160 34904 37194
rect 34938 37160 34994 37194
rect 35028 37160 35084 37194
rect 35118 37160 35195 37194
rect 34233 37141 35195 37160
rect 34233 37137 34305 37141
rect 34233 37103 34252 37137
rect 34286 37103 34305 37137
rect 34233 37047 34305 37103
rect 35123 37118 35195 37141
rect 35123 37084 35142 37118
rect 35176 37084 35195 37118
rect 34233 37013 34252 37047
rect 34286 37013 34305 37047
rect 34233 36957 34305 37013
rect 34233 36923 34252 36957
rect 34286 36923 34305 36957
rect 34233 36867 34305 36923
rect 34233 36833 34252 36867
rect 34286 36833 34305 36867
rect 34233 36777 34305 36833
rect 34233 36743 34252 36777
rect 34286 36743 34305 36777
rect 34233 36687 34305 36743
rect 34233 36653 34252 36687
rect 34286 36653 34305 36687
rect 34233 36597 34305 36653
rect 34233 36563 34252 36597
rect 34286 36563 34305 36597
rect 34233 36507 34305 36563
rect 34233 36473 34252 36507
rect 34286 36473 34305 36507
rect 34233 36417 34305 36473
rect 34233 36383 34252 36417
rect 34286 36383 34305 36417
rect 35123 37028 35195 37084
rect 35123 36994 35142 37028
rect 35176 36994 35195 37028
rect 35123 36938 35195 36994
rect 35123 36904 35142 36938
rect 35176 36904 35195 36938
rect 35123 36848 35195 36904
rect 35123 36814 35142 36848
rect 35176 36814 35195 36848
rect 35123 36758 35195 36814
rect 35123 36724 35142 36758
rect 35176 36724 35195 36758
rect 35123 36668 35195 36724
rect 35123 36634 35142 36668
rect 35176 36634 35195 36668
rect 35123 36578 35195 36634
rect 35123 36544 35142 36578
rect 35176 36544 35195 36578
rect 35123 36488 35195 36544
rect 35123 36454 35142 36488
rect 35176 36454 35195 36488
rect 35123 36398 35195 36454
rect 34233 36323 34305 36383
rect 35123 36364 35142 36398
rect 35176 36364 35195 36398
rect 35123 36323 35195 36364
rect 34233 36304 35195 36323
rect 34233 36270 34330 36304
rect 34364 36270 34420 36304
rect 34454 36270 34510 36304
rect 34544 36270 34600 36304
rect 34634 36270 34690 36304
rect 34724 36270 34780 36304
rect 34814 36270 34870 36304
rect 34904 36270 34960 36304
rect 34994 36270 35050 36304
rect 35084 36270 35195 36304
rect 34233 36251 35195 36270
rect 35573 37194 36535 37213
rect 35573 37160 35704 37194
rect 35738 37160 35794 37194
rect 35828 37160 35884 37194
rect 35918 37160 35974 37194
rect 36008 37160 36064 37194
rect 36098 37160 36154 37194
rect 36188 37160 36244 37194
rect 36278 37160 36334 37194
rect 36368 37160 36424 37194
rect 36458 37160 36535 37194
rect 35573 37141 36535 37160
rect 35573 37137 35645 37141
rect 35573 37103 35592 37137
rect 35626 37103 35645 37137
rect 35573 37047 35645 37103
rect 36463 37118 36535 37141
rect 36463 37084 36482 37118
rect 36516 37084 36535 37118
rect 35573 37013 35592 37047
rect 35626 37013 35645 37047
rect 35573 36957 35645 37013
rect 35573 36923 35592 36957
rect 35626 36923 35645 36957
rect 35573 36867 35645 36923
rect 35573 36833 35592 36867
rect 35626 36833 35645 36867
rect 35573 36777 35645 36833
rect 35573 36743 35592 36777
rect 35626 36743 35645 36777
rect 35573 36687 35645 36743
rect 35573 36653 35592 36687
rect 35626 36653 35645 36687
rect 35573 36597 35645 36653
rect 35573 36563 35592 36597
rect 35626 36563 35645 36597
rect 35573 36507 35645 36563
rect 35573 36473 35592 36507
rect 35626 36473 35645 36507
rect 35573 36417 35645 36473
rect 35573 36383 35592 36417
rect 35626 36383 35645 36417
rect 36463 37028 36535 37084
rect 36463 36994 36482 37028
rect 36516 36994 36535 37028
rect 36463 36938 36535 36994
rect 36463 36904 36482 36938
rect 36516 36904 36535 36938
rect 36463 36848 36535 36904
rect 36463 36814 36482 36848
rect 36516 36814 36535 36848
rect 36463 36758 36535 36814
rect 36463 36724 36482 36758
rect 36516 36724 36535 36758
rect 36463 36668 36535 36724
rect 36463 36634 36482 36668
rect 36516 36634 36535 36668
rect 36463 36578 36535 36634
rect 36463 36544 36482 36578
rect 36516 36544 36535 36578
rect 36463 36488 36535 36544
rect 36463 36454 36482 36488
rect 36516 36454 36535 36488
rect 36463 36398 36535 36454
rect 35573 36323 35645 36383
rect 36463 36364 36482 36398
rect 36516 36364 36535 36398
rect 36463 36323 36535 36364
rect 35573 36304 36535 36323
rect 35573 36270 35670 36304
rect 35704 36270 35760 36304
rect 35794 36270 35850 36304
rect 35884 36270 35940 36304
rect 35974 36270 36030 36304
rect 36064 36270 36120 36304
rect 36154 36270 36210 36304
rect 36244 36270 36300 36304
rect 36334 36270 36390 36304
rect 36424 36270 36535 36304
rect 35573 36251 36535 36270
rect 36913 37194 37875 37213
rect 36913 37160 37044 37194
rect 37078 37160 37134 37194
rect 37168 37160 37224 37194
rect 37258 37160 37314 37194
rect 37348 37160 37404 37194
rect 37438 37160 37494 37194
rect 37528 37160 37584 37194
rect 37618 37160 37674 37194
rect 37708 37160 37764 37194
rect 37798 37160 37875 37194
rect 36913 37141 37875 37160
rect 36913 37137 36985 37141
rect 36913 37103 36932 37137
rect 36966 37103 36985 37137
rect 36913 37047 36985 37103
rect 37803 37118 37875 37141
rect 37803 37084 37822 37118
rect 37856 37084 37875 37118
rect 36913 37013 36932 37047
rect 36966 37013 36985 37047
rect 36913 36957 36985 37013
rect 36913 36923 36932 36957
rect 36966 36923 36985 36957
rect 36913 36867 36985 36923
rect 36913 36833 36932 36867
rect 36966 36833 36985 36867
rect 36913 36777 36985 36833
rect 36913 36743 36932 36777
rect 36966 36743 36985 36777
rect 36913 36687 36985 36743
rect 36913 36653 36932 36687
rect 36966 36653 36985 36687
rect 36913 36597 36985 36653
rect 36913 36563 36932 36597
rect 36966 36563 36985 36597
rect 36913 36507 36985 36563
rect 36913 36473 36932 36507
rect 36966 36473 36985 36507
rect 36913 36417 36985 36473
rect 36913 36383 36932 36417
rect 36966 36383 36985 36417
rect 37803 37028 37875 37084
rect 37803 36994 37822 37028
rect 37856 36994 37875 37028
rect 37803 36938 37875 36994
rect 37803 36904 37822 36938
rect 37856 36904 37875 36938
rect 37803 36848 37875 36904
rect 37803 36814 37822 36848
rect 37856 36814 37875 36848
rect 37803 36758 37875 36814
rect 37803 36724 37822 36758
rect 37856 36724 37875 36758
rect 37803 36668 37875 36724
rect 37803 36634 37822 36668
rect 37856 36634 37875 36668
rect 37803 36578 37875 36634
rect 37803 36544 37822 36578
rect 37856 36544 37875 36578
rect 37803 36488 37875 36544
rect 37803 36454 37822 36488
rect 37856 36454 37875 36488
rect 37803 36398 37875 36454
rect 36913 36323 36985 36383
rect 37803 36364 37822 36398
rect 37856 36364 37875 36398
rect 37803 36323 37875 36364
rect 36913 36304 37875 36323
rect 36913 36270 37010 36304
rect 37044 36270 37100 36304
rect 37134 36270 37190 36304
rect 37224 36270 37280 36304
rect 37314 36270 37370 36304
rect 37404 36270 37460 36304
rect 37494 36270 37550 36304
rect 37584 36270 37640 36304
rect 37674 36270 37730 36304
rect 37764 36270 37875 36304
rect 36913 36251 37875 36270
rect 38253 37194 39215 37213
rect 38253 37160 38384 37194
rect 38418 37160 38474 37194
rect 38508 37160 38564 37194
rect 38598 37160 38654 37194
rect 38688 37160 38744 37194
rect 38778 37160 38834 37194
rect 38868 37160 38924 37194
rect 38958 37160 39014 37194
rect 39048 37160 39104 37194
rect 39138 37160 39215 37194
rect 38253 37141 39215 37160
rect 38253 37137 38325 37141
rect 38253 37103 38272 37137
rect 38306 37103 38325 37137
rect 38253 37047 38325 37103
rect 39143 37118 39215 37141
rect 39143 37084 39162 37118
rect 39196 37084 39215 37118
rect 38253 37013 38272 37047
rect 38306 37013 38325 37047
rect 38253 36957 38325 37013
rect 38253 36923 38272 36957
rect 38306 36923 38325 36957
rect 38253 36867 38325 36923
rect 38253 36833 38272 36867
rect 38306 36833 38325 36867
rect 38253 36777 38325 36833
rect 38253 36743 38272 36777
rect 38306 36743 38325 36777
rect 38253 36687 38325 36743
rect 38253 36653 38272 36687
rect 38306 36653 38325 36687
rect 38253 36597 38325 36653
rect 38253 36563 38272 36597
rect 38306 36563 38325 36597
rect 38253 36507 38325 36563
rect 38253 36473 38272 36507
rect 38306 36473 38325 36507
rect 38253 36417 38325 36473
rect 38253 36383 38272 36417
rect 38306 36383 38325 36417
rect 39143 37028 39215 37084
rect 39143 36994 39162 37028
rect 39196 36994 39215 37028
rect 39143 36938 39215 36994
rect 39143 36904 39162 36938
rect 39196 36904 39215 36938
rect 39143 36848 39215 36904
rect 39143 36814 39162 36848
rect 39196 36814 39215 36848
rect 39143 36758 39215 36814
rect 39143 36724 39162 36758
rect 39196 36724 39215 36758
rect 39143 36668 39215 36724
rect 39143 36634 39162 36668
rect 39196 36634 39215 36668
rect 39143 36578 39215 36634
rect 39143 36544 39162 36578
rect 39196 36544 39215 36578
rect 39143 36488 39215 36544
rect 39143 36454 39162 36488
rect 39196 36454 39215 36488
rect 39143 36398 39215 36454
rect 38253 36323 38325 36383
rect 39143 36364 39162 36398
rect 39196 36364 39215 36398
rect 39143 36323 39215 36364
rect 38253 36304 39215 36323
rect 38253 36270 38350 36304
rect 38384 36270 38440 36304
rect 38474 36270 38530 36304
rect 38564 36270 38620 36304
rect 38654 36270 38710 36304
rect 38744 36270 38800 36304
rect 38834 36270 38890 36304
rect 38924 36270 38980 36304
rect 39014 36270 39070 36304
rect 39104 36270 39215 36304
rect 38253 36251 39215 36270
rect 15146 33839 15266 33842
rect 14088 33789 14128 33832
rect 15146 33805 15191 33839
rect 15225 33805 15266 33839
rect 15146 33802 15266 33805
rect 16446 33839 16566 33842
rect 16446 33805 16491 33839
rect 16525 33805 16566 33839
rect 16446 33802 16566 33805
rect 17746 33839 17866 33842
rect 17746 33805 17791 33839
rect 17825 33805 17866 33839
rect 17746 33802 17866 33805
rect 19046 33839 19166 33842
rect 19046 33805 19091 33839
rect 19125 33805 19166 33839
rect 19046 33802 19166 33805
rect 20346 33839 20466 33842
rect 20346 33805 20391 33839
rect 20425 33805 20466 33839
rect 20346 33802 20466 33805
rect 21646 33839 21766 33842
rect 21646 33805 21691 33839
rect 21725 33805 21766 33839
rect 21646 33802 21766 33805
rect 22946 33839 23066 33842
rect 22946 33805 22991 33839
rect 23025 33805 23066 33839
rect 22946 33802 23066 33805
rect 24246 33839 24366 33842
rect 24246 33805 24291 33839
rect 24325 33805 24366 33839
rect 24246 33802 24366 33805
rect 25546 33839 25666 33842
rect 25546 33805 25591 33839
rect 25625 33805 25666 33839
rect 25546 33802 25666 33805
rect 26846 33839 26966 33842
rect 26846 33805 26891 33839
rect 26925 33805 26966 33839
rect 26846 33802 26966 33805
rect 28146 33839 28266 33842
rect 28146 33805 28191 33839
rect 28225 33805 28266 33839
rect 28146 33802 28266 33805
rect 29446 33839 29566 33842
rect 29446 33805 29491 33839
rect 29525 33805 29566 33839
rect 29446 33802 29566 33805
rect 30746 33839 30866 33842
rect 30746 33805 30791 33839
rect 30825 33805 30866 33839
rect 30746 33802 30866 33805
rect 32046 33839 32166 33842
rect 32046 33805 32091 33839
rect 32125 33805 32166 33839
rect 32046 33802 32166 33805
rect 33346 33839 33466 33842
rect 33346 33805 33391 33839
rect 33425 33805 33466 33839
rect 33346 33802 33466 33805
rect 34646 33839 34766 33842
rect 34646 33805 34691 33839
rect 34725 33805 34766 33839
rect 34646 33802 34766 33805
rect 35946 33839 36066 33842
rect 35946 33805 35991 33839
rect 36025 33805 36066 33839
rect 35946 33802 36066 33805
rect 37246 33839 37366 33842
rect 37246 33805 37291 33839
rect 37325 33805 37366 33839
rect 37246 33802 37366 33805
rect 38546 33839 38666 33842
rect 38546 33805 38591 33839
rect 38625 33805 38666 33839
rect 38546 33802 38666 33805
rect 39846 33839 39966 33842
rect 39846 33805 39891 33839
rect 39925 33805 39966 33839
rect 39846 33802 39966 33805
rect 14088 33755 14091 33789
rect 14125 33755 14128 33789
rect 14088 33712 14128 33755
rect 7012 30079 7132 30082
rect 5954 30029 5994 30072
rect 7012 30045 7057 30079
rect 7091 30045 7132 30079
rect 7012 30042 7132 30045
rect 8312 30079 8432 30082
rect 8312 30045 8357 30079
rect 8391 30045 8432 30079
rect 8312 30042 8432 30045
rect 9612 30079 9732 30082
rect 9612 30045 9657 30079
rect 9691 30045 9732 30079
rect 9612 30042 9732 30045
rect 10912 30079 11032 30082
rect 10912 30045 10957 30079
rect 10991 30045 11032 30079
rect 10912 30042 11032 30045
rect 12212 30079 12332 30082
rect 12212 30045 12257 30079
rect 12291 30045 12332 30079
rect 12212 30042 12332 30045
rect 13512 30079 13632 30082
rect 13512 30045 13557 30079
rect 13591 30045 13632 30079
rect 13512 30042 13632 30045
rect 14812 30079 14932 30082
rect 14812 30045 14857 30079
rect 14891 30045 14932 30079
rect 14812 30042 14932 30045
rect 16112 30079 16232 30082
rect 16112 30045 16157 30079
rect 16191 30045 16232 30079
rect 16112 30042 16232 30045
rect 17412 30079 17532 30082
rect 17412 30045 17457 30079
rect 17491 30045 17532 30079
rect 17412 30042 17532 30045
rect 18712 30079 18832 30082
rect 18712 30045 18757 30079
rect 18791 30045 18832 30079
rect 18712 30042 18832 30045
rect 20012 30079 20132 30082
rect 20012 30045 20057 30079
rect 20091 30045 20132 30079
rect 20012 30042 20132 30045
rect 21312 30079 21432 30082
rect 21312 30045 21357 30079
rect 21391 30045 21432 30079
rect 21312 30042 21432 30045
rect 22612 30079 22732 30082
rect 22612 30045 22657 30079
rect 22691 30045 22732 30079
rect 22612 30042 22732 30045
rect 23912 30079 24032 30082
rect 23912 30045 23957 30079
rect 23991 30045 24032 30079
rect 23912 30042 24032 30045
rect 25212 30079 25332 30082
rect 25212 30045 25257 30079
rect 25291 30045 25332 30079
rect 25212 30042 25332 30045
rect 26512 30079 26632 30082
rect 26512 30045 26557 30079
rect 26591 30045 26632 30079
rect 26512 30042 26632 30045
rect 27812 30079 27932 30082
rect 27812 30045 27857 30079
rect 27891 30045 27932 30079
rect 27812 30042 27932 30045
rect 29112 30079 29232 30082
rect 29112 30045 29157 30079
rect 29191 30045 29232 30079
rect 29112 30042 29232 30045
rect 30412 30079 30532 30082
rect 30412 30045 30457 30079
rect 30491 30045 30532 30079
rect 30412 30042 30532 30045
rect 31712 30079 31832 30082
rect 31712 30045 31757 30079
rect 31791 30045 31832 30079
rect 35040 30079 35160 30082
rect 31712 30042 31832 30045
rect 5954 29995 5957 30029
rect 5991 29995 5994 30029
rect 5954 29952 5994 29995
rect 33982 30029 34022 30072
rect 35040 30045 35085 30079
rect 35119 30045 35160 30079
rect 35040 30042 35160 30045
rect 33982 29995 33985 30029
rect 34019 29995 34022 30029
rect 33982 29952 34022 29995
rect 10540 26319 10660 26322
rect 9482 26269 9522 26312
rect 10540 26285 10585 26319
rect 10619 26285 10660 26319
rect 10540 26282 10660 26285
rect 11840 26319 11960 26322
rect 11840 26285 11885 26319
rect 11919 26285 11960 26319
rect 11840 26282 11960 26285
rect 13140 26319 13260 26322
rect 13140 26285 13185 26319
rect 13219 26285 13260 26319
rect 13140 26282 13260 26285
rect 9482 26235 9485 26269
rect 9519 26235 9522 26269
rect 9482 26192 9522 26235
rect 28449 25914 29411 25933
rect 28449 25880 28580 25914
rect 28614 25880 28670 25914
rect 28704 25880 28760 25914
rect 28794 25880 28850 25914
rect 28884 25880 28940 25914
rect 28974 25880 29030 25914
rect 29064 25880 29120 25914
rect 29154 25880 29210 25914
rect 29244 25880 29300 25914
rect 29334 25880 29411 25914
rect 28449 25861 29411 25880
rect 28449 25857 28521 25861
rect 28449 25823 28468 25857
rect 28502 25823 28521 25857
rect 28449 25767 28521 25823
rect 29339 25838 29411 25861
rect 29339 25804 29358 25838
rect 29392 25804 29411 25838
rect 28449 25733 28468 25767
rect 28502 25733 28521 25767
rect 28449 25677 28521 25733
rect 28449 25643 28468 25677
rect 28502 25643 28521 25677
rect 28449 25587 28521 25643
rect 28449 25553 28468 25587
rect 28502 25553 28521 25587
rect 28449 25497 28521 25553
rect 28449 25463 28468 25497
rect 28502 25463 28521 25497
rect 28449 25407 28521 25463
rect 28449 25373 28468 25407
rect 28502 25373 28521 25407
rect 28449 25317 28521 25373
rect 28449 25283 28468 25317
rect 28502 25283 28521 25317
rect 28449 25227 28521 25283
rect 28449 25193 28468 25227
rect 28502 25193 28521 25227
rect 28449 25137 28521 25193
rect 28449 25103 28468 25137
rect 28502 25103 28521 25137
rect 29339 25748 29411 25804
rect 29339 25714 29358 25748
rect 29392 25714 29411 25748
rect 29339 25658 29411 25714
rect 29339 25624 29358 25658
rect 29392 25624 29411 25658
rect 29339 25568 29411 25624
rect 29339 25534 29358 25568
rect 29392 25534 29411 25568
rect 29339 25478 29411 25534
rect 29339 25444 29358 25478
rect 29392 25444 29411 25478
rect 29339 25388 29411 25444
rect 29339 25354 29358 25388
rect 29392 25354 29411 25388
rect 29339 25298 29411 25354
rect 29339 25264 29358 25298
rect 29392 25264 29411 25298
rect 29339 25208 29411 25264
rect 29339 25174 29358 25208
rect 29392 25174 29411 25208
rect 29339 25118 29411 25174
rect 28449 25043 28521 25103
rect 29339 25084 29358 25118
rect 29392 25084 29411 25118
rect 29339 25043 29411 25084
rect 28449 25024 29411 25043
rect 28449 24990 28546 25024
rect 28580 24990 28636 25024
rect 28670 24990 28726 25024
rect 28760 24990 28816 25024
rect 28850 24990 28906 25024
rect 28940 24990 28996 25024
rect 29030 24990 29086 25024
rect 29120 24990 29176 25024
rect 29210 24990 29266 25024
rect 29300 24990 29411 25024
rect 28449 24971 29411 24990
rect 29789 25914 30751 25933
rect 29789 25880 29920 25914
rect 29954 25880 30010 25914
rect 30044 25880 30100 25914
rect 30134 25880 30190 25914
rect 30224 25880 30280 25914
rect 30314 25880 30370 25914
rect 30404 25880 30460 25914
rect 30494 25880 30550 25914
rect 30584 25880 30640 25914
rect 30674 25880 30751 25914
rect 29789 25861 30751 25880
rect 29789 25857 29861 25861
rect 29789 25823 29808 25857
rect 29842 25823 29861 25857
rect 29789 25767 29861 25823
rect 30679 25838 30751 25861
rect 30679 25804 30698 25838
rect 30732 25804 30751 25838
rect 29789 25733 29808 25767
rect 29842 25733 29861 25767
rect 29789 25677 29861 25733
rect 29789 25643 29808 25677
rect 29842 25643 29861 25677
rect 29789 25587 29861 25643
rect 29789 25553 29808 25587
rect 29842 25553 29861 25587
rect 29789 25497 29861 25553
rect 29789 25463 29808 25497
rect 29842 25463 29861 25497
rect 29789 25407 29861 25463
rect 29789 25373 29808 25407
rect 29842 25373 29861 25407
rect 29789 25317 29861 25373
rect 29789 25283 29808 25317
rect 29842 25283 29861 25317
rect 29789 25227 29861 25283
rect 29789 25193 29808 25227
rect 29842 25193 29861 25227
rect 29789 25137 29861 25193
rect 29789 25103 29808 25137
rect 29842 25103 29861 25137
rect 30679 25748 30751 25804
rect 30679 25714 30698 25748
rect 30732 25714 30751 25748
rect 30679 25658 30751 25714
rect 30679 25624 30698 25658
rect 30732 25624 30751 25658
rect 30679 25568 30751 25624
rect 30679 25534 30698 25568
rect 30732 25534 30751 25568
rect 30679 25478 30751 25534
rect 30679 25444 30698 25478
rect 30732 25444 30751 25478
rect 30679 25388 30751 25444
rect 30679 25354 30698 25388
rect 30732 25354 30751 25388
rect 30679 25298 30751 25354
rect 30679 25264 30698 25298
rect 30732 25264 30751 25298
rect 30679 25208 30751 25264
rect 30679 25174 30698 25208
rect 30732 25174 30751 25208
rect 30679 25118 30751 25174
rect 29789 25043 29861 25103
rect 30679 25084 30698 25118
rect 30732 25084 30751 25118
rect 30679 25043 30751 25084
rect 29789 25024 30751 25043
rect 29789 24990 29886 25024
rect 29920 24990 29976 25024
rect 30010 24990 30066 25024
rect 30100 24990 30156 25024
rect 30190 24990 30246 25024
rect 30280 24990 30336 25024
rect 30370 24990 30426 25024
rect 30460 24990 30516 25024
rect 30550 24990 30606 25024
rect 30640 24990 30751 25024
rect 29789 24971 30751 24990
rect 31129 25914 32091 25933
rect 31129 25880 31260 25914
rect 31294 25880 31350 25914
rect 31384 25880 31440 25914
rect 31474 25880 31530 25914
rect 31564 25880 31620 25914
rect 31654 25880 31710 25914
rect 31744 25880 31800 25914
rect 31834 25880 31890 25914
rect 31924 25880 31980 25914
rect 32014 25880 32091 25914
rect 31129 25861 32091 25880
rect 31129 25857 31201 25861
rect 31129 25823 31148 25857
rect 31182 25823 31201 25857
rect 31129 25767 31201 25823
rect 32019 25838 32091 25861
rect 32019 25804 32038 25838
rect 32072 25804 32091 25838
rect 31129 25733 31148 25767
rect 31182 25733 31201 25767
rect 31129 25677 31201 25733
rect 31129 25643 31148 25677
rect 31182 25643 31201 25677
rect 31129 25587 31201 25643
rect 31129 25553 31148 25587
rect 31182 25553 31201 25587
rect 31129 25497 31201 25553
rect 31129 25463 31148 25497
rect 31182 25463 31201 25497
rect 31129 25407 31201 25463
rect 31129 25373 31148 25407
rect 31182 25373 31201 25407
rect 31129 25317 31201 25373
rect 31129 25283 31148 25317
rect 31182 25283 31201 25317
rect 31129 25227 31201 25283
rect 31129 25193 31148 25227
rect 31182 25193 31201 25227
rect 31129 25137 31201 25193
rect 31129 25103 31148 25137
rect 31182 25103 31201 25137
rect 32019 25748 32091 25804
rect 32019 25714 32038 25748
rect 32072 25714 32091 25748
rect 32019 25658 32091 25714
rect 32019 25624 32038 25658
rect 32072 25624 32091 25658
rect 32019 25568 32091 25624
rect 32019 25534 32038 25568
rect 32072 25534 32091 25568
rect 32019 25478 32091 25534
rect 32019 25444 32038 25478
rect 32072 25444 32091 25478
rect 32019 25388 32091 25444
rect 32019 25354 32038 25388
rect 32072 25354 32091 25388
rect 32019 25298 32091 25354
rect 32019 25264 32038 25298
rect 32072 25264 32091 25298
rect 32019 25208 32091 25264
rect 32019 25174 32038 25208
rect 32072 25174 32091 25208
rect 32019 25118 32091 25174
rect 31129 25043 31201 25103
rect 32019 25084 32038 25118
rect 32072 25084 32091 25118
rect 32019 25043 32091 25084
rect 31129 25024 32091 25043
rect 31129 24990 31226 25024
rect 31260 24990 31316 25024
rect 31350 24990 31406 25024
rect 31440 24990 31496 25024
rect 31530 24990 31586 25024
rect 31620 24990 31676 25024
rect 31710 24990 31766 25024
rect 31800 24990 31856 25024
rect 31890 24990 31946 25024
rect 31980 24990 32091 25024
rect 31129 24971 32091 24990
rect 32469 25914 33431 25933
rect 32469 25880 32600 25914
rect 32634 25880 32690 25914
rect 32724 25880 32780 25914
rect 32814 25880 32870 25914
rect 32904 25880 32960 25914
rect 32994 25880 33050 25914
rect 33084 25880 33140 25914
rect 33174 25880 33230 25914
rect 33264 25880 33320 25914
rect 33354 25880 33431 25914
rect 32469 25861 33431 25880
rect 32469 25857 32541 25861
rect 32469 25823 32488 25857
rect 32522 25823 32541 25857
rect 32469 25767 32541 25823
rect 33359 25838 33431 25861
rect 33359 25804 33378 25838
rect 33412 25804 33431 25838
rect 32469 25733 32488 25767
rect 32522 25733 32541 25767
rect 32469 25677 32541 25733
rect 32469 25643 32488 25677
rect 32522 25643 32541 25677
rect 32469 25587 32541 25643
rect 32469 25553 32488 25587
rect 32522 25553 32541 25587
rect 32469 25497 32541 25553
rect 32469 25463 32488 25497
rect 32522 25463 32541 25497
rect 32469 25407 32541 25463
rect 32469 25373 32488 25407
rect 32522 25373 32541 25407
rect 32469 25317 32541 25373
rect 32469 25283 32488 25317
rect 32522 25283 32541 25317
rect 32469 25227 32541 25283
rect 32469 25193 32488 25227
rect 32522 25193 32541 25227
rect 32469 25137 32541 25193
rect 32469 25103 32488 25137
rect 32522 25103 32541 25137
rect 33359 25748 33431 25804
rect 33359 25714 33378 25748
rect 33412 25714 33431 25748
rect 33359 25658 33431 25714
rect 33359 25624 33378 25658
rect 33412 25624 33431 25658
rect 33359 25568 33431 25624
rect 33359 25534 33378 25568
rect 33412 25534 33431 25568
rect 33359 25478 33431 25534
rect 33359 25444 33378 25478
rect 33412 25444 33431 25478
rect 33359 25388 33431 25444
rect 33359 25354 33378 25388
rect 33412 25354 33431 25388
rect 33359 25298 33431 25354
rect 33359 25264 33378 25298
rect 33412 25264 33431 25298
rect 33359 25208 33431 25264
rect 33359 25174 33378 25208
rect 33412 25174 33431 25208
rect 33359 25118 33431 25174
rect 32469 25043 32541 25103
rect 33359 25084 33378 25118
rect 33412 25084 33431 25118
rect 33359 25043 33431 25084
rect 32469 25024 33431 25043
rect 32469 24990 32566 25024
rect 32600 24990 32656 25024
rect 32690 24990 32746 25024
rect 32780 24990 32836 25024
rect 32870 24990 32926 25024
rect 32960 24990 33016 25024
rect 33050 24990 33106 25024
rect 33140 24990 33196 25024
rect 33230 24990 33286 25024
rect 33320 24990 33431 25024
rect 32469 24971 33431 24990
rect 33809 25914 34771 25933
rect 33809 25880 33940 25914
rect 33974 25880 34030 25914
rect 34064 25880 34120 25914
rect 34154 25880 34210 25914
rect 34244 25880 34300 25914
rect 34334 25880 34390 25914
rect 34424 25880 34480 25914
rect 34514 25880 34570 25914
rect 34604 25880 34660 25914
rect 34694 25880 34771 25914
rect 33809 25861 34771 25880
rect 33809 25857 33881 25861
rect 33809 25823 33828 25857
rect 33862 25823 33881 25857
rect 33809 25767 33881 25823
rect 34699 25838 34771 25861
rect 34699 25804 34718 25838
rect 34752 25804 34771 25838
rect 33809 25733 33828 25767
rect 33862 25733 33881 25767
rect 33809 25677 33881 25733
rect 33809 25643 33828 25677
rect 33862 25643 33881 25677
rect 33809 25587 33881 25643
rect 33809 25553 33828 25587
rect 33862 25553 33881 25587
rect 33809 25497 33881 25553
rect 33809 25463 33828 25497
rect 33862 25463 33881 25497
rect 33809 25407 33881 25463
rect 33809 25373 33828 25407
rect 33862 25373 33881 25407
rect 33809 25317 33881 25373
rect 33809 25283 33828 25317
rect 33862 25283 33881 25317
rect 33809 25227 33881 25283
rect 33809 25193 33828 25227
rect 33862 25193 33881 25227
rect 33809 25137 33881 25193
rect 33809 25103 33828 25137
rect 33862 25103 33881 25137
rect 34699 25748 34771 25804
rect 34699 25714 34718 25748
rect 34752 25714 34771 25748
rect 34699 25658 34771 25714
rect 34699 25624 34718 25658
rect 34752 25624 34771 25658
rect 34699 25568 34771 25624
rect 34699 25534 34718 25568
rect 34752 25534 34771 25568
rect 34699 25478 34771 25534
rect 34699 25444 34718 25478
rect 34752 25444 34771 25478
rect 34699 25388 34771 25444
rect 34699 25354 34718 25388
rect 34752 25354 34771 25388
rect 34699 25298 34771 25354
rect 34699 25264 34718 25298
rect 34752 25264 34771 25298
rect 34699 25208 34771 25264
rect 34699 25174 34718 25208
rect 34752 25174 34771 25208
rect 34699 25118 34771 25174
rect 33809 25043 33881 25103
rect 34699 25084 34718 25118
rect 34752 25084 34771 25118
rect 34699 25043 34771 25084
rect 33809 25024 34771 25043
rect 33809 24990 33906 25024
rect 33940 24990 33996 25024
rect 34030 24990 34086 25024
rect 34120 24990 34176 25024
rect 34210 24990 34266 25024
rect 34300 24990 34356 25024
rect 34390 24990 34446 25024
rect 34480 24990 34536 25024
rect 34570 24990 34626 25024
rect 34660 24990 34771 25024
rect 33809 24971 34771 24990
rect 35149 25914 36111 25933
rect 35149 25880 35280 25914
rect 35314 25880 35370 25914
rect 35404 25880 35460 25914
rect 35494 25880 35550 25914
rect 35584 25880 35640 25914
rect 35674 25880 35730 25914
rect 35764 25880 35820 25914
rect 35854 25880 35910 25914
rect 35944 25880 36000 25914
rect 36034 25880 36111 25914
rect 35149 25861 36111 25880
rect 35149 25857 35221 25861
rect 35149 25823 35168 25857
rect 35202 25823 35221 25857
rect 35149 25767 35221 25823
rect 36039 25838 36111 25861
rect 36039 25804 36058 25838
rect 36092 25804 36111 25838
rect 35149 25733 35168 25767
rect 35202 25733 35221 25767
rect 35149 25677 35221 25733
rect 35149 25643 35168 25677
rect 35202 25643 35221 25677
rect 35149 25587 35221 25643
rect 35149 25553 35168 25587
rect 35202 25553 35221 25587
rect 35149 25497 35221 25553
rect 35149 25463 35168 25497
rect 35202 25463 35221 25497
rect 35149 25407 35221 25463
rect 35149 25373 35168 25407
rect 35202 25373 35221 25407
rect 35149 25317 35221 25373
rect 35149 25283 35168 25317
rect 35202 25283 35221 25317
rect 35149 25227 35221 25283
rect 35149 25193 35168 25227
rect 35202 25193 35221 25227
rect 35149 25137 35221 25193
rect 35149 25103 35168 25137
rect 35202 25103 35221 25137
rect 36039 25748 36111 25804
rect 36039 25714 36058 25748
rect 36092 25714 36111 25748
rect 36039 25658 36111 25714
rect 36039 25624 36058 25658
rect 36092 25624 36111 25658
rect 36039 25568 36111 25624
rect 36039 25534 36058 25568
rect 36092 25534 36111 25568
rect 36039 25478 36111 25534
rect 36039 25444 36058 25478
rect 36092 25444 36111 25478
rect 36039 25388 36111 25444
rect 36039 25354 36058 25388
rect 36092 25354 36111 25388
rect 36039 25298 36111 25354
rect 36039 25264 36058 25298
rect 36092 25264 36111 25298
rect 36039 25208 36111 25264
rect 36039 25174 36058 25208
rect 36092 25174 36111 25208
rect 36039 25118 36111 25174
rect 35149 25043 35221 25103
rect 36039 25084 36058 25118
rect 36092 25084 36111 25118
rect 36039 25043 36111 25084
rect 35149 25024 36111 25043
rect 35149 24990 35246 25024
rect 35280 24990 35336 25024
rect 35370 24990 35426 25024
rect 35460 24990 35516 25024
rect 35550 24990 35606 25024
rect 35640 24990 35696 25024
rect 35730 24990 35786 25024
rect 35820 24990 35876 25024
rect 35910 24990 35966 25024
rect 36000 24990 36111 25024
rect 35149 24971 36111 24990
rect 36489 25914 37451 25933
rect 36489 25880 36620 25914
rect 36654 25880 36710 25914
rect 36744 25880 36800 25914
rect 36834 25880 36890 25914
rect 36924 25880 36980 25914
rect 37014 25880 37070 25914
rect 37104 25880 37160 25914
rect 37194 25880 37250 25914
rect 37284 25880 37340 25914
rect 37374 25880 37451 25914
rect 36489 25861 37451 25880
rect 36489 25857 36561 25861
rect 36489 25823 36508 25857
rect 36542 25823 36561 25857
rect 36489 25767 36561 25823
rect 37379 25838 37451 25861
rect 37379 25804 37398 25838
rect 37432 25804 37451 25838
rect 36489 25733 36508 25767
rect 36542 25733 36561 25767
rect 36489 25677 36561 25733
rect 36489 25643 36508 25677
rect 36542 25643 36561 25677
rect 36489 25587 36561 25643
rect 36489 25553 36508 25587
rect 36542 25553 36561 25587
rect 36489 25497 36561 25553
rect 36489 25463 36508 25497
rect 36542 25463 36561 25497
rect 36489 25407 36561 25463
rect 36489 25373 36508 25407
rect 36542 25373 36561 25407
rect 36489 25317 36561 25373
rect 36489 25283 36508 25317
rect 36542 25283 36561 25317
rect 36489 25227 36561 25283
rect 36489 25193 36508 25227
rect 36542 25193 36561 25227
rect 36489 25137 36561 25193
rect 36489 25103 36508 25137
rect 36542 25103 36561 25137
rect 37379 25748 37451 25804
rect 37379 25714 37398 25748
rect 37432 25714 37451 25748
rect 37379 25658 37451 25714
rect 37379 25624 37398 25658
rect 37432 25624 37451 25658
rect 37379 25568 37451 25624
rect 37379 25534 37398 25568
rect 37432 25534 37451 25568
rect 37379 25478 37451 25534
rect 37379 25444 37398 25478
rect 37432 25444 37451 25478
rect 37379 25388 37451 25444
rect 37379 25354 37398 25388
rect 37432 25354 37451 25388
rect 37379 25298 37451 25354
rect 37379 25264 37398 25298
rect 37432 25264 37451 25298
rect 37379 25208 37451 25264
rect 37379 25174 37398 25208
rect 37432 25174 37451 25208
rect 37379 25118 37451 25174
rect 36489 25043 36561 25103
rect 37379 25084 37398 25118
rect 37432 25084 37451 25118
rect 37379 25043 37451 25084
rect 36489 25024 37451 25043
rect 36489 24990 36586 25024
rect 36620 24990 36676 25024
rect 36710 24990 36766 25024
rect 36800 24990 36856 25024
rect 36890 24990 36946 25024
rect 36980 24990 37036 25024
rect 37070 24990 37126 25024
rect 37160 24990 37216 25024
rect 37250 24990 37306 25024
rect 37340 24990 37451 25024
rect 36489 24971 37451 24990
rect 37829 25914 38791 25933
rect 37829 25880 37960 25914
rect 37994 25880 38050 25914
rect 38084 25880 38140 25914
rect 38174 25880 38230 25914
rect 38264 25880 38320 25914
rect 38354 25880 38410 25914
rect 38444 25880 38500 25914
rect 38534 25880 38590 25914
rect 38624 25880 38680 25914
rect 38714 25880 38791 25914
rect 37829 25861 38791 25880
rect 37829 25857 37901 25861
rect 37829 25823 37848 25857
rect 37882 25823 37901 25857
rect 37829 25767 37901 25823
rect 38719 25838 38791 25861
rect 38719 25804 38738 25838
rect 38772 25804 38791 25838
rect 37829 25733 37848 25767
rect 37882 25733 37901 25767
rect 37829 25677 37901 25733
rect 37829 25643 37848 25677
rect 37882 25643 37901 25677
rect 37829 25587 37901 25643
rect 37829 25553 37848 25587
rect 37882 25553 37901 25587
rect 37829 25497 37901 25553
rect 37829 25463 37848 25497
rect 37882 25463 37901 25497
rect 37829 25407 37901 25463
rect 37829 25373 37848 25407
rect 37882 25373 37901 25407
rect 37829 25317 37901 25373
rect 37829 25283 37848 25317
rect 37882 25283 37901 25317
rect 37829 25227 37901 25283
rect 37829 25193 37848 25227
rect 37882 25193 37901 25227
rect 37829 25137 37901 25193
rect 37829 25103 37848 25137
rect 37882 25103 37901 25137
rect 38719 25748 38791 25804
rect 38719 25714 38738 25748
rect 38772 25714 38791 25748
rect 38719 25658 38791 25714
rect 38719 25624 38738 25658
rect 38772 25624 38791 25658
rect 38719 25568 38791 25624
rect 38719 25534 38738 25568
rect 38772 25534 38791 25568
rect 38719 25478 38791 25534
rect 38719 25444 38738 25478
rect 38772 25444 38791 25478
rect 38719 25388 38791 25444
rect 38719 25354 38738 25388
rect 38772 25354 38791 25388
rect 38719 25298 38791 25354
rect 38719 25264 38738 25298
rect 38772 25264 38791 25298
rect 38719 25208 38791 25264
rect 38719 25174 38738 25208
rect 38772 25174 38791 25208
rect 38719 25118 38791 25174
rect 37829 25043 37901 25103
rect 38719 25084 38738 25118
rect 38772 25084 38791 25118
rect 38719 25043 38791 25084
rect 37829 25024 38791 25043
rect 37829 24990 37926 25024
rect 37960 24990 38016 25024
rect 38050 24990 38106 25024
rect 38140 24990 38196 25024
rect 38230 24990 38286 25024
rect 38320 24990 38376 25024
rect 38410 24990 38466 25024
rect 38500 24990 38556 25024
rect 38590 24990 38646 25024
rect 38680 24990 38791 25024
rect 37829 24971 38791 24990
rect 8678 22559 8798 22562
rect 7620 22509 7660 22552
rect 8678 22525 8723 22559
rect 8757 22525 8798 22559
rect 8678 22522 8798 22525
rect 9978 22559 10098 22562
rect 9978 22525 10023 22559
rect 10057 22525 10098 22559
rect 9978 22522 10098 22525
rect 11278 22559 11398 22562
rect 11278 22525 11323 22559
rect 11357 22525 11398 22559
rect 11278 22522 11398 22525
rect 7620 22475 7623 22509
rect 7657 22475 7660 22509
rect 7620 22432 7660 22475
rect 21197 22154 22159 22173
rect 21197 22120 21328 22154
rect 21362 22120 21418 22154
rect 21452 22120 21508 22154
rect 21542 22120 21598 22154
rect 21632 22120 21688 22154
rect 21722 22120 21778 22154
rect 21812 22120 21868 22154
rect 21902 22120 21958 22154
rect 21992 22120 22048 22154
rect 22082 22120 22159 22154
rect 21197 22101 22159 22120
rect 21197 22097 21269 22101
rect 21197 22063 21216 22097
rect 21250 22063 21269 22097
rect 21197 22007 21269 22063
rect 22087 22078 22159 22101
rect 22087 22044 22106 22078
rect 22140 22044 22159 22078
rect 21197 21973 21216 22007
rect 21250 21973 21269 22007
rect 21197 21917 21269 21973
rect 21197 21883 21216 21917
rect 21250 21883 21269 21917
rect 21197 21827 21269 21883
rect 21197 21793 21216 21827
rect 21250 21793 21269 21827
rect 21197 21737 21269 21793
rect 21197 21703 21216 21737
rect 21250 21703 21269 21737
rect 21197 21647 21269 21703
rect 21197 21613 21216 21647
rect 21250 21613 21269 21647
rect 21197 21557 21269 21613
rect 21197 21523 21216 21557
rect 21250 21523 21269 21557
rect 21197 21467 21269 21523
rect 21197 21433 21216 21467
rect 21250 21433 21269 21467
rect 21197 21377 21269 21433
rect 21197 21343 21216 21377
rect 21250 21343 21269 21377
rect 22087 21988 22159 22044
rect 22087 21954 22106 21988
rect 22140 21954 22159 21988
rect 22087 21898 22159 21954
rect 22087 21864 22106 21898
rect 22140 21864 22159 21898
rect 22087 21808 22159 21864
rect 22087 21774 22106 21808
rect 22140 21774 22159 21808
rect 22087 21718 22159 21774
rect 22087 21684 22106 21718
rect 22140 21684 22159 21718
rect 22087 21628 22159 21684
rect 22087 21594 22106 21628
rect 22140 21594 22159 21628
rect 22087 21538 22159 21594
rect 22087 21504 22106 21538
rect 22140 21504 22159 21538
rect 22087 21448 22159 21504
rect 22087 21414 22106 21448
rect 22140 21414 22159 21448
rect 22087 21358 22159 21414
rect 21197 21283 21269 21343
rect 22087 21324 22106 21358
rect 22140 21324 22159 21358
rect 22087 21283 22159 21324
rect 21197 21264 22159 21283
rect 21197 21230 21294 21264
rect 21328 21230 21384 21264
rect 21418 21230 21474 21264
rect 21508 21230 21564 21264
rect 21598 21230 21654 21264
rect 21688 21230 21744 21264
rect 21778 21230 21834 21264
rect 21868 21230 21924 21264
rect 21958 21230 22014 21264
rect 22048 21230 22159 21264
rect 21197 21211 22159 21230
rect 28449 22154 29411 22173
rect 28449 22120 28580 22154
rect 28614 22120 28670 22154
rect 28704 22120 28760 22154
rect 28794 22120 28850 22154
rect 28884 22120 28940 22154
rect 28974 22120 29030 22154
rect 29064 22120 29120 22154
rect 29154 22120 29210 22154
rect 29244 22120 29300 22154
rect 29334 22120 29411 22154
rect 28449 22101 29411 22120
rect 28449 22097 28521 22101
rect 28449 22063 28468 22097
rect 28502 22063 28521 22097
rect 28449 22007 28521 22063
rect 29339 22078 29411 22101
rect 29339 22044 29358 22078
rect 29392 22044 29411 22078
rect 28449 21973 28468 22007
rect 28502 21973 28521 22007
rect 28449 21917 28521 21973
rect 28449 21883 28468 21917
rect 28502 21883 28521 21917
rect 28449 21827 28521 21883
rect 28449 21793 28468 21827
rect 28502 21793 28521 21827
rect 28449 21737 28521 21793
rect 28449 21703 28468 21737
rect 28502 21703 28521 21737
rect 28449 21647 28521 21703
rect 28449 21613 28468 21647
rect 28502 21613 28521 21647
rect 28449 21557 28521 21613
rect 28449 21523 28468 21557
rect 28502 21523 28521 21557
rect 28449 21467 28521 21523
rect 28449 21433 28468 21467
rect 28502 21433 28521 21467
rect 28449 21377 28521 21433
rect 28449 21343 28468 21377
rect 28502 21343 28521 21377
rect 29339 21988 29411 22044
rect 29339 21954 29358 21988
rect 29392 21954 29411 21988
rect 29339 21898 29411 21954
rect 29339 21864 29358 21898
rect 29392 21864 29411 21898
rect 29339 21808 29411 21864
rect 29339 21774 29358 21808
rect 29392 21774 29411 21808
rect 29339 21718 29411 21774
rect 29339 21684 29358 21718
rect 29392 21684 29411 21718
rect 29339 21628 29411 21684
rect 29339 21594 29358 21628
rect 29392 21594 29411 21628
rect 29339 21538 29411 21594
rect 29339 21504 29358 21538
rect 29392 21504 29411 21538
rect 29339 21448 29411 21504
rect 29339 21414 29358 21448
rect 29392 21414 29411 21448
rect 29339 21358 29411 21414
rect 28449 21283 28521 21343
rect 29339 21324 29358 21358
rect 29392 21324 29411 21358
rect 29339 21283 29411 21324
rect 28449 21264 29411 21283
rect 28449 21230 28546 21264
rect 28580 21230 28636 21264
rect 28670 21230 28726 21264
rect 28760 21230 28816 21264
rect 28850 21230 28906 21264
rect 28940 21230 28996 21264
rect 29030 21230 29086 21264
rect 29120 21230 29176 21264
rect 29210 21230 29266 21264
rect 29300 21230 29411 21264
rect 28449 21211 29411 21230
rect 29789 22154 30751 22173
rect 29789 22120 29920 22154
rect 29954 22120 30010 22154
rect 30044 22120 30100 22154
rect 30134 22120 30190 22154
rect 30224 22120 30280 22154
rect 30314 22120 30370 22154
rect 30404 22120 30460 22154
rect 30494 22120 30550 22154
rect 30584 22120 30640 22154
rect 30674 22120 30751 22154
rect 29789 22101 30751 22120
rect 29789 22097 29861 22101
rect 29789 22063 29808 22097
rect 29842 22063 29861 22097
rect 29789 22007 29861 22063
rect 30679 22078 30751 22101
rect 30679 22044 30698 22078
rect 30732 22044 30751 22078
rect 29789 21973 29808 22007
rect 29842 21973 29861 22007
rect 29789 21917 29861 21973
rect 29789 21883 29808 21917
rect 29842 21883 29861 21917
rect 29789 21827 29861 21883
rect 29789 21793 29808 21827
rect 29842 21793 29861 21827
rect 29789 21737 29861 21793
rect 29789 21703 29808 21737
rect 29842 21703 29861 21737
rect 29789 21647 29861 21703
rect 29789 21613 29808 21647
rect 29842 21613 29861 21647
rect 29789 21557 29861 21613
rect 29789 21523 29808 21557
rect 29842 21523 29861 21557
rect 29789 21467 29861 21523
rect 29789 21433 29808 21467
rect 29842 21433 29861 21467
rect 29789 21377 29861 21433
rect 29789 21343 29808 21377
rect 29842 21343 29861 21377
rect 30679 21988 30751 22044
rect 30679 21954 30698 21988
rect 30732 21954 30751 21988
rect 30679 21898 30751 21954
rect 30679 21864 30698 21898
rect 30732 21864 30751 21898
rect 30679 21808 30751 21864
rect 30679 21774 30698 21808
rect 30732 21774 30751 21808
rect 30679 21718 30751 21774
rect 30679 21684 30698 21718
rect 30732 21684 30751 21718
rect 30679 21628 30751 21684
rect 30679 21594 30698 21628
rect 30732 21594 30751 21628
rect 30679 21538 30751 21594
rect 30679 21504 30698 21538
rect 30732 21504 30751 21538
rect 30679 21448 30751 21504
rect 30679 21414 30698 21448
rect 30732 21414 30751 21448
rect 30679 21358 30751 21414
rect 29789 21283 29861 21343
rect 30679 21324 30698 21358
rect 30732 21324 30751 21358
rect 30679 21283 30751 21324
rect 29789 21264 30751 21283
rect 29789 21230 29886 21264
rect 29920 21230 29976 21264
rect 30010 21230 30066 21264
rect 30100 21230 30156 21264
rect 30190 21230 30246 21264
rect 30280 21230 30336 21264
rect 30370 21230 30426 21264
rect 30460 21230 30516 21264
rect 30550 21230 30606 21264
rect 30640 21230 30751 21264
rect 29789 21211 30751 21230
rect 31129 22154 32091 22173
rect 31129 22120 31260 22154
rect 31294 22120 31350 22154
rect 31384 22120 31440 22154
rect 31474 22120 31530 22154
rect 31564 22120 31620 22154
rect 31654 22120 31710 22154
rect 31744 22120 31800 22154
rect 31834 22120 31890 22154
rect 31924 22120 31980 22154
rect 32014 22120 32091 22154
rect 31129 22101 32091 22120
rect 31129 22097 31201 22101
rect 31129 22063 31148 22097
rect 31182 22063 31201 22097
rect 31129 22007 31201 22063
rect 32019 22078 32091 22101
rect 32019 22044 32038 22078
rect 32072 22044 32091 22078
rect 31129 21973 31148 22007
rect 31182 21973 31201 22007
rect 31129 21917 31201 21973
rect 31129 21883 31148 21917
rect 31182 21883 31201 21917
rect 31129 21827 31201 21883
rect 31129 21793 31148 21827
rect 31182 21793 31201 21827
rect 31129 21737 31201 21793
rect 31129 21703 31148 21737
rect 31182 21703 31201 21737
rect 31129 21647 31201 21703
rect 31129 21613 31148 21647
rect 31182 21613 31201 21647
rect 31129 21557 31201 21613
rect 31129 21523 31148 21557
rect 31182 21523 31201 21557
rect 31129 21467 31201 21523
rect 31129 21433 31148 21467
rect 31182 21433 31201 21467
rect 31129 21377 31201 21433
rect 31129 21343 31148 21377
rect 31182 21343 31201 21377
rect 32019 21988 32091 22044
rect 32019 21954 32038 21988
rect 32072 21954 32091 21988
rect 32019 21898 32091 21954
rect 32019 21864 32038 21898
rect 32072 21864 32091 21898
rect 32019 21808 32091 21864
rect 32019 21774 32038 21808
rect 32072 21774 32091 21808
rect 32019 21718 32091 21774
rect 32019 21684 32038 21718
rect 32072 21684 32091 21718
rect 32019 21628 32091 21684
rect 32019 21594 32038 21628
rect 32072 21594 32091 21628
rect 32019 21538 32091 21594
rect 32019 21504 32038 21538
rect 32072 21504 32091 21538
rect 32019 21448 32091 21504
rect 32019 21414 32038 21448
rect 32072 21414 32091 21448
rect 32019 21358 32091 21414
rect 31129 21283 31201 21343
rect 32019 21324 32038 21358
rect 32072 21324 32091 21358
rect 32019 21283 32091 21324
rect 31129 21264 32091 21283
rect 31129 21230 31226 21264
rect 31260 21230 31316 21264
rect 31350 21230 31406 21264
rect 31440 21230 31496 21264
rect 31530 21230 31586 21264
rect 31620 21230 31676 21264
rect 31710 21230 31766 21264
rect 31800 21230 31856 21264
rect 31890 21230 31946 21264
rect 31980 21230 32091 21264
rect 31129 21211 32091 21230
rect 32469 22154 33431 22173
rect 32469 22120 32600 22154
rect 32634 22120 32690 22154
rect 32724 22120 32780 22154
rect 32814 22120 32870 22154
rect 32904 22120 32960 22154
rect 32994 22120 33050 22154
rect 33084 22120 33140 22154
rect 33174 22120 33230 22154
rect 33264 22120 33320 22154
rect 33354 22120 33431 22154
rect 32469 22101 33431 22120
rect 32469 22097 32541 22101
rect 32469 22063 32488 22097
rect 32522 22063 32541 22097
rect 32469 22007 32541 22063
rect 33359 22078 33431 22101
rect 33359 22044 33378 22078
rect 33412 22044 33431 22078
rect 32469 21973 32488 22007
rect 32522 21973 32541 22007
rect 32469 21917 32541 21973
rect 32469 21883 32488 21917
rect 32522 21883 32541 21917
rect 32469 21827 32541 21883
rect 32469 21793 32488 21827
rect 32522 21793 32541 21827
rect 32469 21737 32541 21793
rect 32469 21703 32488 21737
rect 32522 21703 32541 21737
rect 32469 21647 32541 21703
rect 32469 21613 32488 21647
rect 32522 21613 32541 21647
rect 32469 21557 32541 21613
rect 32469 21523 32488 21557
rect 32522 21523 32541 21557
rect 32469 21467 32541 21523
rect 32469 21433 32488 21467
rect 32522 21433 32541 21467
rect 32469 21377 32541 21433
rect 32469 21343 32488 21377
rect 32522 21343 32541 21377
rect 33359 21988 33431 22044
rect 33359 21954 33378 21988
rect 33412 21954 33431 21988
rect 33359 21898 33431 21954
rect 33359 21864 33378 21898
rect 33412 21864 33431 21898
rect 33359 21808 33431 21864
rect 33359 21774 33378 21808
rect 33412 21774 33431 21808
rect 33359 21718 33431 21774
rect 33359 21684 33378 21718
rect 33412 21684 33431 21718
rect 33359 21628 33431 21684
rect 33359 21594 33378 21628
rect 33412 21594 33431 21628
rect 33359 21538 33431 21594
rect 33359 21504 33378 21538
rect 33412 21504 33431 21538
rect 33359 21448 33431 21504
rect 33359 21414 33378 21448
rect 33412 21414 33431 21448
rect 33359 21358 33431 21414
rect 32469 21283 32541 21343
rect 33359 21324 33378 21358
rect 33412 21324 33431 21358
rect 33359 21283 33431 21324
rect 32469 21264 33431 21283
rect 32469 21230 32566 21264
rect 32600 21230 32656 21264
rect 32690 21230 32746 21264
rect 32780 21230 32836 21264
rect 32870 21230 32926 21264
rect 32960 21230 33016 21264
rect 33050 21230 33106 21264
rect 33140 21230 33196 21264
rect 33230 21230 33286 21264
rect 33320 21230 33431 21264
rect 32469 21211 33431 21230
rect 33809 22154 34771 22173
rect 33809 22120 33940 22154
rect 33974 22120 34030 22154
rect 34064 22120 34120 22154
rect 34154 22120 34210 22154
rect 34244 22120 34300 22154
rect 34334 22120 34390 22154
rect 34424 22120 34480 22154
rect 34514 22120 34570 22154
rect 34604 22120 34660 22154
rect 34694 22120 34771 22154
rect 33809 22101 34771 22120
rect 33809 22097 33881 22101
rect 33809 22063 33828 22097
rect 33862 22063 33881 22097
rect 33809 22007 33881 22063
rect 34699 22078 34771 22101
rect 34699 22044 34718 22078
rect 34752 22044 34771 22078
rect 33809 21973 33828 22007
rect 33862 21973 33881 22007
rect 33809 21917 33881 21973
rect 33809 21883 33828 21917
rect 33862 21883 33881 21917
rect 33809 21827 33881 21883
rect 33809 21793 33828 21827
rect 33862 21793 33881 21827
rect 33809 21737 33881 21793
rect 33809 21703 33828 21737
rect 33862 21703 33881 21737
rect 33809 21647 33881 21703
rect 33809 21613 33828 21647
rect 33862 21613 33881 21647
rect 33809 21557 33881 21613
rect 33809 21523 33828 21557
rect 33862 21523 33881 21557
rect 33809 21467 33881 21523
rect 33809 21433 33828 21467
rect 33862 21433 33881 21467
rect 33809 21377 33881 21433
rect 33809 21343 33828 21377
rect 33862 21343 33881 21377
rect 34699 21988 34771 22044
rect 34699 21954 34718 21988
rect 34752 21954 34771 21988
rect 34699 21898 34771 21954
rect 34699 21864 34718 21898
rect 34752 21864 34771 21898
rect 34699 21808 34771 21864
rect 34699 21774 34718 21808
rect 34752 21774 34771 21808
rect 34699 21718 34771 21774
rect 34699 21684 34718 21718
rect 34752 21684 34771 21718
rect 34699 21628 34771 21684
rect 34699 21594 34718 21628
rect 34752 21594 34771 21628
rect 34699 21538 34771 21594
rect 34699 21504 34718 21538
rect 34752 21504 34771 21538
rect 34699 21448 34771 21504
rect 34699 21414 34718 21448
rect 34752 21414 34771 21448
rect 34699 21358 34771 21414
rect 33809 21283 33881 21343
rect 34699 21324 34718 21358
rect 34752 21324 34771 21358
rect 34699 21283 34771 21324
rect 33809 21264 34771 21283
rect 33809 21230 33906 21264
rect 33940 21230 33996 21264
rect 34030 21230 34086 21264
rect 34120 21230 34176 21264
rect 34210 21230 34266 21264
rect 34300 21230 34356 21264
rect 34390 21230 34446 21264
rect 34480 21230 34536 21264
rect 34570 21230 34626 21264
rect 34660 21230 34771 21264
rect 33809 21211 34771 21230
rect 35149 22154 36111 22173
rect 35149 22120 35280 22154
rect 35314 22120 35370 22154
rect 35404 22120 35460 22154
rect 35494 22120 35550 22154
rect 35584 22120 35640 22154
rect 35674 22120 35730 22154
rect 35764 22120 35820 22154
rect 35854 22120 35910 22154
rect 35944 22120 36000 22154
rect 36034 22120 36111 22154
rect 35149 22101 36111 22120
rect 35149 22097 35221 22101
rect 35149 22063 35168 22097
rect 35202 22063 35221 22097
rect 35149 22007 35221 22063
rect 36039 22078 36111 22101
rect 36039 22044 36058 22078
rect 36092 22044 36111 22078
rect 35149 21973 35168 22007
rect 35202 21973 35221 22007
rect 35149 21917 35221 21973
rect 35149 21883 35168 21917
rect 35202 21883 35221 21917
rect 35149 21827 35221 21883
rect 35149 21793 35168 21827
rect 35202 21793 35221 21827
rect 35149 21737 35221 21793
rect 35149 21703 35168 21737
rect 35202 21703 35221 21737
rect 35149 21647 35221 21703
rect 35149 21613 35168 21647
rect 35202 21613 35221 21647
rect 35149 21557 35221 21613
rect 35149 21523 35168 21557
rect 35202 21523 35221 21557
rect 35149 21467 35221 21523
rect 35149 21433 35168 21467
rect 35202 21433 35221 21467
rect 35149 21377 35221 21433
rect 35149 21343 35168 21377
rect 35202 21343 35221 21377
rect 36039 21988 36111 22044
rect 36039 21954 36058 21988
rect 36092 21954 36111 21988
rect 36039 21898 36111 21954
rect 36039 21864 36058 21898
rect 36092 21864 36111 21898
rect 36039 21808 36111 21864
rect 36039 21774 36058 21808
rect 36092 21774 36111 21808
rect 36039 21718 36111 21774
rect 36039 21684 36058 21718
rect 36092 21684 36111 21718
rect 36039 21628 36111 21684
rect 36039 21594 36058 21628
rect 36092 21594 36111 21628
rect 36039 21538 36111 21594
rect 36039 21504 36058 21538
rect 36092 21504 36111 21538
rect 36039 21448 36111 21504
rect 36039 21414 36058 21448
rect 36092 21414 36111 21448
rect 36039 21358 36111 21414
rect 35149 21283 35221 21343
rect 36039 21324 36058 21358
rect 36092 21324 36111 21358
rect 36039 21283 36111 21324
rect 35149 21264 36111 21283
rect 35149 21230 35246 21264
rect 35280 21230 35336 21264
rect 35370 21230 35426 21264
rect 35460 21230 35516 21264
rect 35550 21230 35606 21264
rect 35640 21230 35696 21264
rect 35730 21230 35786 21264
rect 35820 21230 35876 21264
rect 35910 21230 35966 21264
rect 36000 21230 36111 21264
rect 35149 21211 36111 21230
rect 36489 22154 37451 22173
rect 36489 22120 36620 22154
rect 36654 22120 36710 22154
rect 36744 22120 36800 22154
rect 36834 22120 36890 22154
rect 36924 22120 36980 22154
rect 37014 22120 37070 22154
rect 37104 22120 37160 22154
rect 37194 22120 37250 22154
rect 37284 22120 37340 22154
rect 37374 22120 37451 22154
rect 36489 22101 37451 22120
rect 36489 22097 36561 22101
rect 36489 22063 36508 22097
rect 36542 22063 36561 22097
rect 36489 22007 36561 22063
rect 37379 22078 37451 22101
rect 37379 22044 37398 22078
rect 37432 22044 37451 22078
rect 36489 21973 36508 22007
rect 36542 21973 36561 22007
rect 36489 21917 36561 21973
rect 36489 21883 36508 21917
rect 36542 21883 36561 21917
rect 36489 21827 36561 21883
rect 36489 21793 36508 21827
rect 36542 21793 36561 21827
rect 36489 21737 36561 21793
rect 36489 21703 36508 21737
rect 36542 21703 36561 21737
rect 36489 21647 36561 21703
rect 36489 21613 36508 21647
rect 36542 21613 36561 21647
rect 36489 21557 36561 21613
rect 36489 21523 36508 21557
rect 36542 21523 36561 21557
rect 36489 21467 36561 21523
rect 36489 21433 36508 21467
rect 36542 21433 36561 21467
rect 36489 21377 36561 21433
rect 36489 21343 36508 21377
rect 36542 21343 36561 21377
rect 37379 21988 37451 22044
rect 37379 21954 37398 21988
rect 37432 21954 37451 21988
rect 37379 21898 37451 21954
rect 37379 21864 37398 21898
rect 37432 21864 37451 21898
rect 37379 21808 37451 21864
rect 37379 21774 37398 21808
rect 37432 21774 37451 21808
rect 37379 21718 37451 21774
rect 37379 21684 37398 21718
rect 37432 21684 37451 21718
rect 37379 21628 37451 21684
rect 37379 21594 37398 21628
rect 37432 21594 37451 21628
rect 37379 21538 37451 21594
rect 37379 21504 37398 21538
rect 37432 21504 37451 21538
rect 37379 21448 37451 21504
rect 37379 21414 37398 21448
rect 37432 21414 37451 21448
rect 37379 21358 37451 21414
rect 36489 21283 36561 21343
rect 37379 21324 37398 21358
rect 37432 21324 37451 21358
rect 37379 21283 37451 21324
rect 36489 21264 37451 21283
rect 36489 21230 36586 21264
rect 36620 21230 36676 21264
rect 36710 21230 36766 21264
rect 36800 21230 36856 21264
rect 36890 21230 36946 21264
rect 36980 21230 37036 21264
rect 37070 21230 37126 21264
rect 37160 21230 37216 21264
rect 37250 21230 37306 21264
rect 37340 21230 37451 21264
rect 36489 21211 37451 21230
rect 37829 22154 38791 22173
rect 37829 22120 37960 22154
rect 37994 22120 38050 22154
rect 38084 22120 38140 22154
rect 38174 22120 38230 22154
rect 38264 22120 38320 22154
rect 38354 22120 38410 22154
rect 38444 22120 38500 22154
rect 38534 22120 38590 22154
rect 38624 22120 38680 22154
rect 38714 22120 38791 22154
rect 37829 22101 38791 22120
rect 37829 22097 37901 22101
rect 37829 22063 37848 22097
rect 37882 22063 37901 22097
rect 37829 22007 37901 22063
rect 38719 22078 38791 22101
rect 38719 22044 38738 22078
rect 38772 22044 38791 22078
rect 37829 21973 37848 22007
rect 37882 21973 37901 22007
rect 37829 21917 37901 21973
rect 37829 21883 37848 21917
rect 37882 21883 37901 21917
rect 37829 21827 37901 21883
rect 37829 21793 37848 21827
rect 37882 21793 37901 21827
rect 37829 21737 37901 21793
rect 37829 21703 37848 21737
rect 37882 21703 37901 21737
rect 37829 21647 37901 21703
rect 37829 21613 37848 21647
rect 37882 21613 37901 21647
rect 37829 21557 37901 21613
rect 37829 21523 37848 21557
rect 37882 21523 37901 21557
rect 37829 21467 37901 21523
rect 37829 21433 37848 21467
rect 37882 21433 37901 21467
rect 37829 21377 37901 21433
rect 37829 21343 37848 21377
rect 37882 21343 37901 21377
rect 38719 21988 38791 22044
rect 38719 21954 38738 21988
rect 38772 21954 38791 21988
rect 38719 21898 38791 21954
rect 38719 21864 38738 21898
rect 38772 21864 38791 21898
rect 38719 21808 38791 21864
rect 38719 21774 38738 21808
rect 38772 21774 38791 21808
rect 38719 21718 38791 21774
rect 38719 21684 38738 21718
rect 38772 21684 38791 21718
rect 38719 21628 38791 21684
rect 38719 21594 38738 21628
rect 38772 21594 38791 21628
rect 38719 21538 38791 21594
rect 38719 21504 38738 21538
rect 38772 21504 38791 21538
rect 38719 21448 38791 21504
rect 38719 21414 38738 21448
rect 38772 21414 38791 21448
rect 38719 21358 38791 21414
rect 37829 21283 37901 21343
rect 38719 21324 38738 21358
rect 38772 21324 38791 21358
rect 38719 21283 38791 21324
rect 37829 21264 38791 21283
rect 37829 21230 37926 21264
rect 37960 21230 38016 21264
rect 38050 21230 38106 21264
rect 38140 21230 38196 21264
rect 38230 21230 38286 21264
rect 38320 21230 38376 21264
rect 38410 21230 38466 21264
rect 38500 21230 38556 21264
rect 38590 21230 38646 21264
rect 38680 21230 38791 21264
rect 37829 21211 38791 21230
rect 24946 18799 25066 18802
rect 23888 18749 23928 18792
rect 24946 18765 24991 18799
rect 25025 18765 25066 18799
rect 24946 18762 25066 18765
rect 23888 18715 23891 18749
rect 23925 18715 23928 18749
rect 23888 18672 23928 18715
rect 28449 18394 29411 18413
rect 28449 18360 28580 18394
rect 28614 18360 28670 18394
rect 28704 18360 28760 18394
rect 28794 18360 28850 18394
rect 28884 18360 28940 18394
rect 28974 18360 29030 18394
rect 29064 18360 29120 18394
rect 29154 18360 29210 18394
rect 29244 18360 29300 18394
rect 29334 18360 29411 18394
rect 28449 18341 29411 18360
rect 28449 18337 28521 18341
rect 28449 18303 28468 18337
rect 28502 18303 28521 18337
rect 28449 18247 28521 18303
rect 29339 18318 29411 18341
rect 29339 18284 29358 18318
rect 29392 18284 29411 18318
rect 28449 18213 28468 18247
rect 28502 18213 28521 18247
rect 28449 18157 28521 18213
rect 28449 18123 28468 18157
rect 28502 18123 28521 18157
rect 28449 18067 28521 18123
rect 28449 18033 28468 18067
rect 28502 18033 28521 18067
rect 28449 17977 28521 18033
rect 28449 17943 28468 17977
rect 28502 17943 28521 17977
rect 28449 17887 28521 17943
rect 28449 17853 28468 17887
rect 28502 17853 28521 17887
rect 28449 17797 28521 17853
rect 28449 17763 28468 17797
rect 28502 17763 28521 17797
rect 28449 17707 28521 17763
rect 28449 17673 28468 17707
rect 28502 17673 28521 17707
rect 28449 17617 28521 17673
rect 28449 17583 28468 17617
rect 28502 17583 28521 17617
rect 29339 18228 29411 18284
rect 29339 18194 29358 18228
rect 29392 18194 29411 18228
rect 29339 18138 29411 18194
rect 29339 18104 29358 18138
rect 29392 18104 29411 18138
rect 29339 18048 29411 18104
rect 29339 18014 29358 18048
rect 29392 18014 29411 18048
rect 29339 17958 29411 18014
rect 29339 17924 29358 17958
rect 29392 17924 29411 17958
rect 29339 17868 29411 17924
rect 29339 17834 29358 17868
rect 29392 17834 29411 17868
rect 29339 17778 29411 17834
rect 29339 17744 29358 17778
rect 29392 17744 29411 17778
rect 29339 17688 29411 17744
rect 29339 17654 29358 17688
rect 29392 17654 29411 17688
rect 29339 17598 29411 17654
rect 28449 17523 28521 17583
rect 29339 17564 29358 17598
rect 29392 17564 29411 17598
rect 29339 17523 29411 17564
rect 28449 17504 29411 17523
rect 28449 17470 28546 17504
rect 28580 17470 28636 17504
rect 28670 17470 28726 17504
rect 28760 17470 28816 17504
rect 28850 17470 28906 17504
rect 28940 17470 28996 17504
rect 29030 17470 29086 17504
rect 29120 17470 29176 17504
rect 29210 17470 29266 17504
rect 29300 17470 29411 17504
rect 28449 17451 29411 17470
rect 29789 18394 30751 18413
rect 29789 18360 29920 18394
rect 29954 18360 30010 18394
rect 30044 18360 30100 18394
rect 30134 18360 30190 18394
rect 30224 18360 30280 18394
rect 30314 18360 30370 18394
rect 30404 18360 30460 18394
rect 30494 18360 30550 18394
rect 30584 18360 30640 18394
rect 30674 18360 30751 18394
rect 29789 18341 30751 18360
rect 29789 18337 29861 18341
rect 29789 18303 29808 18337
rect 29842 18303 29861 18337
rect 29789 18247 29861 18303
rect 30679 18318 30751 18341
rect 30679 18284 30698 18318
rect 30732 18284 30751 18318
rect 29789 18213 29808 18247
rect 29842 18213 29861 18247
rect 29789 18157 29861 18213
rect 29789 18123 29808 18157
rect 29842 18123 29861 18157
rect 29789 18067 29861 18123
rect 29789 18033 29808 18067
rect 29842 18033 29861 18067
rect 29789 17977 29861 18033
rect 29789 17943 29808 17977
rect 29842 17943 29861 17977
rect 29789 17887 29861 17943
rect 29789 17853 29808 17887
rect 29842 17853 29861 17887
rect 29789 17797 29861 17853
rect 29789 17763 29808 17797
rect 29842 17763 29861 17797
rect 29789 17707 29861 17763
rect 29789 17673 29808 17707
rect 29842 17673 29861 17707
rect 29789 17617 29861 17673
rect 29789 17583 29808 17617
rect 29842 17583 29861 17617
rect 30679 18228 30751 18284
rect 30679 18194 30698 18228
rect 30732 18194 30751 18228
rect 30679 18138 30751 18194
rect 30679 18104 30698 18138
rect 30732 18104 30751 18138
rect 30679 18048 30751 18104
rect 30679 18014 30698 18048
rect 30732 18014 30751 18048
rect 30679 17958 30751 18014
rect 30679 17924 30698 17958
rect 30732 17924 30751 17958
rect 30679 17868 30751 17924
rect 30679 17834 30698 17868
rect 30732 17834 30751 17868
rect 30679 17778 30751 17834
rect 30679 17744 30698 17778
rect 30732 17744 30751 17778
rect 30679 17688 30751 17744
rect 30679 17654 30698 17688
rect 30732 17654 30751 17688
rect 30679 17598 30751 17654
rect 29789 17523 29861 17583
rect 30679 17564 30698 17598
rect 30732 17564 30751 17598
rect 30679 17523 30751 17564
rect 29789 17504 30751 17523
rect 29789 17470 29886 17504
rect 29920 17470 29976 17504
rect 30010 17470 30066 17504
rect 30100 17470 30156 17504
rect 30190 17470 30246 17504
rect 30280 17470 30336 17504
rect 30370 17470 30426 17504
rect 30460 17470 30516 17504
rect 30550 17470 30606 17504
rect 30640 17470 30751 17504
rect 29789 17451 30751 17470
rect 31129 18394 32091 18413
rect 31129 18360 31260 18394
rect 31294 18360 31350 18394
rect 31384 18360 31440 18394
rect 31474 18360 31530 18394
rect 31564 18360 31620 18394
rect 31654 18360 31710 18394
rect 31744 18360 31800 18394
rect 31834 18360 31890 18394
rect 31924 18360 31980 18394
rect 32014 18360 32091 18394
rect 31129 18341 32091 18360
rect 31129 18337 31201 18341
rect 31129 18303 31148 18337
rect 31182 18303 31201 18337
rect 31129 18247 31201 18303
rect 32019 18318 32091 18341
rect 32019 18284 32038 18318
rect 32072 18284 32091 18318
rect 31129 18213 31148 18247
rect 31182 18213 31201 18247
rect 31129 18157 31201 18213
rect 31129 18123 31148 18157
rect 31182 18123 31201 18157
rect 31129 18067 31201 18123
rect 31129 18033 31148 18067
rect 31182 18033 31201 18067
rect 31129 17977 31201 18033
rect 31129 17943 31148 17977
rect 31182 17943 31201 17977
rect 31129 17887 31201 17943
rect 31129 17853 31148 17887
rect 31182 17853 31201 17887
rect 31129 17797 31201 17853
rect 31129 17763 31148 17797
rect 31182 17763 31201 17797
rect 31129 17707 31201 17763
rect 31129 17673 31148 17707
rect 31182 17673 31201 17707
rect 31129 17617 31201 17673
rect 31129 17583 31148 17617
rect 31182 17583 31201 17617
rect 32019 18228 32091 18284
rect 32019 18194 32038 18228
rect 32072 18194 32091 18228
rect 32019 18138 32091 18194
rect 32019 18104 32038 18138
rect 32072 18104 32091 18138
rect 32019 18048 32091 18104
rect 32019 18014 32038 18048
rect 32072 18014 32091 18048
rect 32019 17958 32091 18014
rect 32019 17924 32038 17958
rect 32072 17924 32091 17958
rect 32019 17868 32091 17924
rect 32019 17834 32038 17868
rect 32072 17834 32091 17868
rect 32019 17778 32091 17834
rect 32019 17744 32038 17778
rect 32072 17744 32091 17778
rect 32019 17688 32091 17744
rect 32019 17654 32038 17688
rect 32072 17654 32091 17688
rect 32019 17598 32091 17654
rect 31129 17523 31201 17583
rect 32019 17564 32038 17598
rect 32072 17564 32091 17598
rect 32019 17523 32091 17564
rect 31129 17504 32091 17523
rect 31129 17470 31226 17504
rect 31260 17470 31316 17504
rect 31350 17470 31406 17504
rect 31440 17470 31496 17504
rect 31530 17470 31586 17504
rect 31620 17470 31676 17504
rect 31710 17470 31766 17504
rect 31800 17470 31856 17504
rect 31890 17470 31946 17504
rect 31980 17470 32091 17504
rect 31129 17451 32091 17470
rect 32469 18394 33431 18413
rect 32469 18360 32600 18394
rect 32634 18360 32690 18394
rect 32724 18360 32780 18394
rect 32814 18360 32870 18394
rect 32904 18360 32960 18394
rect 32994 18360 33050 18394
rect 33084 18360 33140 18394
rect 33174 18360 33230 18394
rect 33264 18360 33320 18394
rect 33354 18360 33431 18394
rect 32469 18341 33431 18360
rect 32469 18337 32541 18341
rect 32469 18303 32488 18337
rect 32522 18303 32541 18337
rect 32469 18247 32541 18303
rect 33359 18318 33431 18341
rect 33359 18284 33378 18318
rect 33412 18284 33431 18318
rect 32469 18213 32488 18247
rect 32522 18213 32541 18247
rect 32469 18157 32541 18213
rect 32469 18123 32488 18157
rect 32522 18123 32541 18157
rect 32469 18067 32541 18123
rect 32469 18033 32488 18067
rect 32522 18033 32541 18067
rect 32469 17977 32541 18033
rect 32469 17943 32488 17977
rect 32522 17943 32541 17977
rect 32469 17887 32541 17943
rect 32469 17853 32488 17887
rect 32522 17853 32541 17887
rect 32469 17797 32541 17853
rect 32469 17763 32488 17797
rect 32522 17763 32541 17797
rect 32469 17707 32541 17763
rect 32469 17673 32488 17707
rect 32522 17673 32541 17707
rect 32469 17617 32541 17673
rect 32469 17583 32488 17617
rect 32522 17583 32541 17617
rect 33359 18228 33431 18284
rect 33359 18194 33378 18228
rect 33412 18194 33431 18228
rect 33359 18138 33431 18194
rect 33359 18104 33378 18138
rect 33412 18104 33431 18138
rect 33359 18048 33431 18104
rect 33359 18014 33378 18048
rect 33412 18014 33431 18048
rect 33359 17958 33431 18014
rect 33359 17924 33378 17958
rect 33412 17924 33431 17958
rect 33359 17868 33431 17924
rect 33359 17834 33378 17868
rect 33412 17834 33431 17868
rect 33359 17778 33431 17834
rect 33359 17744 33378 17778
rect 33412 17744 33431 17778
rect 33359 17688 33431 17744
rect 33359 17654 33378 17688
rect 33412 17654 33431 17688
rect 33359 17598 33431 17654
rect 32469 17523 32541 17583
rect 33359 17564 33378 17598
rect 33412 17564 33431 17598
rect 33359 17523 33431 17564
rect 32469 17504 33431 17523
rect 32469 17470 32566 17504
rect 32600 17470 32656 17504
rect 32690 17470 32746 17504
rect 32780 17470 32836 17504
rect 32870 17470 32926 17504
rect 32960 17470 33016 17504
rect 33050 17470 33106 17504
rect 33140 17470 33196 17504
rect 33230 17470 33286 17504
rect 33320 17470 33431 17504
rect 32469 17451 33431 17470
rect 33809 18394 34771 18413
rect 33809 18360 33940 18394
rect 33974 18360 34030 18394
rect 34064 18360 34120 18394
rect 34154 18360 34210 18394
rect 34244 18360 34300 18394
rect 34334 18360 34390 18394
rect 34424 18360 34480 18394
rect 34514 18360 34570 18394
rect 34604 18360 34660 18394
rect 34694 18360 34771 18394
rect 33809 18341 34771 18360
rect 33809 18337 33881 18341
rect 33809 18303 33828 18337
rect 33862 18303 33881 18337
rect 33809 18247 33881 18303
rect 34699 18318 34771 18341
rect 34699 18284 34718 18318
rect 34752 18284 34771 18318
rect 33809 18213 33828 18247
rect 33862 18213 33881 18247
rect 33809 18157 33881 18213
rect 33809 18123 33828 18157
rect 33862 18123 33881 18157
rect 33809 18067 33881 18123
rect 33809 18033 33828 18067
rect 33862 18033 33881 18067
rect 33809 17977 33881 18033
rect 33809 17943 33828 17977
rect 33862 17943 33881 17977
rect 33809 17887 33881 17943
rect 33809 17853 33828 17887
rect 33862 17853 33881 17887
rect 33809 17797 33881 17853
rect 33809 17763 33828 17797
rect 33862 17763 33881 17797
rect 33809 17707 33881 17763
rect 33809 17673 33828 17707
rect 33862 17673 33881 17707
rect 33809 17617 33881 17673
rect 33809 17583 33828 17617
rect 33862 17583 33881 17617
rect 34699 18228 34771 18284
rect 34699 18194 34718 18228
rect 34752 18194 34771 18228
rect 34699 18138 34771 18194
rect 34699 18104 34718 18138
rect 34752 18104 34771 18138
rect 34699 18048 34771 18104
rect 34699 18014 34718 18048
rect 34752 18014 34771 18048
rect 34699 17958 34771 18014
rect 34699 17924 34718 17958
rect 34752 17924 34771 17958
rect 34699 17868 34771 17924
rect 34699 17834 34718 17868
rect 34752 17834 34771 17868
rect 34699 17778 34771 17834
rect 34699 17744 34718 17778
rect 34752 17744 34771 17778
rect 34699 17688 34771 17744
rect 34699 17654 34718 17688
rect 34752 17654 34771 17688
rect 34699 17598 34771 17654
rect 33809 17523 33881 17583
rect 34699 17564 34718 17598
rect 34752 17564 34771 17598
rect 34699 17523 34771 17564
rect 33809 17504 34771 17523
rect 33809 17470 33906 17504
rect 33940 17470 33996 17504
rect 34030 17470 34086 17504
rect 34120 17470 34176 17504
rect 34210 17470 34266 17504
rect 34300 17470 34356 17504
rect 34390 17470 34446 17504
rect 34480 17470 34536 17504
rect 34570 17470 34626 17504
rect 34660 17470 34771 17504
rect 33809 17451 34771 17470
rect 35149 18394 36111 18413
rect 35149 18360 35280 18394
rect 35314 18360 35370 18394
rect 35404 18360 35460 18394
rect 35494 18360 35550 18394
rect 35584 18360 35640 18394
rect 35674 18360 35730 18394
rect 35764 18360 35820 18394
rect 35854 18360 35910 18394
rect 35944 18360 36000 18394
rect 36034 18360 36111 18394
rect 35149 18341 36111 18360
rect 35149 18337 35221 18341
rect 35149 18303 35168 18337
rect 35202 18303 35221 18337
rect 35149 18247 35221 18303
rect 36039 18318 36111 18341
rect 36039 18284 36058 18318
rect 36092 18284 36111 18318
rect 35149 18213 35168 18247
rect 35202 18213 35221 18247
rect 35149 18157 35221 18213
rect 35149 18123 35168 18157
rect 35202 18123 35221 18157
rect 35149 18067 35221 18123
rect 35149 18033 35168 18067
rect 35202 18033 35221 18067
rect 35149 17977 35221 18033
rect 35149 17943 35168 17977
rect 35202 17943 35221 17977
rect 35149 17887 35221 17943
rect 35149 17853 35168 17887
rect 35202 17853 35221 17887
rect 35149 17797 35221 17853
rect 35149 17763 35168 17797
rect 35202 17763 35221 17797
rect 35149 17707 35221 17763
rect 35149 17673 35168 17707
rect 35202 17673 35221 17707
rect 35149 17617 35221 17673
rect 35149 17583 35168 17617
rect 35202 17583 35221 17617
rect 36039 18228 36111 18284
rect 36039 18194 36058 18228
rect 36092 18194 36111 18228
rect 36039 18138 36111 18194
rect 36039 18104 36058 18138
rect 36092 18104 36111 18138
rect 36039 18048 36111 18104
rect 36039 18014 36058 18048
rect 36092 18014 36111 18048
rect 36039 17958 36111 18014
rect 36039 17924 36058 17958
rect 36092 17924 36111 17958
rect 36039 17868 36111 17924
rect 36039 17834 36058 17868
rect 36092 17834 36111 17868
rect 36039 17778 36111 17834
rect 36039 17744 36058 17778
rect 36092 17744 36111 17778
rect 36039 17688 36111 17744
rect 36039 17654 36058 17688
rect 36092 17654 36111 17688
rect 36039 17598 36111 17654
rect 35149 17523 35221 17583
rect 36039 17564 36058 17598
rect 36092 17564 36111 17598
rect 36039 17523 36111 17564
rect 35149 17504 36111 17523
rect 35149 17470 35246 17504
rect 35280 17470 35336 17504
rect 35370 17470 35426 17504
rect 35460 17470 35516 17504
rect 35550 17470 35606 17504
rect 35640 17470 35696 17504
rect 35730 17470 35786 17504
rect 35820 17470 35876 17504
rect 35910 17470 35966 17504
rect 36000 17470 36111 17504
rect 35149 17451 36111 17470
rect 36489 18394 37451 18413
rect 36489 18360 36620 18394
rect 36654 18360 36710 18394
rect 36744 18360 36800 18394
rect 36834 18360 36890 18394
rect 36924 18360 36980 18394
rect 37014 18360 37070 18394
rect 37104 18360 37160 18394
rect 37194 18360 37250 18394
rect 37284 18360 37340 18394
rect 37374 18360 37451 18394
rect 36489 18341 37451 18360
rect 36489 18337 36561 18341
rect 36489 18303 36508 18337
rect 36542 18303 36561 18337
rect 36489 18247 36561 18303
rect 37379 18318 37451 18341
rect 37379 18284 37398 18318
rect 37432 18284 37451 18318
rect 36489 18213 36508 18247
rect 36542 18213 36561 18247
rect 36489 18157 36561 18213
rect 36489 18123 36508 18157
rect 36542 18123 36561 18157
rect 36489 18067 36561 18123
rect 36489 18033 36508 18067
rect 36542 18033 36561 18067
rect 36489 17977 36561 18033
rect 36489 17943 36508 17977
rect 36542 17943 36561 17977
rect 36489 17887 36561 17943
rect 36489 17853 36508 17887
rect 36542 17853 36561 17887
rect 36489 17797 36561 17853
rect 36489 17763 36508 17797
rect 36542 17763 36561 17797
rect 36489 17707 36561 17763
rect 36489 17673 36508 17707
rect 36542 17673 36561 17707
rect 36489 17617 36561 17673
rect 36489 17583 36508 17617
rect 36542 17583 36561 17617
rect 37379 18228 37451 18284
rect 37379 18194 37398 18228
rect 37432 18194 37451 18228
rect 37379 18138 37451 18194
rect 37379 18104 37398 18138
rect 37432 18104 37451 18138
rect 37379 18048 37451 18104
rect 37379 18014 37398 18048
rect 37432 18014 37451 18048
rect 37379 17958 37451 18014
rect 37379 17924 37398 17958
rect 37432 17924 37451 17958
rect 37379 17868 37451 17924
rect 37379 17834 37398 17868
rect 37432 17834 37451 17868
rect 37379 17778 37451 17834
rect 37379 17744 37398 17778
rect 37432 17744 37451 17778
rect 37379 17688 37451 17744
rect 37379 17654 37398 17688
rect 37432 17654 37451 17688
rect 37379 17598 37451 17654
rect 36489 17523 36561 17583
rect 37379 17564 37398 17598
rect 37432 17564 37451 17598
rect 37379 17523 37451 17564
rect 36489 17504 37451 17523
rect 36489 17470 36586 17504
rect 36620 17470 36676 17504
rect 36710 17470 36766 17504
rect 36800 17470 36856 17504
rect 36890 17470 36946 17504
rect 36980 17470 37036 17504
rect 37070 17470 37126 17504
rect 37160 17470 37216 17504
rect 37250 17470 37306 17504
rect 37340 17470 37451 17504
rect 36489 17451 37451 17470
rect 37829 18394 38791 18413
rect 37829 18360 37960 18394
rect 37994 18360 38050 18394
rect 38084 18360 38140 18394
rect 38174 18360 38230 18394
rect 38264 18360 38320 18394
rect 38354 18360 38410 18394
rect 38444 18360 38500 18394
rect 38534 18360 38590 18394
rect 38624 18360 38680 18394
rect 38714 18360 38791 18394
rect 37829 18341 38791 18360
rect 37829 18337 37901 18341
rect 37829 18303 37848 18337
rect 37882 18303 37901 18337
rect 37829 18247 37901 18303
rect 38719 18318 38791 18341
rect 38719 18284 38738 18318
rect 38772 18284 38791 18318
rect 37829 18213 37848 18247
rect 37882 18213 37901 18247
rect 37829 18157 37901 18213
rect 37829 18123 37848 18157
rect 37882 18123 37901 18157
rect 37829 18067 37901 18123
rect 37829 18033 37848 18067
rect 37882 18033 37901 18067
rect 37829 17977 37901 18033
rect 37829 17943 37848 17977
rect 37882 17943 37901 17977
rect 37829 17887 37901 17943
rect 37829 17853 37848 17887
rect 37882 17853 37901 17887
rect 37829 17797 37901 17853
rect 37829 17763 37848 17797
rect 37882 17763 37901 17797
rect 37829 17707 37901 17763
rect 37829 17673 37848 17707
rect 37882 17673 37901 17707
rect 37829 17617 37901 17673
rect 37829 17583 37848 17617
rect 37882 17583 37901 17617
rect 38719 18228 38791 18284
rect 38719 18194 38738 18228
rect 38772 18194 38791 18228
rect 38719 18138 38791 18194
rect 38719 18104 38738 18138
rect 38772 18104 38791 18138
rect 38719 18048 38791 18104
rect 38719 18014 38738 18048
rect 38772 18014 38791 18048
rect 38719 17958 38791 18014
rect 38719 17924 38738 17958
rect 38772 17924 38791 17958
rect 38719 17868 38791 17924
rect 38719 17834 38738 17868
rect 38772 17834 38791 17868
rect 38719 17778 38791 17834
rect 38719 17744 38738 17778
rect 38772 17744 38791 17778
rect 38719 17688 38791 17744
rect 38719 17654 38738 17688
rect 38772 17654 38791 17688
rect 38719 17598 38791 17654
rect 37829 17523 37901 17583
rect 38719 17564 38738 17598
rect 38772 17564 38791 17598
rect 38719 17523 38791 17564
rect 37829 17504 38791 17523
rect 37829 17470 37926 17504
rect 37960 17470 38016 17504
rect 38050 17470 38106 17504
rect 38140 17470 38196 17504
rect 38230 17470 38286 17504
rect 38320 17470 38376 17504
rect 38410 17470 38466 17504
rect 38500 17470 38556 17504
rect 38590 17470 38646 17504
rect 38680 17470 38791 17504
rect 37829 17451 38791 17470
rect 28449 14634 29411 14653
rect 28449 14600 28580 14634
rect 28614 14600 28670 14634
rect 28704 14600 28760 14634
rect 28794 14600 28850 14634
rect 28884 14600 28940 14634
rect 28974 14600 29030 14634
rect 29064 14600 29120 14634
rect 29154 14600 29210 14634
rect 29244 14600 29300 14634
rect 29334 14600 29411 14634
rect 28449 14581 29411 14600
rect 28449 14577 28521 14581
rect 28449 14543 28468 14577
rect 28502 14543 28521 14577
rect 28449 14487 28521 14543
rect 29339 14558 29411 14581
rect 29339 14524 29358 14558
rect 29392 14524 29411 14558
rect 28449 14453 28468 14487
rect 28502 14453 28521 14487
rect 28449 14397 28521 14453
rect 28449 14363 28468 14397
rect 28502 14363 28521 14397
rect 28449 14307 28521 14363
rect 28449 14273 28468 14307
rect 28502 14273 28521 14307
rect 28449 14217 28521 14273
rect 28449 14183 28468 14217
rect 28502 14183 28521 14217
rect 28449 14127 28521 14183
rect 28449 14093 28468 14127
rect 28502 14093 28521 14127
rect 28449 14037 28521 14093
rect 28449 14003 28468 14037
rect 28502 14003 28521 14037
rect 28449 13947 28521 14003
rect 28449 13913 28468 13947
rect 28502 13913 28521 13947
rect 28449 13857 28521 13913
rect 28449 13823 28468 13857
rect 28502 13823 28521 13857
rect 29339 14468 29411 14524
rect 29339 14434 29358 14468
rect 29392 14434 29411 14468
rect 29339 14378 29411 14434
rect 29339 14344 29358 14378
rect 29392 14344 29411 14378
rect 29339 14288 29411 14344
rect 29339 14254 29358 14288
rect 29392 14254 29411 14288
rect 29339 14198 29411 14254
rect 29339 14164 29358 14198
rect 29392 14164 29411 14198
rect 29339 14108 29411 14164
rect 29339 14074 29358 14108
rect 29392 14074 29411 14108
rect 29339 14018 29411 14074
rect 29339 13984 29358 14018
rect 29392 13984 29411 14018
rect 29339 13928 29411 13984
rect 29339 13894 29358 13928
rect 29392 13894 29411 13928
rect 29339 13838 29411 13894
rect 28449 13763 28521 13823
rect 29339 13804 29358 13838
rect 29392 13804 29411 13838
rect 29339 13763 29411 13804
rect 28449 13744 29411 13763
rect 28449 13710 28546 13744
rect 28580 13710 28636 13744
rect 28670 13710 28726 13744
rect 28760 13710 28816 13744
rect 28850 13710 28906 13744
rect 28940 13710 28996 13744
rect 29030 13710 29086 13744
rect 29120 13710 29176 13744
rect 29210 13710 29266 13744
rect 29300 13710 29411 13744
rect 28449 13691 29411 13710
rect 29789 14634 30751 14653
rect 29789 14600 29920 14634
rect 29954 14600 30010 14634
rect 30044 14600 30100 14634
rect 30134 14600 30190 14634
rect 30224 14600 30280 14634
rect 30314 14600 30370 14634
rect 30404 14600 30460 14634
rect 30494 14600 30550 14634
rect 30584 14600 30640 14634
rect 30674 14600 30751 14634
rect 29789 14581 30751 14600
rect 29789 14577 29861 14581
rect 29789 14543 29808 14577
rect 29842 14543 29861 14577
rect 29789 14487 29861 14543
rect 30679 14558 30751 14581
rect 30679 14524 30698 14558
rect 30732 14524 30751 14558
rect 29789 14453 29808 14487
rect 29842 14453 29861 14487
rect 29789 14397 29861 14453
rect 29789 14363 29808 14397
rect 29842 14363 29861 14397
rect 29789 14307 29861 14363
rect 29789 14273 29808 14307
rect 29842 14273 29861 14307
rect 29789 14217 29861 14273
rect 29789 14183 29808 14217
rect 29842 14183 29861 14217
rect 29789 14127 29861 14183
rect 29789 14093 29808 14127
rect 29842 14093 29861 14127
rect 29789 14037 29861 14093
rect 29789 14003 29808 14037
rect 29842 14003 29861 14037
rect 29789 13947 29861 14003
rect 29789 13913 29808 13947
rect 29842 13913 29861 13947
rect 29789 13857 29861 13913
rect 29789 13823 29808 13857
rect 29842 13823 29861 13857
rect 30679 14468 30751 14524
rect 30679 14434 30698 14468
rect 30732 14434 30751 14468
rect 30679 14378 30751 14434
rect 30679 14344 30698 14378
rect 30732 14344 30751 14378
rect 30679 14288 30751 14344
rect 30679 14254 30698 14288
rect 30732 14254 30751 14288
rect 30679 14198 30751 14254
rect 30679 14164 30698 14198
rect 30732 14164 30751 14198
rect 30679 14108 30751 14164
rect 30679 14074 30698 14108
rect 30732 14074 30751 14108
rect 30679 14018 30751 14074
rect 30679 13984 30698 14018
rect 30732 13984 30751 14018
rect 30679 13928 30751 13984
rect 30679 13894 30698 13928
rect 30732 13894 30751 13928
rect 30679 13838 30751 13894
rect 29789 13763 29861 13823
rect 30679 13804 30698 13838
rect 30732 13804 30751 13838
rect 30679 13763 30751 13804
rect 29789 13744 30751 13763
rect 29789 13710 29886 13744
rect 29920 13710 29976 13744
rect 30010 13710 30066 13744
rect 30100 13710 30156 13744
rect 30190 13710 30246 13744
rect 30280 13710 30336 13744
rect 30370 13710 30426 13744
rect 30460 13710 30516 13744
rect 30550 13710 30606 13744
rect 30640 13710 30751 13744
rect 29789 13691 30751 13710
rect 31129 14634 32091 14653
rect 31129 14600 31260 14634
rect 31294 14600 31350 14634
rect 31384 14600 31440 14634
rect 31474 14600 31530 14634
rect 31564 14600 31620 14634
rect 31654 14600 31710 14634
rect 31744 14600 31800 14634
rect 31834 14600 31890 14634
rect 31924 14600 31980 14634
rect 32014 14600 32091 14634
rect 31129 14581 32091 14600
rect 31129 14577 31201 14581
rect 31129 14543 31148 14577
rect 31182 14543 31201 14577
rect 31129 14487 31201 14543
rect 32019 14558 32091 14581
rect 32019 14524 32038 14558
rect 32072 14524 32091 14558
rect 31129 14453 31148 14487
rect 31182 14453 31201 14487
rect 31129 14397 31201 14453
rect 31129 14363 31148 14397
rect 31182 14363 31201 14397
rect 31129 14307 31201 14363
rect 31129 14273 31148 14307
rect 31182 14273 31201 14307
rect 31129 14217 31201 14273
rect 31129 14183 31148 14217
rect 31182 14183 31201 14217
rect 31129 14127 31201 14183
rect 31129 14093 31148 14127
rect 31182 14093 31201 14127
rect 31129 14037 31201 14093
rect 31129 14003 31148 14037
rect 31182 14003 31201 14037
rect 31129 13947 31201 14003
rect 31129 13913 31148 13947
rect 31182 13913 31201 13947
rect 31129 13857 31201 13913
rect 31129 13823 31148 13857
rect 31182 13823 31201 13857
rect 32019 14468 32091 14524
rect 32019 14434 32038 14468
rect 32072 14434 32091 14468
rect 32019 14378 32091 14434
rect 32019 14344 32038 14378
rect 32072 14344 32091 14378
rect 32019 14288 32091 14344
rect 32019 14254 32038 14288
rect 32072 14254 32091 14288
rect 32019 14198 32091 14254
rect 32019 14164 32038 14198
rect 32072 14164 32091 14198
rect 32019 14108 32091 14164
rect 32019 14074 32038 14108
rect 32072 14074 32091 14108
rect 32019 14018 32091 14074
rect 32019 13984 32038 14018
rect 32072 13984 32091 14018
rect 32019 13928 32091 13984
rect 32019 13894 32038 13928
rect 32072 13894 32091 13928
rect 32019 13838 32091 13894
rect 31129 13763 31201 13823
rect 32019 13804 32038 13838
rect 32072 13804 32091 13838
rect 32019 13763 32091 13804
rect 31129 13744 32091 13763
rect 31129 13710 31226 13744
rect 31260 13710 31316 13744
rect 31350 13710 31406 13744
rect 31440 13710 31496 13744
rect 31530 13710 31586 13744
rect 31620 13710 31676 13744
rect 31710 13710 31766 13744
rect 31800 13710 31856 13744
rect 31890 13710 31946 13744
rect 31980 13710 32091 13744
rect 31129 13691 32091 13710
rect 32469 14634 33431 14653
rect 32469 14600 32600 14634
rect 32634 14600 32690 14634
rect 32724 14600 32780 14634
rect 32814 14600 32870 14634
rect 32904 14600 32960 14634
rect 32994 14600 33050 14634
rect 33084 14600 33140 14634
rect 33174 14600 33230 14634
rect 33264 14600 33320 14634
rect 33354 14600 33431 14634
rect 32469 14581 33431 14600
rect 32469 14577 32541 14581
rect 32469 14543 32488 14577
rect 32522 14543 32541 14577
rect 32469 14487 32541 14543
rect 33359 14558 33431 14581
rect 33359 14524 33378 14558
rect 33412 14524 33431 14558
rect 32469 14453 32488 14487
rect 32522 14453 32541 14487
rect 32469 14397 32541 14453
rect 32469 14363 32488 14397
rect 32522 14363 32541 14397
rect 32469 14307 32541 14363
rect 32469 14273 32488 14307
rect 32522 14273 32541 14307
rect 32469 14217 32541 14273
rect 32469 14183 32488 14217
rect 32522 14183 32541 14217
rect 32469 14127 32541 14183
rect 32469 14093 32488 14127
rect 32522 14093 32541 14127
rect 32469 14037 32541 14093
rect 32469 14003 32488 14037
rect 32522 14003 32541 14037
rect 32469 13947 32541 14003
rect 32469 13913 32488 13947
rect 32522 13913 32541 13947
rect 32469 13857 32541 13913
rect 32469 13823 32488 13857
rect 32522 13823 32541 13857
rect 33359 14468 33431 14524
rect 33359 14434 33378 14468
rect 33412 14434 33431 14468
rect 33359 14378 33431 14434
rect 33359 14344 33378 14378
rect 33412 14344 33431 14378
rect 33359 14288 33431 14344
rect 33359 14254 33378 14288
rect 33412 14254 33431 14288
rect 33359 14198 33431 14254
rect 33359 14164 33378 14198
rect 33412 14164 33431 14198
rect 33359 14108 33431 14164
rect 33359 14074 33378 14108
rect 33412 14074 33431 14108
rect 33359 14018 33431 14074
rect 33359 13984 33378 14018
rect 33412 13984 33431 14018
rect 33359 13928 33431 13984
rect 33359 13894 33378 13928
rect 33412 13894 33431 13928
rect 33359 13838 33431 13894
rect 32469 13763 32541 13823
rect 33359 13804 33378 13838
rect 33412 13804 33431 13838
rect 33359 13763 33431 13804
rect 32469 13744 33431 13763
rect 32469 13710 32566 13744
rect 32600 13710 32656 13744
rect 32690 13710 32746 13744
rect 32780 13710 32836 13744
rect 32870 13710 32926 13744
rect 32960 13710 33016 13744
rect 33050 13710 33106 13744
rect 33140 13710 33196 13744
rect 33230 13710 33286 13744
rect 33320 13710 33431 13744
rect 32469 13691 33431 13710
rect 33809 14634 34771 14653
rect 33809 14600 33940 14634
rect 33974 14600 34030 14634
rect 34064 14600 34120 14634
rect 34154 14600 34210 14634
rect 34244 14600 34300 14634
rect 34334 14600 34390 14634
rect 34424 14600 34480 14634
rect 34514 14600 34570 14634
rect 34604 14600 34660 14634
rect 34694 14600 34771 14634
rect 33809 14581 34771 14600
rect 33809 14577 33881 14581
rect 33809 14543 33828 14577
rect 33862 14543 33881 14577
rect 33809 14487 33881 14543
rect 34699 14558 34771 14581
rect 34699 14524 34718 14558
rect 34752 14524 34771 14558
rect 33809 14453 33828 14487
rect 33862 14453 33881 14487
rect 33809 14397 33881 14453
rect 33809 14363 33828 14397
rect 33862 14363 33881 14397
rect 33809 14307 33881 14363
rect 33809 14273 33828 14307
rect 33862 14273 33881 14307
rect 33809 14217 33881 14273
rect 33809 14183 33828 14217
rect 33862 14183 33881 14217
rect 33809 14127 33881 14183
rect 33809 14093 33828 14127
rect 33862 14093 33881 14127
rect 33809 14037 33881 14093
rect 33809 14003 33828 14037
rect 33862 14003 33881 14037
rect 33809 13947 33881 14003
rect 33809 13913 33828 13947
rect 33862 13913 33881 13947
rect 33809 13857 33881 13913
rect 33809 13823 33828 13857
rect 33862 13823 33881 13857
rect 34699 14468 34771 14524
rect 34699 14434 34718 14468
rect 34752 14434 34771 14468
rect 34699 14378 34771 14434
rect 34699 14344 34718 14378
rect 34752 14344 34771 14378
rect 34699 14288 34771 14344
rect 34699 14254 34718 14288
rect 34752 14254 34771 14288
rect 34699 14198 34771 14254
rect 34699 14164 34718 14198
rect 34752 14164 34771 14198
rect 34699 14108 34771 14164
rect 34699 14074 34718 14108
rect 34752 14074 34771 14108
rect 34699 14018 34771 14074
rect 34699 13984 34718 14018
rect 34752 13984 34771 14018
rect 34699 13928 34771 13984
rect 34699 13894 34718 13928
rect 34752 13894 34771 13928
rect 34699 13838 34771 13894
rect 33809 13763 33881 13823
rect 34699 13804 34718 13838
rect 34752 13804 34771 13838
rect 34699 13763 34771 13804
rect 33809 13744 34771 13763
rect 33809 13710 33906 13744
rect 33940 13710 33996 13744
rect 34030 13710 34086 13744
rect 34120 13710 34176 13744
rect 34210 13710 34266 13744
rect 34300 13710 34356 13744
rect 34390 13710 34446 13744
rect 34480 13710 34536 13744
rect 34570 13710 34626 13744
rect 34660 13710 34771 13744
rect 33809 13691 34771 13710
rect 35149 14634 36111 14653
rect 35149 14600 35280 14634
rect 35314 14600 35370 14634
rect 35404 14600 35460 14634
rect 35494 14600 35550 14634
rect 35584 14600 35640 14634
rect 35674 14600 35730 14634
rect 35764 14600 35820 14634
rect 35854 14600 35910 14634
rect 35944 14600 36000 14634
rect 36034 14600 36111 14634
rect 35149 14581 36111 14600
rect 35149 14577 35221 14581
rect 35149 14543 35168 14577
rect 35202 14543 35221 14577
rect 35149 14487 35221 14543
rect 36039 14558 36111 14581
rect 36039 14524 36058 14558
rect 36092 14524 36111 14558
rect 35149 14453 35168 14487
rect 35202 14453 35221 14487
rect 35149 14397 35221 14453
rect 35149 14363 35168 14397
rect 35202 14363 35221 14397
rect 35149 14307 35221 14363
rect 35149 14273 35168 14307
rect 35202 14273 35221 14307
rect 35149 14217 35221 14273
rect 35149 14183 35168 14217
rect 35202 14183 35221 14217
rect 35149 14127 35221 14183
rect 35149 14093 35168 14127
rect 35202 14093 35221 14127
rect 35149 14037 35221 14093
rect 35149 14003 35168 14037
rect 35202 14003 35221 14037
rect 35149 13947 35221 14003
rect 35149 13913 35168 13947
rect 35202 13913 35221 13947
rect 35149 13857 35221 13913
rect 35149 13823 35168 13857
rect 35202 13823 35221 13857
rect 36039 14468 36111 14524
rect 36039 14434 36058 14468
rect 36092 14434 36111 14468
rect 36039 14378 36111 14434
rect 36039 14344 36058 14378
rect 36092 14344 36111 14378
rect 36039 14288 36111 14344
rect 36039 14254 36058 14288
rect 36092 14254 36111 14288
rect 36039 14198 36111 14254
rect 36039 14164 36058 14198
rect 36092 14164 36111 14198
rect 36039 14108 36111 14164
rect 36039 14074 36058 14108
rect 36092 14074 36111 14108
rect 36039 14018 36111 14074
rect 36039 13984 36058 14018
rect 36092 13984 36111 14018
rect 36039 13928 36111 13984
rect 36039 13894 36058 13928
rect 36092 13894 36111 13928
rect 36039 13838 36111 13894
rect 35149 13763 35221 13823
rect 36039 13804 36058 13838
rect 36092 13804 36111 13838
rect 36039 13763 36111 13804
rect 35149 13744 36111 13763
rect 35149 13710 35246 13744
rect 35280 13710 35336 13744
rect 35370 13710 35426 13744
rect 35460 13710 35516 13744
rect 35550 13710 35606 13744
rect 35640 13710 35696 13744
rect 35730 13710 35786 13744
rect 35820 13710 35876 13744
rect 35910 13710 35966 13744
rect 36000 13710 36111 13744
rect 35149 13691 36111 13710
rect 36489 14634 37451 14653
rect 36489 14600 36620 14634
rect 36654 14600 36710 14634
rect 36744 14600 36800 14634
rect 36834 14600 36890 14634
rect 36924 14600 36980 14634
rect 37014 14600 37070 14634
rect 37104 14600 37160 14634
rect 37194 14600 37250 14634
rect 37284 14600 37340 14634
rect 37374 14600 37451 14634
rect 36489 14581 37451 14600
rect 36489 14577 36561 14581
rect 36489 14543 36508 14577
rect 36542 14543 36561 14577
rect 36489 14487 36561 14543
rect 37379 14558 37451 14581
rect 37379 14524 37398 14558
rect 37432 14524 37451 14558
rect 36489 14453 36508 14487
rect 36542 14453 36561 14487
rect 36489 14397 36561 14453
rect 36489 14363 36508 14397
rect 36542 14363 36561 14397
rect 36489 14307 36561 14363
rect 36489 14273 36508 14307
rect 36542 14273 36561 14307
rect 36489 14217 36561 14273
rect 36489 14183 36508 14217
rect 36542 14183 36561 14217
rect 36489 14127 36561 14183
rect 36489 14093 36508 14127
rect 36542 14093 36561 14127
rect 36489 14037 36561 14093
rect 36489 14003 36508 14037
rect 36542 14003 36561 14037
rect 36489 13947 36561 14003
rect 36489 13913 36508 13947
rect 36542 13913 36561 13947
rect 36489 13857 36561 13913
rect 36489 13823 36508 13857
rect 36542 13823 36561 13857
rect 37379 14468 37451 14524
rect 37379 14434 37398 14468
rect 37432 14434 37451 14468
rect 37379 14378 37451 14434
rect 37379 14344 37398 14378
rect 37432 14344 37451 14378
rect 37379 14288 37451 14344
rect 37379 14254 37398 14288
rect 37432 14254 37451 14288
rect 37379 14198 37451 14254
rect 37379 14164 37398 14198
rect 37432 14164 37451 14198
rect 37379 14108 37451 14164
rect 37379 14074 37398 14108
rect 37432 14074 37451 14108
rect 37379 14018 37451 14074
rect 37379 13984 37398 14018
rect 37432 13984 37451 14018
rect 37379 13928 37451 13984
rect 37379 13894 37398 13928
rect 37432 13894 37451 13928
rect 37379 13838 37451 13894
rect 36489 13763 36561 13823
rect 37379 13804 37398 13838
rect 37432 13804 37451 13838
rect 37379 13763 37451 13804
rect 36489 13744 37451 13763
rect 36489 13710 36586 13744
rect 36620 13710 36676 13744
rect 36710 13710 36766 13744
rect 36800 13710 36856 13744
rect 36890 13710 36946 13744
rect 36980 13710 37036 13744
rect 37070 13710 37126 13744
rect 37160 13710 37216 13744
rect 37250 13710 37306 13744
rect 37340 13710 37451 13744
rect 36489 13691 37451 13710
rect 37829 14634 38791 14653
rect 37829 14600 37960 14634
rect 37994 14600 38050 14634
rect 38084 14600 38140 14634
rect 38174 14600 38230 14634
rect 38264 14600 38320 14634
rect 38354 14600 38410 14634
rect 38444 14600 38500 14634
rect 38534 14600 38590 14634
rect 38624 14600 38680 14634
rect 38714 14600 38791 14634
rect 37829 14581 38791 14600
rect 37829 14577 37901 14581
rect 37829 14543 37848 14577
rect 37882 14543 37901 14577
rect 37829 14487 37901 14543
rect 38719 14558 38791 14581
rect 38719 14524 38738 14558
rect 38772 14524 38791 14558
rect 37829 14453 37848 14487
rect 37882 14453 37901 14487
rect 37829 14397 37901 14453
rect 37829 14363 37848 14397
rect 37882 14363 37901 14397
rect 37829 14307 37901 14363
rect 37829 14273 37848 14307
rect 37882 14273 37901 14307
rect 37829 14217 37901 14273
rect 37829 14183 37848 14217
rect 37882 14183 37901 14217
rect 37829 14127 37901 14183
rect 37829 14093 37848 14127
rect 37882 14093 37901 14127
rect 37829 14037 37901 14093
rect 37829 14003 37848 14037
rect 37882 14003 37901 14037
rect 37829 13947 37901 14003
rect 37829 13913 37848 13947
rect 37882 13913 37901 13947
rect 37829 13857 37901 13913
rect 37829 13823 37848 13857
rect 37882 13823 37901 13857
rect 38719 14468 38791 14524
rect 38719 14434 38738 14468
rect 38772 14434 38791 14468
rect 38719 14378 38791 14434
rect 38719 14344 38738 14378
rect 38772 14344 38791 14378
rect 38719 14288 38791 14344
rect 38719 14254 38738 14288
rect 38772 14254 38791 14288
rect 38719 14198 38791 14254
rect 38719 14164 38738 14198
rect 38772 14164 38791 14198
rect 38719 14108 38791 14164
rect 38719 14074 38738 14108
rect 38772 14074 38791 14108
rect 38719 14018 38791 14074
rect 38719 13984 38738 14018
rect 38772 13984 38791 14018
rect 38719 13928 38791 13984
rect 38719 13894 38738 13928
rect 38772 13894 38791 13928
rect 38719 13838 38791 13894
rect 37829 13763 37901 13823
rect 38719 13804 38738 13838
rect 38772 13804 38791 13838
rect 38719 13763 38791 13804
rect 37829 13744 38791 13763
rect 37829 13710 37926 13744
rect 37960 13710 38016 13744
rect 38050 13710 38106 13744
rect 38140 13710 38196 13744
rect 38230 13710 38286 13744
rect 38320 13710 38376 13744
rect 38410 13710 38466 13744
rect 38500 13710 38556 13744
rect 38590 13710 38646 13744
rect 38680 13710 38791 13744
rect 37829 13691 38791 13710
<< psubdiffcont >>
rect 5927 39675 5961 39709
rect 30084 37284 30118 37318
rect 30180 37307 30214 37341
rect 30270 37307 30304 37341
rect 30360 37307 30394 37341
rect 30450 37307 30484 37341
rect 30540 37307 30574 37341
rect 30630 37307 30664 37341
rect 30720 37307 30754 37341
rect 30810 37307 30844 37341
rect 30900 37307 30934 37341
rect 30990 37307 31024 37341
rect 31080 37307 31114 37341
rect 31170 37307 31204 37341
rect 31271 37284 31305 37318
rect 31424 37284 31458 37318
rect 31520 37307 31554 37341
rect 31610 37307 31644 37341
rect 31700 37307 31734 37341
rect 31790 37307 31824 37341
rect 31880 37307 31914 37341
rect 31970 37307 32004 37341
rect 32060 37307 32094 37341
rect 32150 37307 32184 37341
rect 32240 37307 32274 37341
rect 32330 37307 32364 37341
rect 32420 37307 32454 37341
rect 32510 37307 32544 37341
rect 32611 37284 32645 37318
rect 32764 37284 32798 37318
rect 32860 37307 32894 37341
rect 32950 37307 32984 37341
rect 33040 37307 33074 37341
rect 33130 37307 33164 37341
rect 33220 37307 33254 37341
rect 33310 37307 33344 37341
rect 33400 37307 33434 37341
rect 33490 37307 33524 37341
rect 33580 37307 33614 37341
rect 33670 37307 33704 37341
rect 33760 37307 33794 37341
rect 33850 37307 33884 37341
rect 33951 37284 33985 37318
rect 34104 37284 34138 37318
rect 34200 37307 34234 37341
rect 34290 37307 34324 37341
rect 34380 37307 34414 37341
rect 34470 37307 34504 37341
rect 34560 37307 34594 37341
rect 34650 37307 34684 37341
rect 34740 37307 34774 37341
rect 34830 37307 34864 37341
rect 34920 37307 34954 37341
rect 35010 37307 35044 37341
rect 35100 37307 35134 37341
rect 35190 37307 35224 37341
rect 35291 37284 35325 37318
rect 35444 37284 35478 37318
rect 35540 37307 35574 37341
rect 35630 37307 35664 37341
rect 35720 37307 35754 37341
rect 35810 37307 35844 37341
rect 35900 37307 35934 37341
rect 35990 37307 36024 37341
rect 36080 37307 36114 37341
rect 36170 37307 36204 37341
rect 36260 37307 36294 37341
rect 36350 37307 36384 37341
rect 36440 37307 36474 37341
rect 36530 37307 36564 37341
rect 36631 37284 36665 37318
rect 36784 37284 36818 37318
rect 36880 37307 36914 37341
rect 36970 37307 37004 37341
rect 37060 37307 37094 37341
rect 37150 37307 37184 37341
rect 37240 37307 37274 37341
rect 37330 37307 37364 37341
rect 37420 37307 37454 37341
rect 37510 37307 37544 37341
rect 37600 37307 37634 37341
rect 37690 37307 37724 37341
rect 37780 37307 37814 37341
rect 37870 37307 37904 37341
rect 37971 37284 38005 37318
rect 38124 37284 38158 37318
rect 38220 37307 38254 37341
rect 38310 37307 38344 37341
rect 38400 37307 38434 37341
rect 38490 37307 38524 37341
rect 38580 37307 38614 37341
rect 38670 37307 38704 37341
rect 38760 37307 38794 37341
rect 38850 37307 38884 37341
rect 38940 37307 38974 37341
rect 39030 37307 39064 37341
rect 39120 37307 39154 37341
rect 39210 37307 39244 37341
rect 39311 37284 39345 37318
rect 30084 37194 30118 37228
rect 30084 37104 30118 37138
rect 30084 37014 30118 37048
rect 30084 36924 30118 36958
rect 30084 36834 30118 36868
rect 30084 36744 30118 36778
rect 30084 36654 30118 36688
rect 30084 36564 30118 36598
rect 30084 36474 30118 36508
rect 30084 36384 30118 36418
rect 30084 36294 30118 36328
rect 31271 37194 31305 37228
rect 31424 37194 31458 37228
rect 31271 37104 31305 37138
rect 31424 37104 31458 37138
rect 31271 37014 31305 37048
rect 31424 37014 31458 37048
rect 31271 36924 31305 36958
rect 31424 36924 31458 36958
rect 31271 36834 31305 36868
rect 31424 36834 31458 36868
rect 31271 36744 31305 36778
rect 31424 36744 31458 36778
rect 31271 36654 31305 36688
rect 31424 36654 31458 36688
rect 31271 36564 31305 36598
rect 31424 36564 31458 36598
rect 31271 36474 31305 36508
rect 31424 36474 31458 36508
rect 31271 36384 31305 36418
rect 31424 36384 31458 36418
rect 31271 36294 31305 36328
rect 31424 36294 31458 36328
rect 30084 36204 30118 36238
rect 32611 37194 32645 37228
rect 32764 37194 32798 37228
rect 32611 37104 32645 37138
rect 32764 37104 32798 37138
rect 32611 37014 32645 37048
rect 32764 37014 32798 37048
rect 32611 36924 32645 36958
rect 32764 36924 32798 36958
rect 32611 36834 32645 36868
rect 32764 36834 32798 36868
rect 32611 36744 32645 36778
rect 32764 36744 32798 36778
rect 32611 36654 32645 36688
rect 32764 36654 32798 36688
rect 32611 36564 32645 36598
rect 32764 36564 32798 36598
rect 32611 36474 32645 36508
rect 32764 36474 32798 36508
rect 32611 36384 32645 36418
rect 32764 36384 32798 36418
rect 32611 36294 32645 36328
rect 32764 36294 32798 36328
rect 31271 36204 31305 36238
rect 31424 36204 31458 36238
rect 33951 37194 33985 37228
rect 34104 37194 34138 37228
rect 33951 37104 33985 37138
rect 34104 37104 34138 37138
rect 33951 37014 33985 37048
rect 34104 37014 34138 37048
rect 33951 36924 33985 36958
rect 34104 36924 34138 36958
rect 33951 36834 33985 36868
rect 34104 36834 34138 36868
rect 33951 36744 33985 36778
rect 34104 36744 34138 36778
rect 33951 36654 33985 36688
rect 34104 36654 34138 36688
rect 33951 36564 33985 36598
rect 34104 36564 34138 36598
rect 33951 36474 33985 36508
rect 34104 36474 34138 36508
rect 33951 36384 33985 36418
rect 34104 36384 34138 36418
rect 33951 36294 33985 36328
rect 34104 36294 34138 36328
rect 32611 36204 32645 36238
rect 32764 36204 32798 36238
rect 35291 37194 35325 37228
rect 35444 37194 35478 37228
rect 35291 37104 35325 37138
rect 35444 37104 35478 37138
rect 35291 37014 35325 37048
rect 35444 37014 35478 37048
rect 35291 36924 35325 36958
rect 35444 36924 35478 36958
rect 35291 36834 35325 36868
rect 35444 36834 35478 36868
rect 35291 36744 35325 36778
rect 35444 36744 35478 36778
rect 35291 36654 35325 36688
rect 35444 36654 35478 36688
rect 35291 36564 35325 36598
rect 35444 36564 35478 36598
rect 35291 36474 35325 36508
rect 35444 36474 35478 36508
rect 35291 36384 35325 36418
rect 35444 36384 35478 36418
rect 35291 36294 35325 36328
rect 35444 36294 35478 36328
rect 33951 36204 33985 36238
rect 34104 36204 34138 36238
rect 36631 37194 36665 37228
rect 36784 37194 36818 37228
rect 36631 37104 36665 37138
rect 36784 37104 36818 37138
rect 36631 37014 36665 37048
rect 36784 37014 36818 37048
rect 36631 36924 36665 36958
rect 36784 36924 36818 36958
rect 36631 36834 36665 36868
rect 36784 36834 36818 36868
rect 36631 36744 36665 36778
rect 36784 36744 36818 36778
rect 36631 36654 36665 36688
rect 36784 36654 36818 36688
rect 36631 36564 36665 36598
rect 36784 36564 36818 36598
rect 36631 36474 36665 36508
rect 36784 36474 36818 36508
rect 36631 36384 36665 36418
rect 36784 36384 36818 36418
rect 36631 36294 36665 36328
rect 36784 36294 36818 36328
rect 35291 36204 35325 36238
rect 35444 36204 35478 36238
rect 37971 37194 38005 37228
rect 38124 37194 38158 37228
rect 37971 37104 38005 37138
rect 38124 37104 38158 37138
rect 37971 37014 38005 37048
rect 38124 37014 38158 37048
rect 37971 36924 38005 36958
rect 38124 36924 38158 36958
rect 37971 36834 38005 36868
rect 38124 36834 38158 36868
rect 37971 36744 38005 36778
rect 38124 36744 38158 36778
rect 37971 36654 38005 36688
rect 38124 36654 38158 36688
rect 37971 36564 38005 36598
rect 38124 36564 38158 36598
rect 37971 36474 38005 36508
rect 38124 36474 38158 36508
rect 37971 36384 38005 36418
rect 38124 36384 38158 36418
rect 37971 36294 38005 36328
rect 38124 36294 38158 36328
rect 36631 36204 36665 36238
rect 36784 36204 36818 36238
rect 39311 37194 39345 37228
rect 39311 37104 39345 37138
rect 39311 37014 39345 37048
rect 39311 36924 39345 36958
rect 39311 36834 39345 36868
rect 39311 36744 39345 36778
rect 39311 36654 39345 36688
rect 39311 36564 39345 36598
rect 40745 36621 41187 36723
rect 39311 36474 39345 36508
rect 39311 36384 39345 36418
rect 39311 36294 39345 36328
rect 37971 36204 38005 36238
rect 38124 36204 38158 36238
rect 39311 36204 39345 36238
rect 30180 36120 30214 36154
rect 30270 36120 30304 36154
rect 30360 36120 30394 36154
rect 30450 36120 30484 36154
rect 30540 36120 30574 36154
rect 30630 36120 30664 36154
rect 30720 36120 30754 36154
rect 30810 36120 30844 36154
rect 30900 36120 30934 36154
rect 30990 36120 31024 36154
rect 31080 36120 31114 36154
rect 31170 36120 31204 36154
rect 31520 36120 31554 36154
rect 31610 36120 31644 36154
rect 31700 36120 31734 36154
rect 31790 36120 31824 36154
rect 31880 36120 31914 36154
rect 31970 36120 32004 36154
rect 32060 36120 32094 36154
rect 32150 36120 32184 36154
rect 32240 36120 32274 36154
rect 32330 36120 32364 36154
rect 32420 36120 32454 36154
rect 32510 36120 32544 36154
rect 32860 36120 32894 36154
rect 32950 36120 32984 36154
rect 33040 36120 33074 36154
rect 33130 36120 33164 36154
rect 33220 36120 33254 36154
rect 33310 36120 33344 36154
rect 33400 36120 33434 36154
rect 33490 36120 33524 36154
rect 33580 36120 33614 36154
rect 33670 36120 33704 36154
rect 33760 36120 33794 36154
rect 33850 36120 33884 36154
rect 34200 36120 34234 36154
rect 34290 36120 34324 36154
rect 34380 36120 34414 36154
rect 34470 36120 34504 36154
rect 34560 36120 34594 36154
rect 34650 36120 34684 36154
rect 34740 36120 34774 36154
rect 34830 36120 34864 36154
rect 34920 36120 34954 36154
rect 35010 36120 35044 36154
rect 35100 36120 35134 36154
rect 35190 36120 35224 36154
rect 35540 36120 35574 36154
rect 35630 36120 35664 36154
rect 35720 36120 35754 36154
rect 35810 36120 35844 36154
rect 35900 36120 35934 36154
rect 35990 36120 36024 36154
rect 36080 36120 36114 36154
rect 36170 36120 36204 36154
rect 36260 36120 36294 36154
rect 36350 36120 36384 36154
rect 36440 36120 36474 36154
rect 36530 36120 36564 36154
rect 36880 36120 36914 36154
rect 36970 36120 37004 36154
rect 37060 36120 37094 36154
rect 37150 36120 37184 36154
rect 37240 36120 37274 36154
rect 37330 36120 37364 36154
rect 37420 36120 37454 36154
rect 37510 36120 37544 36154
rect 37600 36120 37634 36154
rect 37690 36120 37724 36154
rect 37780 36120 37814 36154
rect 37870 36120 37904 36154
rect 38220 36120 38254 36154
rect 38310 36120 38344 36154
rect 38400 36120 38434 36154
rect 38490 36120 38524 36154
rect 38580 36120 38614 36154
rect 38670 36120 38704 36154
rect 38760 36120 38794 36154
rect 38850 36120 38884 36154
rect 38940 36120 38974 36154
rect 39030 36120 39064 36154
rect 39120 36120 39154 36154
rect 39210 36120 39244 36154
rect 28271 35915 28305 35949
rect 38393 29101 38835 29203
rect 41137 29101 41579 29203
rect 7719 25341 8161 25443
rect 28320 26004 28354 26038
rect 28416 26027 28450 26061
rect 28506 26027 28540 26061
rect 28596 26027 28630 26061
rect 28686 26027 28720 26061
rect 28776 26027 28810 26061
rect 28866 26027 28900 26061
rect 28956 26027 28990 26061
rect 29046 26027 29080 26061
rect 29136 26027 29170 26061
rect 29226 26027 29260 26061
rect 29316 26027 29350 26061
rect 29406 26027 29440 26061
rect 29507 26004 29541 26038
rect 29660 26004 29694 26038
rect 29756 26027 29790 26061
rect 29846 26027 29880 26061
rect 29936 26027 29970 26061
rect 30026 26027 30060 26061
rect 30116 26027 30150 26061
rect 30206 26027 30240 26061
rect 30296 26027 30330 26061
rect 30386 26027 30420 26061
rect 30476 26027 30510 26061
rect 30566 26027 30600 26061
rect 30656 26027 30690 26061
rect 30746 26027 30780 26061
rect 30847 26004 30881 26038
rect 31000 26004 31034 26038
rect 31096 26027 31130 26061
rect 31186 26027 31220 26061
rect 31276 26027 31310 26061
rect 31366 26027 31400 26061
rect 31456 26027 31490 26061
rect 31546 26027 31580 26061
rect 31636 26027 31670 26061
rect 31726 26027 31760 26061
rect 31816 26027 31850 26061
rect 31906 26027 31940 26061
rect 31996 26027 32030 26061
rect 32086 26027 32120 26061
rect 32187 26004 32221 26038
rect 32340 26004 32374 26038
rect 32436 26027 32470 26061
rect 32526 26027 32560 26061
rect 32616 26027 32650 26061
rect 32706 26027 32740 26061
rect 32796 26027 32830 26061
rect 32886 26027 32920 26061
rect 32976 26027 33010 26061
rect 33066 26027 33100 26061
rect 33156 26027 33190 26061
rect 33246 26027 33280 26061
rect 33336 26027 33370 26061
rect 33426 26027 33460 26061
rect 33527 26004 33561 26038
rect 33680 26004 33714 26038
rect 33776 26027 33810 26061
rect 33866 26027 33900 26061
rect 33956 26027 33990 26061
rect 34046 26027 34080 26061
rect 34136 26027 34170 26061
rect 34226 26027 34260 26061
rect 34316 26027 34350 26061
rect 34406 26027 34440 26061
rect 34496 26027 34530 26061
rect 34586 26027 34620 26061
rect 34676 26027 34710 26061
rect 34766 26027 34800 26061
rect 34867 26004 34901 26038
rect 35020 26004 35054 26038
rect 35116 26027 35150 26061
rect 35206 26027 35240 26061
rect 35296 26027 35330 26061
rect 35386 26027 35420 26061
rect 35476 26027 35510 26061
rect 35566 26027 35600 26061
rect 35656 26027 35690 26061
rect 35746 26027 35780 26061
rect 35836 26027 35870 26061
rect 35926 26027 35960 26061
rect 36016 26027 36050 26061
rect 36106 26027 36140 26061
rect 36207 26004 36241 26038
rect 36360 26004 36394 26038
rect 36456 26027 36490 26061
rect 36546 26027 36580 26061
rect 36636 26027 36670 26061
rect 36726 26027 36760 26061
rect 36816 26027 36850 26061
rect 36906 26027 36940 26061
rect 36996 26027 37030 26061
rect 37086 26027 37120 26061
rect 37176 26027 37210 26061
rect 37266 26027 37300 26061
rect 37356 26027 37390 26061
rect 37446 26027 37480 26061
rect 37547 26004 37581 26038
rect 37700 26004 37734 26038
rect 37796 26027 37830 26061
rect 37886 26027 37920 26061
rect 37976 26027 38010 26061
rect 38066 26027 38100 26061
rect 38156 26027 38190 26061
rect 38246 26027 38280 26061
rect 38336 26027 38370 26061
rect 38426 26027 38460 26061
rect 38516 26027 38550 26061
rect 38606 26027 38640 26061
rect 38696 26027 38730 26061
rect 38786 26027 38820 26061
rect 38887 26004 38921 26038
rect 28320 25914 28354 25948
rect 28320 25824 28354 25858
rect 28320 25734 28354 25768
rect 28320 25644 28354 25678
rect 28320 25554 28354 25588
rect 28320 25464 28354 25498
rect 28320 25374 28354 25408
rect 28320 25284 28354 25318
rect 28320 25194 28354 25228
rect 28320 25104 28354 25138
rect 28320 25014 28354 25048
rect 29507 25914 29541 25948
rect 29660 25914 29694 25948
rect 29507 25824 29541 25858
rect 29660 25824 29694 25858
rect 29507 25734 29541 25768
rect 29660 25734 29694 25768
rect 29507 25644 29541 25678
rect 29660 25644 29694 25678
rect 29507 25554 29541 25588
rect 29660 25554 29694 25588
rect 29507 25464 29541 25498
rect 29660 25464 29694 25498
rect 29507 25374 29541 25408
rect 29660 25374 29694 25408
rect 29507 25284 29541 25318
rect 29660 25284 29694 25318
rect 29507 25194 29541 25228
rect 29660 25194 29694 25228
rect 29507 25104 29541 25138
rect 29660 25104 29694 25138
rect 29507 25014 29541 25048
rect 29660 25014 29694 25048
rect 28320 24924 28354 24958
rect 30847 25914 30881 25948
rect 31000 25914 31034 25948
rect 30847 25824 30881 25858
rect 31000 25824 31034 25858
rect 30847 25734 30881 25768
rect 31000 25734 31034 25768
rect 30847 25644 30881 25678
rect 31000 25644 31034 25678
rect 30847 25554 30881 25588
rect 31000 25554 31034 25588
rect 30847 25464 30881 25498
rect 31000 25464 31034 25498
rect 30847 25374 30881 25408
rect 31000 25374 31034 25408
rect 30847 25284 30881 25318
rect 31000 25284 31034 25318
rect 30847 25194 30881 25228
rect 31000 25194 31034 25228
rect 30847 25104 30881 25138
rect 31000 25104 31034 25138
rect 30847 25014 30881 25048
rect 31000 25014 31034 25048
rect 29507 24924 29541 24958
rect 29660 24924 29694 24958
rect 32187 25914 32221 25948
rect 32340 25914 32374 25948
rect 32187 25824 32221 25858
rect 32340 25824 32374 25858
rect 32187 25734 32221 25768
rect 32340 25734 32374 25768
rect 32187 25644 32221 25678
rect 32340 25644 32374 25678
rect 32187 25554 32221 25588
rect 32340 25554 32374 25588
rect 32187 25464 32221 25498
rect 32340 25464 32374 25498
rect 32187 25374 32221 25408
rect 32340 25374 32374 25408
rect 32187 25284 32221 25318
rect 32340 25284 32374 25318
rect 32187 25194 32221 25228
rect 32340 25194 32374 25228
rect 32187 25104 32221 25138
rect 32340 25104 32374 25138
rect 32187 25014 32221 25048
rect 32340 25014 32374 25048
rect 30847 24924 30881 24958
rect 31000 24924 31034 24958
rect 33527 25914 33561 25948
rect 33680 25914 33714 25948
rect 33527 25824 33561 25858
rect 33680 25824 33714 25858
rect 33527 25734 33561 25768
rect 33680 25734 33714 25768
rect 33527 25644 33561 25678
rect 33680 25644 33714 25678
rect 33527 25554 33561 25588
rect 33680 25554 33714 25588
rect 33527 25464 33561 25498
rect 33680 25464 33714 25498
rect 33527 25374 33561 25408
rect 33680 25374 33714 25408
rect 33527 25284 33561 25318
rect 33680 25284 33714 25318
rect 33527 25194 33561 25228
rect 33680 25194 33714 25228
rect 33527 25104 33561 25138
rect 33680 25104 33714 25138
rect 33527 25014 33561 25048
rect 33680 25014 33714 25048
rect 32187 24924 32221 24958
rect 32340 24924 32374 24958
rect 34867 25914 34901 25948
rect 35020 25914 35054 25948
rect 34867 25824 34901 25858
rect 35020 25824 35054 25858
rect 34867 25734 34901 25768
rect 35020 25734 35054 25768
rect 34867 25644 34901 25678
rect 35020 25644 35054 25678
rect 34867 25554 34901 25588
rect 35020 25554 35054 25588
rect 34867 25464 34901 25498
rect 35020 25464 35054 25498
rect 34867 25374 34901 25408
rect 35020 25374 35054 25408
rect 34867 25284 34901 25318
rect 35020 25284 35054 25318
rect 34867 25194 34901 25228
rect 35020 25194 35054 25228
rect 34867 25104 34901 25138
rect 35020 25104 35054 25138
rect 34867 25014 34901 25048
rect 35020 25014 35054 25048
rect 33527 24924 33561 24958
rect 33680 24924 33714 24958
rect 36207 25914 36241 25948
rect 36360 25914 36394 25948
rect 36207 25824 36241 25858
rect 36360 25824 36394 25858
rect 36207 25734 36241 25768
rect 36360 25734 36394 25768
rect 36207 25644 36241 25678
rect 36360 25644 36394 25678
rect 36207 25554 36241 25588
rect 36360 25554 36394 25588
rect 36207 25464 36241 25498
rect 36360 25464 36394 25498
rect 36207 25374 36241 25408
rect 36360 25374 36394 25408
rect 36207 25284 36241 25318
rect 36360 25284 36394 25318
rect 36207 25194 36241 25228
rect 36360 25194 36394 25228
rect 36207 25104 36241 25138
rect 36360 25104 36394 25138
rect 36207 25014 36241 25048
rect 36360 25014 36394 25048
rect 34867 24924 34901 24958
rect 35020 24924 35054 24958
rect 37547 25914 37581 25948
rect 37700 25914 37734 25948
rect 37547 25824 37581 25858
rect 37700 25824 37734 25858
rect 37547 25734 37581 25768
rect 37700 25734 37734 25768
rect 37547 25644 37581 25678
rect 37700 25644 37734 25678
rect 37547 25554 37581 25588
rect 37700 25554 37734 25588
rect 37547 25464 37581 25498
rect 37700 25464 37734 25498
rect 37547 25374 37581 25408
rect 37700 25374 37734 25408
rect 37547 25284 37581 25318
rect 37700 25284 37734 25318
rect 37547 25194 37581 25228
rect 37700 25194 37734 25228
rect 37547 25104 37581 25138
rect 37700 25104 37734 25138
rect 37547 25014 37581 25048
rect 37700 25014 37734 25048
rect 36207 24924 36241 24958
rect 36360 24924 36394 24958
rect 38887 25914 38921 25948
rect 38887 25824 38921 25858
rect 38887 25734 38921 25768
rect 38887 25644 38921 25678
rect 38887 25554 38921 25588
rect 38887 25464 38921 25498
rect 38887 25374 38921 25408
rect 38887 25284 38921 25318
rect 40745 25341 41187 25443
rect 38887 25194 38921 25228
rect 38887 25104 38921 25138
rect 38887 25014 38921 25048
rect 37547 24924 37581 24958
rect 37700 24924 37734 24958
rect 38887 24924 38921 24958
rect 28416 24840 28450 24874
rect 28506 24840 28540 24874
rect 28596 24840 28630 24874
rect 28686 24840 28720 24874
rect 28776 24840 28810 24874
rect 28866 24840 28900 24874
rect 28956 24840 28990 24874
rect 29046 24840 29080 24874
rect 29136 24840 29170 24874
rect 29226 24840 29260 24874
rect 29316 24840 29350 24874
rect 29406 24840 29440 24874
rect 29756 24840 29790 24874
rect 29846 24840 29880 24874
rect 29936 24840 29970 24874
rect 30026 24840 30060 24874
rect 30116 24840 30150 24874
rect 30206 24840 30240 24874
rect 30296 24840 30330 24874
rect 30386 24840 30420 24874
rect 30476 24840 30510 24874
rect 30566 24840 30600 24874
rect 30656 24840 30690 24874
rect 30746 24840 30780 24874
rect 31096 24840 31130 24874
rect 31186 24840 31220 24874
rect 31276 24840 31310 24874
rect 31366 24840 31400 24874
rect 31456 24840 31490 24874
rect 31546 24840 31580 24874
rect 31636 24840 31670 24874
rect 31726 24840 31760 24874
rect 31816 24840 31850 24874
rect 31906 24840 31940 24874
rect 31996 24840 32030 24874
rect 32086 24840 32120 24874
rect 32436 24840 32470 24874
rect 32526 24840 32560 24874
rect 32616 24840 32650 24874
rect 32706 24840 32740 24874
rect 32796 24840 32830 24874
rect 32886 24840 32920 24874
rect 32976 24840 33010 24874
rect 33066 24840 33100 24874
rect 33156 24840 33190 24874
rect 33246 24840 33280 24874
rect 33336 24840 33370 24874
rect 33426 24840 33460 24874
rect 33776 24840 33810 24874
rect 33866 24840 33900 24874
rect 33956 24840 33990 24874
rect 34046 24840 34080 24874
rect 34136 24840 34170 24874
rect 34226 24840 34260 24874
rect 34316 24840 34350 24874
rect 34406 24840 34440 24874
rect 34496 24840 34530 24874
rect 34586 24840 34620 24874
rect 34676 24840 34710 24874
rect 34766 24840 34800 24874
rect 35116 24840 35150 24874
rect 35206 24840 35240 24874
rect 35296 24840 35330 24874
rect 35386 24840 35420 24874
rect 35476 24840 35510 24874
rect 35566 24840 35600 24874
rect 35656 24840 35690 24874
rect 35746 24840 35780 24874
rect 35836 24840 35870 24874
rect 35926 24840 35960 24874
rect 36016 24840 36050 24874
rect 36106 24840 36140 24874
rect 36456 24840 36490 24874
rect 36546 24840 36580 24874
rect 36636 24840 36670 24874
rect 36726 24840 36760 24874
rect 36816 24840 36850 24874
rect 36906 24840 36940 24874
rect 36996 24840 37030 24874
rect 37086 24840 37120 24874
rect 37176 24840 37210 24874
rect 37266 24840 37300 24874
rect 37356 24840 37390 24874
rect 37446 24840 37480 24874
rect 37796 24840 37830 24874
rect 37886 24840 37920 24874
rect 37976 24840 38010 24874
rect 38066 24840 38100 24874
rect 38156 24840 38190 24874
rect 38246 24840 38280 24874
rect 38336 24840 38370 24874
rect 38426 24840 38460 24874
rect 38516 24840 38550 24874
rect 38606 24840 38640 24874
rect 38696 24840 38730 24874
rect 38786 24840 38820 24874
rect 22911 24635 22945 24669
rect 24013 24605 24047 24639
rect 25313 24605 25347 24639
rect 21068 22244 21102 22278
rect 21164 22267 21198 22301
rect 21254 22267 21288 22301
rect 21344 22267 21378 22301
rect 21434 22267 21468 22301
rect 21524 22267 21558 22301
rect 21614 22267 21648 22301
rect 21704 22267 21738 22301
rect 21794 22267 21828 22301
rect 21884 22267 21918 22301
rect 21974 22267 22008 22301
rect 22064 22267 22098 22301
rect 22154 22267 22188 22301
rect 22255 22244 22289 22278
rect 21068 22154 21102 22188
rect 21068 22064 21102 22098
rect 21068 21974 21102 22008
rect 21068 21884 21102 21918
rect 21068 21794 21102 21828
rect 21068 21704 21102 21738
rect 21068 21614 21102 21648
rect 21068 21524 21102 21558
rect 21068 21434 21102 21468
rect 21068 21344 21102 21378
rect 21068 21254 21102 21288
rect 22255 22154 22289 22188
rect 28320 22244 28354 22278
rect 28416 22267 28450 22301
rect 28506 22267 28540 22301
rect 28596 22267 28630 22301
rect 28686 22267 28720 22301
rect 28776 22267 28810 22301
rect 28866 22267 28900 22301
rect 28956 22267 28990 22301
rect 29046 22267 29080 22301
rect 29136 22267 29170 22301
rect 29226 22267 29260 22301
rect 29316 22267 29350 22301
rect 29406 22267 29440 22301
rect 29507 22244 29541 22278
rect 29660 22244 29694 22278
rect 29756 22267 29790 22301
rect 29846 22267 29880 22301
rect 29936 22267 29970 22301
rect 30026 22267 30060 22301
rect 30116 22267 30150 22301
rect 30206 22267 30240 22301
rect 30296 22267 30330 22301
rect 30386 22267 30420 22301
rect 30476 22267 30510 22301
rect 30566 22267 30600 22301
rect 30656 22267 30690 22301
rect 30746 22267 30780 22301
rect 30847 22244 30881 22278
rect 31000 22244 31034 22278
rect 31096 22267 31130 22301
rect 31186 22267 31220 22301
rect 31276 22267 31310 22301
rect 31366 22267 31400 22301
rect 31456 22267 31490 22301
rect 31546 22267 31580 22301
rect 31636 22267 31670 22301
rect 31726 22267 31760 22301
rect 31816 22267 31850 22301
rect 31906 22267 31940 22301
rect 31996 22267 32030 22301
rect 32086 22267 32120 22301
rect 32187 22244 32221 22278
rect 32340 22244 32374 22278
rect 32436 22267 32470 22301
rect 32526 22267 32560 22301
rect 32616 22267 32650 22301
rect 32706 22267 32740 22301
rect 32796 22267 32830 22301
rect 32886 22267 32920 22301
rect 32976 22267 33010 22301
rect 33066 22267 33100 22301
rect 33156 22267 33190 22301
rect 33246 22267 33280 22301
rect 33336 22267 33370 22301
rect 33426 22267 33460 22301
rect 33527 22244 33561 22278
rect 33680 22244 33714 22278
rect 33776 22267 33810 22301
rect 33866 22267 33900 22301
rect 33956 22267 33990 22301
rect 34046 22267 34080 22301
rect 34136 22267 34170 22301
rect 34226 22267 34260 22301
rect 34316 22267 34350 22301
rect 34406 22267 34440 22301
rect 34496 22267 34530 22301
rect 34586 22267 34620 22301
rect 34676 22267 34710 22301
rect 34766 22267 34800 22301
rect 34867 22244 34901 22278
rect 35020 22244 35054 22278
rect 35116 22267 35150 22301
rect 35206 22267 35240 22301
rect 35296 22267 35330 22301
rect 35386 22267 35420 22301
rect 35476 22267 35510 22301
rect 35566 22267 35600 22301
rect 35656 22267 35690 22301
rect 35746 22267 35780 22301
rect 35836 22267 35870 22301
rect 35926 22267 35960 22301
rect 36016 22267 36050 22301
rect 36106 22267 36140 22301
rect 36207 22244 36241 22278
rect 36360 22244 36394 22278
rect 36456 22267 36490 22301
rect 36546 22267 36580 22301
rect 36636 22267 36670 22301
rect 36726 22267 36760 22301
rect 36816 22267 36850 22301
rect 36906 22267 36940 22301
rect 36996 22267 37030 22301
rect 37086 22267 37120 22301
rect 37176 22267 37210 22301
rect 37266 22267 37300 22301
rect 37356 22267 37390 22301
rect 37446 22267 37480 22301
rect 37547 22244 37581 22278
rect 37700 22244 37734 22278
rect 37796 22267 37830 22301
rect 37886 22267 37920 22301
rect 37976 22267 38010 22301
rect 38066 22267 38100 22301
rect 38156 22267 38190 22301
rect 38246 22267 38280 22301
rect 38336 22267 38370 22301
rect 38426 22267 38460 22301
rect 38516 22267 38550 22301
rect 38606 22267 38640 22301
rect 38696 22267 38730 22301
rect 38786 22267 38820 22301
rect 38887 22244 38921 22278
rect 28320 22154 28354 22188
rect 22255 22064 22289 22098
rect 22255 21974 22289 22008
rect 22255 21884 22289 21918
rect 22255 21794 22289 21828
rect 22255 21704 22289 21738
rect 22255 21614 22289 21648
rect 22255 21524 22289 21558
rect 22255 21434 22289 21468
rect 22255 21344 22289 21378
rect 28320 22064 28354 22098
rect 28320 21974 28354 22008
rect 28320 21884 28354 21918
rect 28320 21794 28354 21828
rect 28320 21704 28354 21738
rect 28320 21614 28354 21648
rect 28320 21524 28354 21558
rect 28320 21434 28354 21468
rect 28320 21344 28354 21378
rect 22255 21254 22289 21288
rect 21068 21164 21102 21198
rect 22255 21164 22289 21198
rect 28320 21254 28354 21288
rect 29507 22154 29541 22188
rect 29660 22154 29694 22188
rect 29507 22064 29541 22098
rect 29660 22064 29694 22098
rect 29507 21974 29541 22008
rect 29660 21974 29694 22008
rect 29507 21884 29541 21918
rect 29660 21884 29694 21918
rect 29507 21794 29541 21828
rect 29660 21794 29694 21828
rect 29507 21704 29541 21738
rect 29660 21704 29694 21738
rect 29507 21614 29541 21648
rect 29660 21614 29694 21648
rect 29507 21524 29541 21558
rect 29660 21524 29694 21558
rect 29507 21434 29541 21468
rect 29660 21434 29694 21468
rect 29507 21344 29541 21378
rect 29660 21344 29694 21378
rect 29507 21254 29541 21288
rect 29660 21254 29694 21288
rect 28320 21164 28354 21198
rect 30847 22154 30881 22188
rect 31000 22154 31034 22188
rect 30847 22064 30881 22098
rect 31000 22064 31034 22098
rect 30847 21974 30881 22008
rect 31000 21974 31034 22008
rect 30847 21884 30881 21918
rect 31000 21884 31034 21918
rect 30847 21794 30881 21828
rect 31000 21794 31034 21828
rect 30847 21704 30881 21738
rect 31000 21704 31034 21738
rect 30847 21614 30881 21648
rect 31000 21614 31034 21648
rect 30847 21524 30881 21558
rect 31000 21524 31034 21558
rect 30847 21434 30881 21468
rect 31000 21434 31034 21468
rect 30847 21344 30881 21378
rect 31000 21344 31034 21378
rect 30847 21254 30881 21288
rect 31000 21254 31034 21288
rect 29507 21164 29541 21198
rect 29660 21164 29694 21198
rect 32187 22154 32221 22188
rect 32340 22154 32374 22188
rect 32187 22064 32221 22098
rect 32340 22064 32374 22098
rect 32187 21974 32221 22008
rect 32340 21974 32374 22008
rect 32187 21884 32221 21918
rect 32340 21884 32374 21918
rect 32187 21794 32221 21828
rect 32340 21794 32374 21828
rect 32187 21704 32221 21738
rect 32340 21704 32374 21738
rect 32187 21614 32221 21648
rect 32340 21614 32374 21648
rect 32187 21524 32221 21558
rect 32340 21524 32374 21558
rect 32187 21434 32221 21468
rect 32340 21434 32374 21468
rect 32187 21344 32221 21378
rect 32340 21344 32374 21378
rect 32187 21254 32221 21288
rect 32340 21254 32374 21288
rect 30847 21164 30881 21198
rect 31000 21164 31034 21198
rect 33527 22154 33561 22188
rect 33680 22154 33714 22188
rect 33527 22064 33561 22098
rect 33680 22064 33714 22098
rect 33527 21974 33561 22008
rect 33680 21974 33714 22008
rect 33527 21884 33561 21918
rect 33680 21884 33714 21918
rect 33527 21794 33561 21828
rect 33680 21794 33714 21828
rect 33527 21704 33561 21738
rect 33680 21704 33714 21738
rect 33527 21614 33561 21648
rect 33680 21614 33714 21648
rect 33527 21524 33561 21558
rect 33680 21524 33714 21558
rect 33527 21434 33561 21468
rect 33680 21434 33714 21468
rect 33527 21344 33561 21378
rect 33680 21344 33714 21378
rect 33527 21254 33561 21288
rect 33680 21254 33714 21288
rect 32187 21164 32221 21198
rect 32340 21164 32374 21198
rect 34867 22154 34901 22188
rect 35020 22154 35054 22188
rect 34867 22064 34901 22098
rect 35020 22064 35054 22098
rect 34867 21974 34901 22008
rect 35020 21974 35054 22008
rect 34867 21884 34901 21918
rect 35020 21884 35054 21918
rect 34867 21794 34901 21828
rect 35020 21794 35054 21828
rect 34867 21704 34901 21738
rect 35020 21704 35054 21738
rect 34867 21614 34901 21648
rect 35020 21614 35054 21648
rect 34867 21524 34901 21558
rect 35020 21524 35054 21558
rect 34867 21434 34901 21468
rect 35020 21434 35054 21468
rect 34867 21344 34901 21378
rect 35020 21344 35054 21378
rect 34867 21254 34901 21288
rect 35020 21254 35054 21288
rect 33527 21164 33561 21198
rect 33680 21164 33714 21198
rect 36207 22154 36241 22188
rect 36360 22154 36394 22188
rect 36207 22064 36241 22098
rect 36360 22064 36394 22098
rect 36207 21974 36241 22008
rect 36360 21974 36394 22008
rect 36207 21884 36241 21918
rect 36360 21884 36394 21918
rect 36207 21794 36241 21828
rect 36360 21794 36394 21828
rect 36207 21704 36241 21738
rect 36360 21704 36394 21738
rect 36207 21614 36241 21648
rect 36360 21614 36394 21648
rect 36207 21524 36241 21558
rect 36360 21524 36394 21558
rect 36207 21434 36241 21468
rect 36360 21434 36394 21468
rect 36207 21344 36241 21378
rect 36360 21344 36394 21378
rect 36207 21254 36241 21288
rect 36360 21254 36394 21288
rect 34867 21164 34901 21198
rect 35020 21164 35054 21198
rect 37547 22154 37581 22188
rect 37700 22154 37734 22188
rect 37547 22064 37581 22098
rect 37700 22064 37734 22098
rect 37547 21974 37581 22008
rect 37700 21974 37734 22008
rect 37547 21884 37581 21918
rect 37700 21884 37734 21918
rect 37547 21794 37581 21828
rect 37700 21794 37734 21828
rect 37547 21704 37581 21738
rect 37700 21704 37734 21738
rect 37547 21614 37581 21648
rect 37700 21614 37734 21648
rect 37547 21524 37581 21558
rect 37700 21524 37734 21558
rect 37547 21434 37581 21468
rect 37700 21434 37734 21468
rect 37547 21344 37581 21378
rect 37700 21344 37734 21378
rect 37547 21254 37581 21288
rect 37700 21254 37734 21288
rect 36207 21164 36241 21198
rect 36360 21164 36394 21198
rect 38887 22154 38921 22188
rect 38887 22064 38921 22098
rect 38887 21974 38921 22008
rect 38887 21884 38921 21918
rect 38887 21794 38921 21828
rect 38887 21704 38921 21738
rect 38887 21614 38921 21648
rect 38887 21524 38921 21558
rect 40745 21581 41187 21683
rect 38887 21434 38921 21468
rect 38887 21344 38921 21378
rect 38887 21254 38921 21288
rect 37547 21164 37581 21198
rect 37700 21164 37734 21198
rect 38887 21164 38921 21198
rect 21164 21080 21198 21114
rect 21254 21080 21288 21114
rect 21344 21080 21378 21114
rect 21434 21080 21468 21114
rect 21524 21080 21558 21114
rect 21614 21080 21648 21114
rect 21704 21080 21738 21114
rect 21794 21080 21828 21114
rect 21884 21080 21918 21114
rect 21974 21080 22008 21114
rect 22064 21080 22098 21114
rect 22154 21080 22188 21114
rect 28416 21080 28450 21114
rect 28506 21080 28540 21114
rect 28596 21080 28630 21114
rect 28686 21080 28720 21114
rect 28776 21080 28810 21114
rect 28866 21080 28900 21114
rect 28956 21080 28990 21114
rect 29046 21080 29080 21114
rect 29136 21080 29170 21114
rect 29226 21080 29260 21114
rect 29316 21080 29350 21114
rect 29406 21080 29440 21114
rect 29756 21080 29790 21114
rect 29846 21080 29880 21114
rect 29936 21080 29970 21114
rect 30026 21080 30060 21114
rect 30116 21080 30150 21114
rect 30206 21080 30240 21114
rect 30296 21080 30330 21114
rect 30386 21080 30420 21114
rect 30476 21080 30510 21114
rect 30566 21080 30600 21114
rect 30656 21080 30690 21114
rect 30746 21080 30780 21114
rect 31096 21080 31130 21114
rect 31186 21080 31220 21114
rect 31276 21080 31310 21114
rect 31366 21080 31400 21114
rect 31456 21080 31490 21114
rect 31546 21080 31580 21114
rect 31636 21080 31670 21114
rect 31726 21080 31760 21114
rect 31816 21080 31850 21114
rect 31906 21080 31940 21114
rect 31996 21080 32030 21114
rect 32086 21080 32120 21114
rect 32436 21080 32470 21114
rect 32526 21080 32560 21114
rect 32616 21080 32650 21114
rect 32706 21080 32740 21114
rect 32796 21080 32830 21114
rect 32886 21080 32920 21114
rect 32976 21080 33010 21114
rect 33066 21080 33100 21114
rect 33156 21080 33190 21114
rect 33246 21080 33280 21114
rect 33336 21080 33370 21114
rect 33426 21080 33460 21114
rect 33776 21080 33810 21114
rect 33866 21080 33900 21114
rect 33956 21080 33990 21114
rect 34046 21080 34080 21114
rect 34136 21080 34170 21114
rect 34226 21080 34260 21114
rect 34316 21080 34350 21114
rect 34406 21080 34440 21114
rect 34496 21080 34530 21114
rect 34586 21080 34620 21114
rect 34676 21080 34710 21114
rect 34766 21080 34800 21114
rect 35116 21080 35150 21114
rect 35206 21080 35240 21114
rect 35296 21080 35330 21114
rect 35386 21080 35420 21114
rect 35476 21080 35510 21114
rect 35566 21080 35600 21114
rect 35656 21080 35690 21114
rect 35746 21080 35780 21114
rect 35836 21080 35870 21114
rect 35926 21080 35960 21114
rect 36016 21080 36050 21114
rect 36106 21080 36140 21114
rect 36456 21080 36490 21114
rect 36546 21080 36580 21114
rect 36636 21080 36670 21114
rect 36726 21080 36760 21114
rect 36816 21080 36850 21114
rect 36906 21080 36940 21114
rect 36996 21080 37030 21114
rect 37086 21080 37120 21114
rect 37176 21080 37210 21114
rect 37266 21080 37300 21114
rect 37356 21080 37390 21114
rect 37446 21080 37480 21114
rect 37796 21080 37830 21114
rect 37886 21080 37920 21114
rect 37976 21080 38010 21114
rect 38066 21080 38100 21114
rect 38156 21080 38190 21114
rect 38246 21080 38280 21114
rect 38336 21080 38370 21114
rect 38426 21080 38460 21114
rect 38516 21080 38550 21114
rect 38606 21080 38640 21114
rect 38696 21080 38730 21114
rect 38786 21080 38820 21114
rect 22911 20875 22945 20909
rect 24013 20845 24047 20879
rect 25313 20845 25347 20879
rect 11639 17821 12081 17923
rect 14383 17821 14825 17923
rect 5957 17115 5991 17149
rect 7059 17085 7093 17119
rect 8359 17085 8393 17119
rect 28320 18484 28354 18518
rect 28416 18507 28450 18541
rect 28506 18507 28540 18541
rect 28596 18507 28630 18541
rect 28686 18507 28720 18541
rect 28776 18507 28810 18541
rect 28866 18507 28900 18541
rect 28956 18507 28990 18541
rect 29046 18507 29080 18541
rect 29136 18507 29170 18541
rect 29226 18507 29260 18541
rect 29316 18507 29350 18541
rect 29406 18507 29440 18541
rect 29507 18484 29541 18518
rect 29660 18484 29694 18518
rect 29756 18507 29790 18541
rect 29846 18507 29880 18541
rect 29936 18507 29970 18541
rect 30026 18507 30060 18541
rect 30116 18507 30150 18541
rect 30206 18507 30240 18541
rect 30296 18507 30330 18541
rect 30386 18507 30420 18541
rect 30476 18507 30510 18541
rect 30566 18507 30600 18541
rect 30656 18507 30690 18541
rect 30746 18507 30780 18541
rect 30847 18484 30881 18518
rect 31000 18484 31034 18518
rect 31096 18507 31130 18541
rect 31186 18507 31220 18541
rect 31276 18507 31310 18541
rect 31366 18507 31400 18541
rect 31456 18507 31490 18541
rect 31546 18507 31580 18541
rect 31636 18507 31670 18541
rect 31726 18507 31760 18541
rect 31816 18507 31850 18541
rect 31906 18507 31940 18541
rect 31996 18507 32030 18541
rect 32086 18507 32120 18541
rect 32187 18484 32221 18518
rect 32340 18484 32374 18518
rect 32436 18507 32470 18541
rect 32526 18507 32560 18541
rect 32616 18507 32650 18541
rect 32706 18507 32740 18541
rect 32796 18507 32830 18541
rect 32886 18507 32920 18541
rect 32976 18507 33010 18541
rect 33066 18507 33100 18541
rect 33156 18507 33190 18541
rect 33246 18507 33280 18541
rect 33336 18507 33370 18541
rect 33426 18507 33460 18541
rect 33527 18484 33561 18518
rect 33680 18484 33714 18518
rect 33776 18507 33810 18541
rect 33866 18507 33900 18541
rect 33956 18507 33990 18541
rect 34046 18507 34080 18541
rect 34136 18507 34170 18541
rect 34226 18507 34260 18541
rect 34316 18507 34350 18541
rect 34406 18507 34440 18541
rect 34496 18507 34530 18541
rect 34586 18507 34620 18541
rect 34676 18507 34710 18541
rect 34766 18507 34800 18541
rect 34867 18484 34901 18518
rect 35020 18484 35054 18518
rect 35116 18507 35150 18541
rect 35206 18507 35240 18541
rect 35296 18507 35330 18541
rect 35386 18507 35420 18541
rect 35476 18507 35510 18541
rect 35566 18507 35600 18541
rect 35656 18507 35690 18541
rect 35746 18507 35780 18541
rect 35836 18507 35870 18541
rect 35926 18507 35960 18541
rect 36016 18507 36050 18541
rect 36106 18507 36140 18541
rect 36207 18484 36241 18518
rect 36360 18484 36394 18518
rect 36456 18507 36490 18541
rect 36546 18507 36580 18541
rect 36636 18507 36670 18541
rect 36726 18507 36760 18541
rect 36816 18507 36850 18541
rect 36906 18507 36940 18541
rect 36996 18507 37030 18541
rect 37086 18507 37120 18541
rect 37176 18507 37210 18541
rect 37266 18507 37300 18541
rect 37356 18507 37390 18541
rect 37446 18507 37480 18541
rect 37547 18484 37581 18518
rect 37700 18484 37734 18518
rect 37796 18507 37830 18541
rect 37886 18507 37920 18541
rect 37976 18507 38010 18541
rect 38066 18507 38100 18541
rect 38156 18507 38190 18541
rect 38246 18507 38280 18541
rect 38336 18507 38370 18541
rect 38426 18507 38460 18541
rect 38516 18507 38550 18541
rect 38606 18507 38640 18541
rect 38696 18507 38730 18541
rect 38786 18507 38820 18541
rect 38887 18484 38921 18518
rect 28320 18394 28354 18428
rect 28320 18304 28354 18338
rect 28320 18214 28354 18248
rect 28320 18124 28354 18158
rect 28320 18034 28354 18068
rect 28320 17944 28354 17978
rect 28320 17854 28354 17888
rect 28320 17764 28354 17798
rect 28320 17674 28354 17708
rect 28320 17584 28354 17618
rect 28320 17494 28354 17528
rect 29507 18394 29541 18428
rect 29660 18394 29694 18428
rect 29507 18304 29541 18338
rect 29660 18304 29694 18338
rect 29507 18214 29541 18248
rect 29660 18214 29694 18248
rect 29507 18124 29541 18158
rect 29660 18124 29694 18158
rect 29507 18034 29541 18068
rect 29660 18034 29694 18068
rect 29507 17944 29541 17978
rect 29660 17944 29694 17978
rect 29507 17854 29541 17888
rect 29660 17854 29694 17888
rect 29507 17764 29541 17798
rect 29660 17764 29694 17798
rect 29507 17674 29541 17708
rect 29660 17674 29694 17708
rect 29507 17584 29541 17618
rect 29660 17584 29694 17618
rect 29507 17494 29541 17528
rect 29660 17494 29694 17528
rect 28320 17404 28354 17438
rect 30847 18394 30881 18428
rect 31000 18394 31034 18428
rect 30847 18304 30881 18338
rect 31000 18304 31034 18338
rect 30847 18214 30881 18248
rect 31000 18214 31034 18248
rect 30847 18124 30881 18158
rect 31000 18124 31034 18158
rect 30847 18034 30881 18068
rect 31000 18034 31034 18068
rect 30847 17944 30881 17978
rect 31000 17944 31034 17978
rect 30847 17854 30881 17888
rect 31000 17854 31034 17888
rect 30847 17764 30881 17798
rect 31000 17764 31034 17798
rect 30847 17674 30881 17708
rect 31000 17674 31034 17708
rect 30847 17584 30881 17618
rect 31000 17584 31034 17618
rect 30847 17494 30881 17528
rect 31000 17494 31034 17528
rect 29507 17404 29541 17438
rect 29660 17404 29694 17438
rect 32187 18394 32221 18428
rect 32340 18394 32374 18428
rect 32187 18304 32221 18338
rect 32340 18304 32374 18338
rect 32187 18214 32221 18248
rect 32340 18214 32374 18248
rect 32187 18124 32221 18158
rect 32340 18124 32374 18158
rect 32187 18034 32221 18068
rect 32340 18034 32374 18068
rect 32187 17944 32221 17978
rect 32340 17944 32374 17978
rect 32187 17854 32221 17888
rect 32340 17854 32374 17888
rect 32187 17764 32221 17798
rect 32340 17764 32374 17798
rect 32187 17674 32221 17708
rect 32340 17674 32374 17708
rect 32187 17584 32221 17618
rect 32340 17584 32374 17618
rect 32187 17494 32221 17528
rect 32340 17494 32374 17528
rect 30847 17404 30881 17438
rect 31000 17404 31034 17438
rect 33527 18394 33561 18428
rect 33680 18394 33714 18428
rect 33527 18304 33561 18338
rect 33680 18304 33714 18338
rect 33527 18214 33561 18248
rect 33680 18214 33714 18248
rect 33527 18124 33561 18158
rect 33680 18124 33714 18158
rect 33527 18034 33561 18068
rect 33680 18034 33714 18068
rect 33527 17944 33561 17978
rect 33680 17944 33714 17978
rect 33527 17854 33561 17888
rect 33680 17854 33714 17888
rect 33527 17764 33561 17798
rect 33680 17764 33714 17798
rect 33527 17674 33561 17708
rect 33680 17674 33714 17708
rect 33527 17584 33561 17618
rect 33680 17584 33714 17618
rect 33527 17494 33561 17528
rect 33680 17494 33714 17528
rect 32187 17404 32221 17438
rect 32340 17404 32374 17438
rect 34867 18394 34901 18428
rect 35020 18394 35054 18428
rect 34867 18304 34901 18338
rect 35020 18304 35054 18338
rect 34867 18214 34901 18248
rect 35020 18214 35054 18248
rect 34867 18124 34901 18158
rect 35020 18124 35054 18158
rect 34867 18034 34901 18068
rect 35020 18034 35054 18068
rect 34867 17944 34901 17978
rect 35020 17944 35054 17978
rect 34867 17854 34901 17888
rect 35020 17854 35054 17888
rect 34867 17764 34901 17798
rect 35020 17764 35054 17798
rect 34867 17674 34901 17708
rect 35020 17674 35054 17708
rect 34867 17584 34901 17618
rect 35020 17584 35054 17618
rect 34867 17494 34901 17528
rect 35020 17494 35054 17528
rect 33527 17404 33561 17438
rect 33680 17404 33714 17438
rect 36207 18394 36241 18428
rect 36360 18394 36394 18428
rect 36207 18304 36241 18338
rect 36360 18304 36394 18338
rect 36207 18214 36241 18248
rect 36360 18214 36394 18248
rect 36207 18124 36241 18158
rect 36360 18124 36394 18158
rect 36207 18034 36241 18068
rect 36360 18034 36394 18068
rect 36207 17944 36241 17978
rect 36360 17944 36394 17978
rect 36207 17854 36241 17888
rect 36360 17854 36394 17888
rect 36207 17764 36241 17798
rect 36360 17764 36394 17798
rect 36207 17674 36241 17708
rect 36360 17674 36394 17708
rect 36207 17584 36241 17618
rect 36360 17584 36394 17618
rect 36207 17494 36241 17528
rect 36360 17494 36394 17528
rect 34867 17404 34901 17438
rect 35020 17404 35054 17438
rect 37547 18394 37581 18428
rect 37700 18394 37734 18428
rect 37547 18304 37581 18338
rect 37700 18304 37734 18338
rect 37547 18214 37581 18248
rect 37700 18214 37734 18248
rect 37547 18124 37581 18158
rect 37700 18124 37734 18158
rect 37547 18034 37581 18068
rect 37700 18034 37734 18068
rect 37547 17944 37581 17978
rect 37700 17944 37734 17978
rect 37547 17854 37581 17888
rect 37700 17854 37734 17888
rect 37547 17764 37581 17798
rect 37700 17764 37734 17798
rect 37547 17674 37581 17708
rect 37700 17674 37734 17708
rect 37547 17584 37581 17618
rect 37700 17584 37734 17618
rect 37547 17494 37581 17528
rect 37700 17494 37734 17528
rect 36207 17404 36241 17438
rect 36360 17404 36394 17438
rect 38887 18394 38921 18428
rect 38887 18304 38921 18338
rect 38887 18214 38921 18248
rect 38887 18124 38921 18158
rect 38887 18034 38921 18068
rect 38887 17944 38921 17978
rect 38887 17854 38921 17888
rect 38887 17764 38921 17798
rect 40255 17821 40697 17923
rect 38887 17674 38921 17708
rect 38887 17584 38921 17618
rect 38887 17494 38921 17528
rect 37547 17404 37581 17438
rect 37700 17404 37734 17438
rect 38887 17404 38921 17438
rect 28416 17320 28450 17354
rect 28506 17320 28540 17354
rect 28596 17320 28630 17354
rect 28686 17320 28720 17354
rect 28776 17320 28810 17354
rect 28866 17320 28900 17354
rect 28956 17320 28990 17354
rect 29046 17320 29080 17354
rect 29136 17320 29170 17354
rect 29226 17320 29260 17354
rect 29316 17320 29350 17354
rect 29406 17320 29440 17354
rect 29756 17320 29790 17354
rect 29846 17320 29880 17354
rect 29936 17320 29970 17354
rect 30026 17320 30060 17354
rect 30116 17320 30150 17354
rect 30206 17320 30240 17354
rect 30296 17320 30330 17354
rect 30386 17320 30420 17354
rect 30476 17320 30510 17354
rect 30566 17320 30600 17354
rect 30656 17320 30690 17354
rect 30746 17320 30780 17354
rect 31096 17320 31130 17354
rect 31186 17320 31220 17354
rect 31276 17320 31310 17354
rect 31366 17320 31400 17354
rect 31456 17320 31490 17354
rect 31546 17320 31580 17354
rect 31636 17320 31670 17354
rect 31726 17320 31760 17354
rect 31816 17320 31850 17354
rect 31906 17320 31940 17354
rect 31996 17320 32030 17354
rect 32086 17320 32120 17354
rect 32436 17320 32470 17354
rect 32526 17320 32560 17354
rect 32616 17320 32650 17354
rect 32706 17320 32740 17354
rect 32796 17320 32830 17354
rect 32886 17320 32920 17354
rect 32976 17320 33010 17354
rect 33066 17320 33100 17354
rect 33156 17320 33190 17354
rect 33246 17320 33280 17354
rect 33336 17320 33370 17354
rect 33426 17320 33460 17354
rect 33776 17320 33810 17354
rect 33866 17320 33900 17354
rect 33956 17320 33990 17354
rect 34046 17320 34080 17354
rect 34136 17320 34170 17354
rect 34226 17320 34260 17354
rect 34316 17320 34350 17354
rect 34406 17320 34440 17354
rect 34496 17320 34530 17354
rect 34586 17320 34620 17354
rect 34676 17320 34710 17354
rect 34766 17320 34800 17354
rect 35116 17320 35150 17354
rect 35206 17320 35240 17354
rect 35296 17320 35330 17354
rect 35386 17320 35420 17354
rect 35476 17320 35510 17354
rect 35566 17320 35600 17354
rect 35656 17320 35690 17354
rect 35746 17320 35780 17354
rect 35836 17320 35870 17354
rect 35926 17320 35960 17354
rect 36016 17320 36050 17354
rect 36106 17320 36140 17354
rect 36456 17320 36490 17354
rect 36546 17320 36580 17354
rect 36636 17320 36670 17354
rect 36726 17320 36760 17354
rect 36816 17320 36850 17354
rect 36906 17320 36940 17354
rect 36996 17320 37030 17354
rect 37086 17320 37120 17354
rect 37176 17320 37210 17354
rect 37266 17320 37300 17354
rect 37356 17320 37390 17354
rect 37446 17320 37480 17354
rect 37796 17320 37830 17354
rect 37886 17320 37920 17354
rect 37976 17320 38010 17354
rect 38066 17320 38100 17354
rect 38156 17320 38190 17354
rect 38246 17320 38280 17354
rect 38336 17320 38370 17354
rect 38426 17320 38460 17354
rect 38516 17320 38550 17354
rect 38606 17320 38640 17354
rect 38696 17320 38730 17354
rect 38786 17320 38820 17354
rect 28320 14724 28354 14758
rect 28416 14747 28450 14781
rect 28506 14747 28540 14781
rect 28596 14747 28630 14781
rect 28686 14747 28720 14781
rect 28776 14747 28810 14781
rect 28866 14747 28900 14781
rect 28956 14747 28990 14781
rect 29046 14747 29080 14781
rect 29136 14747 29170 14781
rect 29226 14747 29260 14781
rect 29316 14747 29350 14781
rect 29406 14747 29440 14781
rect 29507 14724 29541 14758
rect 29660 14724 29694 14758
rect 29756 14747 29790 14781
rect 29846 14747 29880 14781
rect 29936 14747 29970 14781
rect 30026 14747 30060 14781
rect 30116 14747 30150 14781
rect 30206 14747 30240 14781
rect 30296 14747 30330 14781
rect 30386 14747 30420 14781
rect 30476 14747 30510 14781
rect 30566 14747 30600 14781
rect 30656 14747 30690 14781
rect 30746 14747 30780 14781
rect 30847 14724 30881 14758
rect 31000 14724 31034 14758
rect 31096 14747 31130 14781
rect 31186 14747 31220 14781
rect 31276 14747 31310 14781
rect 31366 14747 31400 14781
rect 31456 14747 31490 14781
rect 31546 14747 31580 14781
rect 31636 14747 31670 14781
rect 31726 14747 31760 14781
rect 31816 14747 31850 14781
rect 31906 14747 31940 14781
rect 31996 14747 32030 14781
rect 32086 14747 32120 14781
rect 32187 14724 32221 14758
rect 32340 14724 32374 14758
rect 32436 14747 32470 14781
rect 32526 14747 32560 14781
rect 32616 14747 32650 14781
rect 32706 14747 32740 14781
rect 32796 14747 32830 14781
rect 32886 14747 32920 14781
rect 32976 14747 33010 14781
rect 33066 14747 33100 14781
rect 33156 14747 33190 14781
rect 33246 14747 33280 14781
rect 33336 14747 33370 14781
rect 33426 14747 33460 14781
rect 33527 14724 33561 14758
rect 33680 14724 33714 14758
rect 33776 14747 33810 14781
rect 33866 14747 33900 14781
rect 33956 14747 33990 14781
rect 34046 14747 34080 14781
rect 34136 14747 34170 14781
rect 34226 14747 34260 14781
rect 34316 14747 34350 14781
rect 34406 14747 34440 14781
rect 34496 14747 34530 14781
rect 34586 14747 34620 14781
rect 34676 14747 34710 14781
rect 34766 14747 34800 14781
rect 34867 14724 34901 14758
rect 35020 14724 35054 14758
rect 35116 14747 35150 14781
rect 35206 14747 35240 14781
rect 35296 14747 35330 14781
rect 35386 14747 35420 14781
rect 35476 14747 35510 14781
rect 35566 14747 35600 14781
rect 35656 14747 35690 14781
rect 35746 14747 35780 14781
rect 35836 14747 35870 14781
rect 35926 14747 35960 14781
rect 36016 14747 36050 14781
rect 36106 14747 36140 14781
rect 36207 14724 36241 14758
rect 36360 14724 36394 14758
rect 36456 14747 36490 14781
rect 36546 14747 36580 14781
rect 36636 14747 36670 14781
rect 36726 14747 36760 14781
rect 36816 14747 36850 14781
rect 36906 14747 36940 14781
rect 36996 14747 37030 14781
rect 37086 14747 37120 14781
rect 37176 14747 37210 14781
rect 37266 14747 37300 14781
rect 37356 14747 37390 14781
rect 37446 14747 37480 14781
rect 37547 14724 37581 14758
rect 37700 14724 37734 14758
rect 37796 14747 37830 14781
rect 37886 14747 37920 14781
rect 37976 14747 38010 14781
rect 38066 14747 38100 14781
rect 38156 14747 38190 14781
rect 38246 14747 38280 14781
rect 38336 14747 38370 14781
rect 38426 14747 38460 14781
rect 38516 14747 38550 14781
rect 38606 14747 38640 14781
rect 38696 14747 38730 14781
rect 38786 14747 38820 14781
rect 38887 14724 38921 14758
rect 28320 14634 28354 14668
rect 28320 14544 28354 14578
rect 28320 14454 28354 14488
rect 28320 14364 28354 14398
rect 28320 14274 28354 14308
rect 8895 14061 9337 14163
rect 11639 14061 12081 14163
rect 14383 14061 14825 14163
rect 24575 14061 25017 14163
rect 28320 14184 28354 14218
rect 28320 14094 28354 14128
rect 28320 14004 28354 14038
rect 28320 13914 28354 13948
rect 28320 13824 28354 13858
rect 28320 13734 28354 13768
rect 29507 14634 29541 14668
rect 29660 14634 29694 14668
rect 29507 14544 29541 14578
rect 29660 14544 29694 14578
rect 29507 14454 29541 14488
rect 29660 14454 29694 14488
rect 29507 14364 29541 14398
rect 29660 14364 29694 14398
rect 29507 14274 29541 14308
rect 29660 14274 29694 14308
rect 29507 14184 29541 14218
rect 29660 14184 29694 14218
rect 29507 14094 29541 14128
rect 29660 14094 29694 14128
rect 29507 14004 29541 14038
rect 29660 14004 29694 14038
rect 29507 13914 29541 13948
rect 29660 13914 29694 13948
rect 29507 13824 29541 13858
rect 29660 13824 29694 13858
rect 29507 13734 29541 13768
rect 29660 13734 29694 13768
rect 28320 13644 28354 13678
rect 30847 14634 30881 14668
rect 31000 14634 31034 14668
rect 30847 14544 30881 14578
rect 31000 14544 31034 14578
rect 30847 14454 30881 14488
rect 31000 14454 31034 14488
rect 30847 14364 30881 14398
rect 31000 14364 31034 14398
rect 30847 14274 30881 14308
rect 31000 14274 31034 14308
rect 30847 14184 30881 14218
rect 31000 14184 31034 14218
rect 30847 14094 30881 14128
rect 31000 14094 31034 14128
rect 30847 14004 30881 14038
rect 31000 14004 31034 14038
rect 30847 13914 30881 13948
rect 31000 13914 31034 13948
rect 30847 13824 30881 13858
rect 31000 13824 31034 13858
rect 30847 13734 30881 13768
rect 31000 13734 31034 13768
rect 29507 13644 29541 13678
rect 29660 13644 29694 13678
rect 32187 14634 32221 14668
rect 32340 14634 32374 14668
rect 32187 14544 32221 14578
rect 32340 14544 32374 14578
rect 32187 14454 32221 14488
rect 32340 14454 32374 14488
rect 32187 14364 32221 14398
rect 32340 14364 32374 14398
rect 32187 14274 32221 14308
rect 32340 14274 32374 14308
rect 32187 14184 32221 14218
rect 32340 14184 32374 14218
rect 32187 14094 32221 14128
rect 32340 14094 32374 14128
rect 32187 14004 32221 14038
rect 32340 14004 32374 14038
rect 32187 13914 32221 13948
rect 32340 13914 32374 13948
rect 32187 13824 32221 13858
rect 32340 13824 32374 13858
rect 32187 13734 32221 13768
rect 32340 13734 32374 13768
rect 30847 13644 30881 13678
rect 31000 13644 31034 13678
rect 33527 14634 33561 14668
rect 33680 14634 33714 14668
rect 33527 14544 33561 14578
rect 33680 14544 33714 14578
rect 33527 14454 33561 14488
rect 33680 14454 33714 14488
rect 33527 14364 33561 14398
rect 33680 14364 33714 14398
rect 33527 14274 33561 14308
rect 33680 14274 33714 14308
rect 33527 14184 33561 14218
rect 33680 14184 33714 14218
rect 33527 14094 33561 14128
rect 33680 14094 33714 14128
rect 33527 14004 33561 14038
rect 33680 14004 33714 14038
rect 33527 13914 33561 13948
rect 33680 13914 33714 13948
rect 33527 13824 33561 13858
rect 33680 13824 33714 13858
rect 33527 13734 33561 13768
rect 33680 13734 33714 13768
rect 32187 13644 32221 13678
rect 32340 13644 32374 13678
rect 34867 14634 34901 14668
rect 35020 14634 35054 14668
rect 34867 14544 34901 14578
rect 35020 14544 35054 14578
rect 34867 14454 34901 14488
rect 35020 14454 35054 14488
rect 34867 14364 34901 14398
rect 35020 14364 35054 14398
rect 34867 14274 34901 14308
rect 35020 14274 35054 14308
rect 34867 14184 34901 14218
rect 35020 14184 35054 14218
rect 34867 14094 34901 14128
rect 35020 14094 35054 14128
rect 34867 14004 34901 14038
rect 35020 14004 35054 14038
rect 34867 13914 34901 13948
rect 35020 13914 35054 13948
rect 34867 13824 34901 13858
rect 35020 13824 35054 13858
rect 34867 13734 34901 13768
rect 35020 13734 35054 13768
rect 33527 13644 33561 13678
rect 33680 13644 33714 13678
rect 36207 14634 36241 14668
rect 36360 14634 36394 14668
rect 36207 14544 36241 14578
rect 36360 14544 36394 14578
rect 36207 14454 36241 14488
rect 36360 14454 36394 14488
rect 36207 14364 36241 14398
rect 36360 14364 36394 14398
rect 36207 14274 36241 14308
rect 36360 14274 36394 14308
rect 36207 14184 36241 14218
rect 36360 14184 36394 14218
rect 36207 14094 36241 14128
rect 36360 14094 36394 14128
rect 36207 14004 36241 14038
rect 36360 14004 36394 14038
rect 36207 13914 36241 13948
rect 36360 13914 36394 13948
rect 36207 13824 36241 13858
rect 36360 13824 36394 13858
rect 36207 13734 36241 13768
rect 36360 13734 36394 13768
rect 34867 13644 34901 13678
rect 35020 13644 35054 13678
rect 37547 14634 37581 14668
rect 37700 14634 37734 14668
rect 37547 14544 37581 14578
rect 37700 14544 37734 14578
rect 37547 14454 37581 14488
rect 37700 14454 37734 14488
rect 37547 14364 37581 14398
rect 37700 14364 37734 14398
rect 37547 14274 37581 14308
rect 37700 14274 37734 14308
rect 37547 14184 37581 14218
rect 37700 14184 37734 14218
rect 37547 14094 37581 14128
rect 37700 14094 37734 14128
rect 37547 14004 37581 14038
rect 37700 14004 37734 14038
rect 37547 13914 37581 13948
rect 37700 13914 37734 13948
rect 37547 13824 37581 13858
rect 37700 13824 37734 13858
rect 37547 13734 37581 13768
rect 37700 13734 37734 13768
rect 36207 13644 36241 13678
rect 36360 13644 36394 13678
rect 38887 14634 38921 14668
rect 38887 14544 38921 14578
rect 38887 14454 38921 14488
rect 38887 14364 38921 14398
rect 38887 14274 38921 14308
rect 38887 14184 38921 14218
rect 38887 14094 38921 14128
rect 38887 14004 38921 14038
rect 40255 14061 40697 14163
rect 38887 13914 38921 13948
rect 38887 13824 38921 13858
rect 38887 13734 38921 13768
rect 37547 13644 37581 13678
rect 37700 13644 37734 13678
rect 38887 13644 38921 13678
rect 28416 13560 28450 13594
rect 28506 13560 28540 13594
rect 28596 13560 28630 13594
rect 28686 13560 28720 13594
rect 28776 13560 28810 13594
rect 28866 13560 28900 13594
rect 28956 13560 28990 13594
rect 29046 13560 29080 13594
rect 29136 13560 29170 13594
rect 29226 13560 29260 13594
rect 29316 13560 29350 13594
rect 29406 13560 29440 13594
rect 29756 13560 29790 13594
rect 29846 13560 29880 13594
rect 29936 13560 29970 13594
rect 30026 13560 30060 13594
rect 30116 13560 30150 13594
rect 30206 13560 30240 13594
rect 30296 13560 30330 13594
rect 30386 13560 30420 13594
rect 30476 13560 30510 13594
rect 30566 13560 30600 13594
rect 30656 13560 30690 13594
rect 30746 13560 30780 13594
rect 31096 13560 31130 13594
rect 31186 13560 31220 13594
rect 31276 13560 31310 13594
rect 31366 13560 31400 13594
rect 31456 13560 31490 13594
rect 31546 13560 31580 13594
rect 31636 13560 31670 13594
rect 31726 13560 31760 13594
rect 31816 13560 31850 13594
rect 31906 13560 31940 13594
rect 31996 13560 32030 13594
rect 32086 13560 32120 13594
rect 32436 13560 32470 13594
rect 32526 13560 32560 13594
rect 32616 13560 32650 13594
rect 32706 13560 32740 13594
rect 32796 13560 32830 13594
rect 32886 13560 32920 13594
rect 32976 13560 33010 13594
rect 33066 13560 33100 13594
rect 33156 13560 33190 13594
rect 33246 13560 33280 13594
rect 33336 13560 33370 13594
rect 33426 13560 33460 13594
rect 33776 13560 33810 13594
rect 33866 13560 33900 13594
rect 33956 13560 33990 13594
rect 34046 13560 34080 13594
rect 34136 13560 34170 13594
rect 34226 13560 34260 13594
rect 34316 13560 34350 13594
rect 34406 13560 34440 13594
rect 34496 13560 34530 13594
rect 34586 13560 34620 13594
rect 34676 13560 34710 13594
rect 34766 13560 34800 13594
rect 35116 13560 35150 13594
rect 35206 13560 35240 13594
rect 35296 13560 35330 13594
rect 35386 13560 35420 13594
rect 35476 13560 35510 13594
rect 35566 13560 35600 13594
rect 35656 13560 35690 13594
rect 35746 13560 35780 13594
rect 35836 13560 35870 13594
rect 35926 13560 35960 13594
rect 36016 13560 36050 13594
rect 36106 13560 36140 13594
rect 36456 13560 36490 13594
rect 36546 13560 36580 13594
rect 36636 13560 36670 13594
rect 36726 13560 36760 13594
rect 36816 13560 36850 13594
rect 36906 13560 36940 13594
rect 36996 13560 37030 13594
rect 37086 13560 37120 13594
rect 37176 13560 37210 13594
rect 37266 13560 37300 13594
rect 37356 13560 37390 13594
rect 37446 13560 37480 13594
rect 37796 13560 37830 13594
rect 37886 13560 37920 13594
rect 37976 13560 38010 13594
rect 38066 13560 38100 13594
rect 38156 13560 38190 13594
rect 38246 13560 38280 13594
rect 38336 13560 38370 13594
rect 38426 13560 38460 13594
rect 38516 13560 38550 13594
rect 38606 13560 38640 13594
rect 38696 13560 38730 13594
rect 38786 13560 38820 13594
rect 8895 10301 9337 10403
rect 11639 10301 12081 10403
rect 14383 10301 14825 10403
rect 24863 10301 25305 10403
rect 27907 10301 28349 10403
rect 30651 10301 31093 10403
rect 33395 10301 33837 10403
rect 36139 10301 36581 10403
rect 38883 10301 39325 10403
rect 8895 6541 9337 6643
rect 15553 6541 15995 6643
rect 18597 6541 19039 6643
rect 21341 6541 21783 6643
rect 24085 6541 24527 6643
rect 26829 6541 27271 6643
rect 29573 6541 30015 6643
rect 32317 6541 32759 6643
rect 36139 6541 36581 6643
rect 38883 6541 39325 6643
<< nsubdiffcont >>
rect 16073 41325 16107 41359
rect 17373 41325 17407 41359
rect 18673 41325 18707 41359
rect 19973 41325 20007 41359
rect 21273 41325 21307 41359
rect 22573 41325 22607 41359
rect 23873 41325 23907 41359
rect 25173 41325 25207 41359
rect 26473 41325 26507 41359
rect 27773 41325 27807 41359
rect 29073 41325 29107 41359
rect 30373 41325 30407 41359
rect 31673 41325 31707 41359
rect 32973 41325 33007 41359
rect 34273 41325 34307 41359
rect 35573 41325 35607 41359
rect 36873 41325 36907 41359
rect 38173 41325 38207 41359
rect 39473 41325 39507 41359
rect 40773 41325 40807 41359
rect 14973 41275 15007 41309
rect 30344 37160 30378 37194
rect 30434 37160 30468 37194
rect 30524 37160 30558 37194
rect 30614 37160 30648 37194
rect 30704 37160 30738 37194
rect 30794 37160 30828 37194
rect 30884 37160 30918 37194
rect 30974 37160 31008 37194
rect 31064 37160 31098 37194
rect 30232 37103 30266 37137
rect 31122 37084 31156 37118
rect 30232 37013 30266 37047
rect 30232 36923 30266 36957
rect 30232 36833 30266 36867
rect 30232 36743 30266 36777
rect 30232 36653 30266 36687
rect 30232 36563 30266 36597
rect 30232 36473 30266 36507
rect 30232 36383 30266 36417
rect 31122 36994 31156 37028
rect 31122 36904 31156 36938
rect 31122 36814 31156 36848
rect 31122 36724 31156 36758
rect 31122 36634 31156 36668
rect 31122 36544 31156 36578
rect 31122 36454 31156 36488
rect 31122 36364 31156 36398
rect 30310 36270 30344 36304
rect 30400 36270 30434 36304
rect 30490 36270 30524 36304
rect 30580 36270 30614 36304
rect 30670 36270 30704 36304
rect 30760 36270 30794 36304
rect 30850 36270 30884 36304
rect 30940 36270 30974 36304
rect 31030 36270 31064 36304
rect 31684 37160 31718 37194
rect 31774 37160 31808 37194
rect 31864 37160 31898 37194
rect 31954 37160 31988 37194
rect 32044 37160 32078 37194
rect 32134 37160 32168 37194
rect 32224 37160 32258 37194
rect 32314 37160 32348 37194
rect 32404 37160 32438 37194
rect 31572 37103 31606 37137
rect 32462 37084 32496 37118
rect 31572 37013 31606 37047
rect 31572 36923 31606 36957
rect 31572 36833 31606 36867
rect 31572 36743 31606 36777
rect 31572 36653 31606 36687
rect 31572 36563 31606 36597
rect 31572 36473 31606 36507
rect 31572 36383 31606 36417
rect 32462 36994 32496 37028
rect 32462 36904 32496 36938
rect 32462 36814 32496 36848
rect 32462 36724 32496 36758
rect 32462 36634 32496 36668
rect 32462 36544 32496 36578
rect 32462 36454 32496 36488
rect 32462 36364 32496 36398
rect 31650 36270 31684 36304
rect 31740 36270 31774 36304
rect 31830 36270 31864 36304
rect 31920 36270 31954 36304
rect 32010 36270 32044 36304
rect 32100 36270 32134 36304
rect 32190 36270 32224 36304
rect 32280 36270 32314 36304
rect 32370 36270 32404 36304
rect 33024 37160 33058 37194
rect 33114 37160 33148 37194
rect 33204 37160 33238 37194
rect 33294 37160 33328 37194
rect 33384 37160 33418 37194
rect 33474 37160 33508 37194
rect 33564 37160 33598 37194
rect 33654 37160 33688 37194
rect 33744 37160 33778 37194
rect 32912 37103 32946 37137
rect 33802 37084 33836 37118
rect 32912 37013 32946 37047
rect 32912 36923 32946 36957
rect 32912 36833 32946 36867
rect 32912 36743 32946 36777
rect 32912 36653 32946 36687
rect 32912 36563 32946 36597
rect 32912 36473 32946 36507
rect 32912 36383 32946 36417
rect 33802 36994 33836 37028
rect 33802 36904 33836 36938
rect 33802 36814 33836 36848
rect 33802 36724 33836 36758
rect 33802 36634 33836 36668
rect 33802 36544 33836 36578
rect 33802 36454 33836 36488
rect 33802 36364 33836 36398
rect 32990 36270 33024 36304
rect 33080 36270 33114 36304
rect 33170 36270 33204 36304
rect 33260 36270 33294 36304
rect 33350 36270 33384 36304
rect 33440 36270 33474 36304
rect 33530 36270 33564 36304
rect 33620 36270 33654 36304
rect 33710 36270 33744 36304
rect 34364 37160 34398 37194
rect 34454 37160 34488 37194
rect 34544 37160 34578 37194
rect 34634 37160 34668 37194
rect 34724 37160 34758 37194
rect 34814 37160 34848 37194
rect 34904 37160 34938 37194
rect 34994 37160 35028 37194
rect 35084 37160 35118 37194
rect 34252 37103 34286 37137
rect 35142 37084 35176 37118
rect 34252 37013 34286 37047
rect 34252 36923 34286 36957
rect 34252 36833 34286 36867
rect 34252 36743 34286 36777
rect 34252 36653 34286 36687
rect 34252 36563 34286 36597
rect 34252 36473 34286 36507
rect 34252 36383 34286 36417
rect 35142 36994 35176 37028
rect 35142 36904 35176 36938
rect 35142 36814 35176 36848
rect 35142 36724 35176 36758
rect 35142 36634 35176 36668
rect 35142 36544 35176 36578
rect 35142 36454 35176 36488
rect 35142 36364 35176 36398
rect 34330 36270 34364 36304
rect 34420 36270 34454 36304
rect 34510 36270 34544 36304
rect 34600 36270 34634 36304
rect 34690 36270 34724 36304
rect 34780 36270 34814 36304
rect 34870 36270 34904 36304
rect 34960 36270 34994 36304
rect 35050 36270 35084 36304
rect 35704 37160 35738 37194
rect 35794 37160 35828 37194
rect 35884 37160 35918 37194
rect 35974 37160 36008 37194
rect 36064 37160 36098 37194
rect 36154 37160 36188 37194
rect 36244 37160 36278 37194
rect 36334 37160 36368 37194
rect 36424 37160 36458 37194
rect 35592 37103 35626 37137
rect 36482 37084 36516 37118
rect 35592 37013 35626 37047
rect 35592 36923 35626 36957
rect 35592 36833 35626 36867
rect 35592 36743 35626 36777
rect 35592 36653 35626 36687
rect 35592 36563 35626 36597
rect 35592 36473 35626 36507
rect 35592 36383 35626 36417
rect 36482 36994 36516 37028
rect 36482 36904 36516 36938
rect 36482 36814 36516 36848
rect 36482 36724 36516 36758
rect 36482 36634 36516 36668
rect 36482 36544 36516 36578
rect 36482 36454 36516 36488
rect 36482 36364 36516 36398
rect 35670 36270 35704 36304
rect 35760 36270 35794 36304
rect 35850 36270 35884 36304
rect 35940 36270 35974 36304
rect 36030 36270 36064 36304
rect 36120 36270 36154 36304
rect 36210 36270 36244 36304
rect 36300 36270 36334 36304
rect 36390 36270 36424 36304
rect 37044 37160 37078 37194
rect 37134 37160 37168 37194
rect 37224 37160 37258 37194
rect 37314 37160 37348 37194
rect 37404 37160 37438 37194
rect 37494 37160 37528 37194
rect 37584 37160 37618 37194
rect 37674 37160 37708 37194
rect 37764 37160 37798 37194
rect 36932 37103 36966 37137
rect 37822 37084 37856 37118
rect 36932 37013 36966 37047
rect 36932 36923 36966 36957
rect 36932 36833 36966 36867
rect 36932 36743 36966 36777
rect 36932 36653 36966 36687
rect 36932 36563 36966 36597
rect 36932 36473 36966 36507
rect 36932 36383 36966 36417
rect 37822 36994 37856 37028
rect 37822 36904 37856 36938
rect 37822 36814 37856 36848
rect 37822 36724 37856 36758
rect 37822 36634 37856 36668
rect 37822 36544 37856 36578
rect 37822 36454 37856 36488
rect 37822 36364 37856 36398
rect 37010 36270 37044 36304
rect 37100 36270 37134 36304
rect 37190 36270 37224 36304
rect 37280 36270 37314 36304
rect 37370 36270 37404 36304
rect 37460 36270 37494 36304
rect 37550 36270 37584 36304
rect 37640 36270 37674 36304
rect 37730 36270 37764 36304
rect 38384 37160 38418 37194
rect 38474 37160 38508 37194
rect 38564 37160 38598 37194
rect 38654 37160 38688 37194
rect 38744 37160 38778 37194
rect 38834 37160 38868 37194
rect 38924 37160 38958 37194
rect 39014 37160 39048 37194
rect 39104 37160 39138 37194
rect 38272 37103 38306 37137
rect 39162 37084 39196 37118
rect 38272 37013 38306 37047
rect 38272 36923 38306 36957
rect 38272 36833 38306 36867
rect 38272 36743 38306 36777
rect 38272 36653 38306 36687
rect 38272 36563 38306 36597
rect 38272 36473 38306 36507
rect 38272 36383 38306 36417
rect 39162 36994 39196 37028
rect 39162 36904 39196 36938
rect 39162 36814 39196 36848
rect 39162 36724 39196 36758
rect 39162 36634 39196 36668
rect 39162 36544 39196 36578
rect 39162 36454 39196 36488
rect 39162 36364 39196 36398
rect 38350 36270 38384 36304
rect 38440 36270 38474 36304
rect 38530 36270 38564 36304
rect 38620 36270 38654 36304
rect 38710 36270 38744 36304
rect 38800 36270 38834 36304
rect 38890 36270 38924 36304
rect 38980 36270 39014 36304
rect 39070 36270 39104 36304
rect 15191 33805 15225 33839
rect 16491 33805 16525 33839
rect 17791 33805 17825 33839
rect 19091 33805 19125 33839
rect 20391 33805 20425 33839
rect 21691 33805 21725 33839
rect 22991 33805 23025 33839
rect 24291 33805 24325 33839
rect 25591 33805 25625 33839
rect 26891 33805 26925 33839
rect 28191 33805 28225 33839
rect 29491 33805 29525 33839
rect 30791 33805 30825 33839
rect 32091 33805 32125 33839
rect 33391 33805 33425 33839
rect 34691 33805 34725 33839
rect 35991 33805 36025 33839
rect 37291 33805 37325 33839
rect 38591 33805 38625 33839
rect 39891 33805 39925 33839
rect 14091 33755 14125 33789
rect 7057 30045 7091 30079
rect 8357 30045 8391 30079
rect 9657 30045 9691 30079
rect 10957 30045 10991 30079
rect 12257 30045 12291 30079
rect 13557 30045 13591 30079
rect 14857 30045 14891 30079
rect 16157 30045 16191 30079
rect 17457 30045 17491 30079
rect 18757 30045 18791 30079
rect 20057 30045 20091 30079
rect 21357 30045 21391 30079
rect 22657 30045 22691 30079
rect 23957 30045 23991 30079
rect 25257 30045 25291 30079
rect 26557 30045 26591 30079
rect 27857 30045 27891 30079
rect 29157 30045 29191 30079
rect 30457 30045 30491 30079
rect 31757 30045 31791 30079
rect 5957 29995 5991 30029
rect 35085 30045 35119 30079
rect 33985 29995 34019 30029
rect 10585 26285 10619 26319
rect 11885 26285 11919 26319
rect 13185 26285 13219 26319
rect 9485 26235 9519 26269
rect 28580 25880 28614 25914
rect 28670 25880 28704 25914
rect 28760 25880 28794 25914
rect 28850 25880 28884 25914
rect 28940 25880 28974 25914
rect 29030 25880 29064 25914
rect 29120 25880 29154 25914
rect 29210 25880 29244 25914
rect 29300 25880 29334 25914
rect 28468 25823 28502 25857
rect 29358 25804 29392 25838
rect 28468 25733 28502 25767
rect 28468 25643 28502 25677
rect 28468 25553 28502 25587
rect 28468 25463 28502 25497
rect 28468 25373 28502 25407
rect 28468 25283 28502 25317
rect 28468 25193 28502 25227
rect 28468 25103 28502 25137
rect 29358 25714 29392 25748
rect 29358 25624 29392 25658
rect 29358 25534 29392 25568
rect 29358 25444 29392 25478
rect 29358 25354 29392 25388
rect 29358 25264 29392 25298
rect 29358 25174 29392 25208
rect 29358 25084 29392 25118
rect 28546 24990 28580 25024
rect 28636 24990 28670 25024
rect 28726 24990 28760 25024
rect 28816 24990 28850 25024
rect 28906 24990 28940 25024
rect 28996 24990 29030 25024
rect 29086 24990 29120 25024
rect 29176 24990 29210 25024
rect 29266 24990 29300 25024
rect 29920 25880 29954 25914
rect 30010 25880 30044 25914
rect 30100 25880 30134 25914
rect 30190 25880 30224 25914
rect 30280 25880 30314 25914
rect 30370 25880 30404 25914
rect 30460 25880 30494 25914
rect 30550 25880 30584 25914
rect 30640 25880 30674 25914
rect 29808 25823 29842 25857
rect 30698 25804 30732 25838
rect 29808 25733 29842 25767
rect 29808 25643 29842 25677
rect 29808 25553 29842 25587
rect 29808 25463 29842 25497
rect 29808 25373 29842 25407
rect 29808 25283 29842 25317
rect 29808 25193 29842 25227
rect 29808 25103 29842 25137
rect 30698 25714 30732 25748
rect 30698 25624 30732 25658
rect 30698 25534 30732 25568
rect 30698 25444 30732 25478
rect 30698 25354 30732 25388
rect 30698 25264 30732 25298
rect 30698 25174 30732 25208
rect 30698 25084 30732 25118
rect 29886 24990 29920 25024
rect 29976 24990 30010 25024
rect 30066 24990 30100 25024
rect 30156 24990 30190 25024
rect 30246 24990 30280 25024
rect 30336 24990 30370 25024
rect 30426 24990 30460 25024
rect 30516 24990 30550 25024
rect 30606 24990 30640 25024
rect 31260 25880 31294 25914
rect 31350 25880 31384 25914
rect 31440 25880 31474 25914
rect 31530 25880 31564 25914
rect 31620 25880 31654 25914
rect 31710 25880 31744 25914
rect 31800 25880 31834 25914
rect 31890 25880 31924 25914
rect 31980 25880 32014 25914
rect 31148 25823 31182 25857
rect 32038 25804 32072 25838
rect 31148 25733 31182 25767
rect 31148 25643 31182 25677
rect 31148 25553 31182 25587
rect 31148 25463 31182 25497
rect 31148 25373 31182 25407
rect 31148 25283 31182 25317
rect 31148 25193 31182 25227
rect 31148 25103 31182 25137
rect 32038 25714 32072 25748
rect 32038 25624 32072 25658
rect 32038 25534 32072 25568
rect 32038 25444 32072 25478
rect 32038 25354 32072 25388
rect 32038 25264 32072 25298
rect 32038 25174 32072 25208
rect 32038 25084 32072 25118
rect 31226 24990 31260 25024
rect 31316 24990 31350 25024
rect 31406 24990 31440 25024
rect 31496 24990 31530 25024
rect 31586 24990 31620 25024
rect 31676 24990 31710 25024
rect 31766 24990 31800 25024
rect 31856 24990 31890 25024
rect 31946 24990 31980 25024
rect 32600 25880 32634 25914
rect 32690 25880 32724 25914
rect 32780 25880 32814 25914
rect 32870 25880 32904 25914
rect 32960 25880 32994 25914
rect 33050 25880 33084 25914
rect 33140 25880 33174 25914
rect 33230 25880 33264 25914
rect 33320 25880 33354 25914
rect 32488 25823 32522 25857
rect 33378 25804 33412 25838
rect 32488 25733 32522 25767
rect 32488 25643 32522 25677
rect 32488 25553 32522 25587
rect 32488 25463 32522 25497
rect 32488 25373 32522 25407
rect 32488 25283 32522 25317
rect 32488 25193 32522 25227
rect 32488 25103 32522 25137
rect 33378 25714 33412 25748
rect 33378 25624 33412 25658
rect 33378 25534 33412 25568
rect 33378 25444 33412 25478
rect 33378 25354 33412 25388
rect 33378 25264 33412 25298
rect 33378 25174 33412 25208
rect 33378 25084 33412 25118
rect 32566 24990 32600 25024
rect 32656 24990 32690 25024
rect 32746 24990 32780 25024
rect 32836 24990 32870 25024
rect 32926 24990 32960 25024
rect 33016 24990 33050 25024
rect 33106 24990 33140 25024
rect 33196 24990 33230 25024
rect 33286 24990 33320 25024
rect 33940 25880 33974 25914
rect 34030 25880 34064 25914
rect 34120 25880 34154 25914
rect 34210 25880 34244 25914
rect 34300 25880 34334 25914
rect 34390 25880 34424 25914
rect 34480 25880 34514 25914
rect 34570 25880 34604 25914
rect 34660 25880 34694 25914
rect 33828 25823 33862 25857
rect 34718 25804 34752 25838
rect 33828 25733 33862 25767
rect 33828 25643 33862 25677
rect 33828 25553 33862 25587
rect 33828 25463 33862 25497
rect 33828 25373 33862 25407
rect 33828 25283 33862 25317
rect 33828 25193 33862 25227
rect 33828 25103 33862 25137
rect 34718 25714 34752 25748
rect 34718 25624 34752 25658
rect 34718 25534 34752 25568
rect 34718 25444 34752 25478
rect 34718 25354 34752 25388
rect 34718 25264 34752 25298
rect 34718 25174 34752 25208
rect 34718 25084 34752 25118
rect 33906 24990 33940 25024
rect 33996 24990 34030 25024
rect 34086 24990 34120 25024
rect 34176 24990 34210 25024
rect 34266 24990 34300 25024
rect 34356 24990 34390 25024
rect 34446 24990 34480 25024
rect 34536 24990 34570 25024
rect 34626 24990 34660 25024
rect 35280 25880 35314 25914
rect 35370 25880 35404 25914
rect 35460 25880 35494 25914
rect 35550 25880 35584 25914
rect 35640 25880 35674 25914
rect 35730 25880 35764 25914
rect 35820 25880 35854 25914
rect 35910 25880 35944 25914
rect 36000 25880 36034 25914
rect 35168 25823 35202 25857
rect 36058 25804 36092 25838
rect 35168 25733 35202 25767
rect 35168 25643 35202 25677
rect 35168 25553 35202 25587
rect 35168 25463 35202 25497
rect 35168 25373 35202 25407
rect 35168 25283 35202 25317
rect 35168 25193 35202 25227
rect 35168 25103 35202 25137
rect 36058 25714 36092 25748
rect 36058 25624 36092 25658
rect 36058 25534 36092 25568
rect 36058 25444 36092 25478
rect 36058 25354 36092 25388
rect 36058 25264 36092 25298
rect 36058 25174 36092 25208
rect 36058 25084 36092 25118
rect 35246 24990 35280 25024
rect 35336 24990 35370 25024
rect 35426 24990 35460 25024
rect 35516 24990 35550 25024
rect 35606 24990 35640 25024
rect 35696 24990 35730 25024
rect 35786 24990 35820 25024
rect 35876 24990 35910 25024
rect 35966 24990 36000 25024
rect 36620 25880 36654 25914
rect 36710 25880 36744 25914
rect 36800 25880 36834 25914
rect 36890 25880 36924 25914
rect 36980 25880 37014 25914
rect 37070 25880 37104 25914
rect 37160 25880 37194 25914
rect 37250 25880 37284 25914
rect 37340 25880 37374 25914
rect 36508 25823 36542 25857
rect 37398 25804 37432 25838
rect 36508 25733 36542 25767
rect 36508 25643 36542 25677
rect 36508 25553 36542 25587
rect 36508 25463 36542 25497
rect 36508 25373 36542 25407
rect 36508 25283 36542 25317
rect 36508 25193 36542 25227
rect 36508 25103 36542 25137
rect 37398 25714 37432 25748
rect 37398 25624 37432 25658
rect 37398 25534 37432 25568
rect 37398 25444 37432 25478
rect 37398 25354 37432 25388
rect 37398 25264 37432 25298
rect 37398 25174 37432 25208
rect 37398 25084 37432 25118
rect 36586 24990 36620 25024
rect 36676 24990 36710 25024
rect 36766 24990 36800 25024
rect 36856 24990 36890 25024
rect 36946 24990 36980 25024
rect 37036 24990 37070 25024
rect 37126 24990 37160 25024
rect 37216 24990 37250 25024
rect 37306 24990 37340 25024
rect 37960 25880 37994 25914
rect 38050 25880 38084 25914
rect 38140 25880 38174 25914
rect 38230 25880 38264 25914
rect 38320 25880 38354 25914
rect 38410 25880 38444 25914
rect 38500 25880 38534 25914
rect 38590 25880 38624 25914
rect 38680 25880 38714 25914
rect 37848 25823 37882 25857
rect 38738 25804 38772 25838
rect 37848 25733 37882 25767
rect 37848 25643 37882 25677
rect 37848 25553 37882 25587
rect 37848 25463 37882 25497
rect 37848 25373 37882 25407
rect 37848 25283 37882 25317
rect 37848 25193 37882 25227
rect 37848 25103 37882 25137
rect 38738 25714 38772 25748
rect 38738 25624 38772 25658
rect 38738 25534 38772 25568
rect 38738 25444 38772 25478
rect 38738 25354 38772 25388
rect 38738 25264 38772 25298
rect 38738 25174 38772 25208
rect 38738 25084 38772 25118
rect 37926 24990 37960 25024
rect 38016 24990 38050 25024
rect 38106 24990 38140 25024
rect 38196 24990 38230 25024
rect 38286 24990 38320 25024
rect 38376 24990 38410 25024
rect 38466 24990 38500 25024
rect 38556 24990 38590 25024
rect 38646 24990 38680 25024
rect 8723 22525 8757 22559
rect 10023 22525 10057 22559
rect 11323 22525 11357 22559
rect 7623 22475 7657 22509
rect 21328 22120 21362 22154
rect 21418 22120 21452 22154
rect 21508 22120 21542 22154
rect 21598 22120 21632 22154
rect 21688 22120 21722 22154
rect 21778 22120 21812 22154
rect 21868 22120 21902 22154
rect 21958 22120 21992 22154
rect 22048 22120 22082 22154
rect 21216 22063 21250 22097
rect 22106 22044 22140 22078
rect 21216 21973 21250 22007
rect 21216 21883 21250 21917
rect 21216 21793 21250 21827
rect 21216 21703 21250 21737
rect 21216 21613 21250 21647
rect 21216 21523 21250 21557
rect 21216 21433 21250 21467
rect 21216 21343 21250 21377
rect 22106 21954 22140 21988
rect 22106 21864 22140 21898
rect 22106 21774 22140 21808
rect 22106 21684 22140 21718
rect 22106 21594 22140 21628
rect 22106 21504 22140 21538
rect 22106 21414 22140 21448
rect 22106 21324 22140 21358
rect 21294 21230 21328 21264
rect 21384 21230 21418 21264
rect 21474 21230 21508 21264
rect 21564 21230 21598 21264
rect 21654 21230 21688 21264
rect 21744 21230 21778 21264
rect 21834 21230 21868 21264
rect 21924 21230 21958 21264
rect 22014 21230 22048 21264
rect 28580 22120 28614 22154
rect 28670 22120 28704 22154
rect 28760 22120 28794 22154
rect 28850 22120 28884 22154
rect 28940 22120 28974 22154
rect 29030 22120 29064 22154
rect 29120 22120 29154 22154
rect 29210 22120 29244 22154
rect 29300 22120 29334 22154
rect 28468 22063 28502 22097
rect 29358 22044 29392 22078
rect 28468 21973 28502 22007
rect 28468 21883 28502 21917
rect 28468 21793 28502 21827
rect 28468 21703 28502 21737
rect 28468 21613 28502 21647
rect 28468 21523 28502 21557
rect 28468 21433 28502 21467
rect 28468 21343 28502 21377
rect 29358 21954 29392 21988
rect 29358 21864 29392 21898
rect 29358 21774 29392 21808
rect 29358 21684 29392 21718
rect 29358 21594 29392 21628
rect 29358 21504 29392 21538
rect 29358 21414 29392 21448
rect 29358 21324 29392 21358
rect 28546 21230 28580 21264
rect 28636 21230 28670 21264
rect 28726 21230 28760 21264
rect 28816 21230 28850 21264
rect 28906 21230 28940 21264
rect 28996 21230 29030 21264
rect 29086 21230 29120 21264
rect 29176 21230 29210 21264
rect 29266 21230 29300 21264
rect 29920 22120 29954 22154
rect 30010 22120 30044 22154
rect 30100 22120 30134 22154
rect 30190 22120 30224 22154
rect 30280 22120 30314 22154
rect 30370 22120 30404 22154
rect 30460 22120 30494 22154
rect 30550 22120 30584 22154
rect 30640 22120 30674 22154
rect 29808 22063 29842 22097
rect 30698 22044 30732 22078
rect 29808 21973 29842 22007
rect 29808 21883 29842 21917
rect 29808 21793 29842 21827
rect 29808 21703 29842 21737
rect 29808 21613 29842 21647
rect 29808 21523 29842 21557
rect 29808 21433 29842 21467
rect 29808 21343 29842 21377
rect 30698 21954 30732 21988
rect 30698 21864 30732 21898
rect 30698 21774 30732 21808
rect 30698 21684 30732 21718
rect 30698 21594 30732 21628
rect 30698 21504 30732 21538
rect 30698 21414 30732 21448
rect 30698 21324 30732 21358
rect 29886 21230 29920 21264
rect 29976 21230 30010 21264
rect 30066 21230 30100 21264
rect 30156 21230 30190 21264
rect 30246 21230 30280 21264
rect 30336 21230 30370 21264
rect 30426 21230 30460 21264
rect 30516 21230 30550 21264
rect 30606 21230 30640 21264
rect 31260 22120 31294 22154
rect 31350 22120 31384 22154
rect 31440 22120 31474 22154
rect 31530 22120 31564 22154
rect 31620 22120 31654 22154
rect 31710 22120 31744 22154
rect 31800 22120 31834 22154
rect 31890 22120 31924 22154
rect 31980 22120 32014 22154
rect 31148 22063 31182 22097
rect 32038 22044 32072 22078
rect 31148 21973 31182 22007
rect 31148 21883 31182 21917
rect 31148 21793 31182 21827
rect 31148 21703 31182 21737
rect 31148 21613 31182 21647
rect 31148 21523 31182 21557
rect 31148 21433 31182 21467
rect 31148 21343 31182 21377
rect 32038 21954 32072 21988
rect 32038 21864 32072 21898
rect 32038 21774 32072 21808
rect 32038 21684 32072 21718
rect 32038 21594 32072 21628
rect 32038 21504 32072 21538
rect 32038 21414 32072 21448
rect 32038 21324 32072 21358
rect 31226 21230 31260 21264
rect 31316 21230 31350 21264
rect 31406 21230 31440 21264
rect 31496 21230 31530 21264
rect 31586 21230 31620 21264
rect 31676 21230 31710 21264
rect 31766 21230 31800 21264
rect 31856 21230 31890 21264
rect 31946 21230 31980 21264
rect 32600 22120 32634 22154
rect 32690 22120 32724 22154
rect 32780 22120 32814 22154
rect 32870 22120 32904 22154
rect 32960 22120 32994 22154
rect 33050 22120 33084 22154
rect 33140 22120 33174 22154
rect 33230 22120 33264 22154
rect 33320 22120 33354 22154
rect 32488 22063 32522 22097
rect 33378 22044 33412 22078
rect 32488 21973 32522 22007
rect 32488 21883 32522 21917
rect 32488 21793 32522 21827
rect 32488 21703 32522 21737
rect 32488 21613 32522 21647
rect 32488 21523 32522 21557
rect 32488 21433 32522 21467
rect 32488 21343 32522 21377
rect 33378 21954 33412 21988
rect 33378 21864 33412 21898
rect 33378 21774 33412 21808
rect 33378 21684 33412 21718
rect 33378 21594 33412 21628
rect 33378 21504 33412 21538
rect 33378 21414 33412 21448
rect 33378 21324 33412 21358
rect 32566 21230 32600 21264
rect 32656 21230 32690 21264
rect 32746 21230 32780 21264
rect 32836 21230 32870 21264
rect 32926 21230 32960 21264
rect 33016 21230 33050 21264
rect 33106 21230 33140 21264
rect 33196 21230 33230 21264
rect 33286 21230 33320 21264
rect 33940 22120 33974 22154
rect 34030 22120 34064 22154
rect 34120 22120 34154 22154
rect 34210 22120 34244 22154
rect 34300 22120 34334 22154
rect 34390 22120 34424 22154
rect 34480 22120 34514 22154
rect 34570 22120 34604 22154
rect 34660 22120 34694 22154
rect 33828 22063 33862 22097
rect 34718 22044 34752 22078
rect 33828 21973 33862 22007
rect 33828 21883 33862 21917
rect 33828 21793 33862 21827
rect 33828 21703 33862 21737
rect 33828 21613 33862 21647
rect 33828 21523 33862 21557
rect 33828 21433 33862 21467
rect 33828 21343 33862 21377
rect 34718 21954 34752 21988
rect 34718 21864 34752 21898
rect 34718 21774 34752 21808
rect 34718 21684 34752 21718
rect 34718 21594 34752 21628
rect 34718 21504 34752 21538
rect 34718 21414 34752 21448
rect 34718 21324 34752 21358
rect 33906 21230 33940 21264
rect 33996 21230 34030 21264
rect 34086 21230 34120 21264
rect 34176 21230 34210 21264
rect 34266 21230 34300 21264
rect 34356 21230 34390 21264
rect 34446 21230 34480 21264
rect 34536 21230 34570 21264
rect 34626 21230 34660 21264
rect 35280 22120 35314 22154
rect 35370 22120 35404 22154
rect 35460 22120 35494 22154
rect 35550 22120 35584 22154
rect 35640 22120 35674 22154
rect 35730 22120 35764 22154
rect 35820 22120 35854 22154
rect 35910 22120 35944 22154
rect 36000 22120 36034 22154
rect 35168 22063 35202 22097
rect 36058 22044 36092 22078
rect 35168 21973 35202 22007
rect 35168 21883 35202 21917
rect 35168 21793 35202 21827
rect 35168 21703 35202 21737
rect 35168 21613 35202 21647
rect 35168 21523 35202 21557
rect 35168 21433 35202 21467
rect 35168 21343 35202 21377
rect 36058 21954 36092 21988
rect 36058 21864 36092 21898
rect 36058 21774 36092 21808
rect 36058 21684 36092 21718
rect 36058 21594 36092 21628
rect 36058 21504 36092 21538
rect 36058 21414 36092 21448
rect 36058 21324 36092 21358
rect 35246 21230 35280 21264
rect 35336 21230 35370 21264
rect 35426 21230 35460 21264
rect 35516 21230 35550 21264
rect 35606 21230 35640 21264
rect 35696 21230 35730 21264
rect 35786 21230 35820 21264
rect 35876 21230 35910 21264
rect 35966 21230 36000 21264
rect 36620 22120 36654 22154
rect 36710 22120 36744 22154
rect 36800 22120 36834 22154
rect 36890 22120 36924 22154
rect 36980 22120 37014 22154
rect 37070 22120 37104 22154
rect 37160 22120 37194 22154
rect 37250 22120 37284 22154
rect 37340 22120 37374 22154
rect 36508 22063 36542 22097
rect 37398 22044 37432 22078
rect 36508 21973 36542 22007
rect 36508 21883 36542 21917
rect 36508 21793 36542 21827
rect 36508 21703 36542 21737
rect 36508 21613 36542 21647
rect 36508 21523 36542 21557
rect 36508 21433 36542 21467
rect 36508 21343 36542 21377
rect 37398 21954 37432 21988
rect 37398 21864 37432 21898
rect 37398 21774 37432 21808
rect 37398 21684 37432 21718
rect 37398 21594 37432 21628
rect 37398 21504 37432 21538
rect 37398 21414 37432 21448
rect 37398 21324 37432 21358
rect 36586 21230 36620 21264
rect 36676 21230 36710 21264
rect 36766 21230 36800 21264
rect 36856 21230 36890 21264
rect 36946 21230 36980 21264
rect 37036 21230 37070 21264
rect 37126 21230 37160 21264
rect 37216 21230 37250 21264
rect 37306 21230 37340 21264
rect 37960 22120 37994 22154
rect 38050 22120 38084 22154
rect 38140 22120 38174 22154
rect 38230 22120 38264 22154
rect 38320 22120 38354 22154
rect 38410 22120 38444 22154
rect 38500 22120 38534 22154
rect 38590 22120 38624 22154
rect 38680 22120 38714 22154
rect 37848 22063 37882 22097
rect 38738 22044 38772 22078
rect 37848 21973 37882 22007
rect 37848 21883 37882 21917
rect 37848 21793 37882 21827
rect 37848 21703 37882 21737
rect 37848 21613 37882 21647
rect 37848 21523 37882 21557
rect 37848 21433 37882 21467
rect 37848 21343 37882 21377
rect 38738 21954 38772 21988
rect 38738 21864 38772 21898
rect 38738 21774 38772 21808
rect 38738 21684 38772 21718
rect 38738 21594 38772 21628
rect 38738 21504 38772 21538
rect 38738 21414 38772 21448
rect 38738 21324 38772 21358
rect 37926 21230 37960 21264
rect 38016 21230 38050 21264
rect 38106 21230 38140 21264
rect 38196 21230 38230 21264
rect 38286 21230 38320 21264
rect 38376 21230 38410 21264
rect 38466 21230 38500 21264
rect 38556 21230 38590 21264
rect 38646 21230 38680 21264
rect 24991 18765 25025 18799
rect 23891 18715 23925 18749
rect 28580 18360 28614 18394
rect 28670 18360 28704 18394
rect 28760 18360 28794 18394
rect 28850 18360 28884 18394
rect 28940 18360 28974 18394
rect 29030 18360 29064 18394
rect 29120 18360 29154 18394
rect 29210 18360 29244 18394
rect 29300 18360 29334 18394
rect 28468 18303 28502 18337
rect 29358 18284 29392 18318
rect 28468 18213 28502 18247
rect 28468 18123 28502 18157
rect 28468 18033 28502 18067
rect 28468 17943 28502 17977
rect 28468 17853 28502 17887
rect 28468 17763 28502 17797
rect 28468 17673 28502 17707
rect 28468 17583 28502 17617
rect 29358 18194 29392 18228
rect 29358 18104 29392 18138
rect 29358 18014 29392 18048
rect 29358 17924 29392 17958
rect 29358 17834 29392 17868
rect 29358 17744 29392 17778
rect 29358 17654 29392 17688
rect 29358 17564 29392 17598
rect 28546 17470 28580 17504
rect 28636 17470 28670 17504
rect 28726 17470 28760 17504
rect 28816 17470 28850 17504
rect 28906 17470 28940 17504
rect 28996 17470 29030 17504
rect 29086 17470 29120 17504
rect 29176 17470 29210 17504
rect 29266 17470 29300 17504
rect 29920 18360 29954 18394
rect 30010 18360 30044 18394
rect 30100 18360 30134 18394
rect 30190 18360 30224 18394
rect 30280 18360 30314 18394
rect 30370 18360 30404 18394
rect 30460 18360 30494 18394
rect 30550 18360 30584 18394
rect 30640 18360 30674 18394
rect 29808 18303 29842 18337
rect 30698 18284 30732 18318
rect 29808 18213 29842 18247
rect 29808 18123 29842 18157
rect 29808 18033 29842 18067
rect 29808 17943 29842 17977
rect 29808 17853 29842 17887
rect 29808 17763 29842 17797
rect 29808 17673 29842 17707
rect 29808 17583 29842 17617
rect 30698 18194 30732 18228
rect 30698 18104 30732 18138
rect 30698 18014 30732 18048
rect 30698 17924 30732 17958
rect 30698 17834 30732 17868
rect 30698 17744 30732 17778
rect 30698 17654 30732 17688
rect 30698 17564 30732 17598
rect 29886 17470 29920 17504
rect 29976 17470 30010 17504
rect 30066 17470 30100 17504
rect 30156 17470 30190 17504
rect 30246 17470 30280 17504
rect 30336 17470 30370 17504
rect 30426 17470 30460 17504
rect 30516 17470 30550 17504
rect 30606 17470 30640 17504
rect 31260 18360 31294 18394
rect 31350 18360 31384 18394
rect 31440 18360 31474 18394
rect 31530 18360 31564 18394
rect 31620 18360 31654 18394
rect 31710 18360 31744 18394
rect 31800 18360 31834 18394
rect 31890 18360 31924 18394
rect 31980 18360 32014 18394
rect 31148 18303 31182 18337
rect 32038 18284 32072 18318
rect 31148 18213 31182 18247
rect 31148 18123 31182 18157
rect 31148 18033 31182 18067
rect 31148 17943 31182 17977
rect 31148 17853 31182 17887
rect 31148 17763 31182 17797
rect 31148 17673 31182 17707
rect 31148 17583 31182 17617
rect 32038 18194 32072 18228
rect 32038 18104 32072 18138
rect 32038 18014 32072 18048
rect 32038 17924 32072 17958
rect 32038 17834 32072 17868
rect 32038 17744 32072 17778
rect 32038 17654 32072 17688
rect 32038 17564 32072 17598
rect 31226 17470 31260 17504
rect 31316 17470 31350 17504
rect 31406 17470 31440 17504
rect 31496 17470 31530 17504
rect 31586 17470 31620 17504
rect 31676 17470 31710 17504
rect 31766 17470 31800 17504
rect 31856 17470 31890 17504
rect 31946 17470 31980 17504
rect 32600 18360 32634 18394
rect 32690 18360 32724 18394
rect 32780 18360 32814 18394
rect 32870 18360 32904 18394
rect 32960 18360 32994 18394
rect 33050 18360 33084 18394
rect 33140 18360 33174 18394
rect 33230 18360 33264 18394
rect 33320 18360 33354 18394
rect 32488 18303 32522 18337
rect 33378 18284 33412 18318
rect 32488 18213 32522 18247
rect 32488 18123 32522 18157
rect 32488 18033 32522 18067
rect 32488 17943 32522 17977
rect 32488 17853 32522 17887
rect 32488 17763 32522 17797
rect 32488 17673 32522 17707
rect 32488 17583 32522 17617
rect 33378 18194 33412 18228
rect 33378 18104 33412 18138
rect 33378 18014 33412 18048
rect 33378 17924 33412 17958
rect 33378 17834 33412 17868
rect 33378 17744 33412 17778
rect 33378 17654 33412 17688
rect 33378 17564 33412 17598
rect 32566 17470 32600 17504
rect 32656 17470 32690 17504
rect 32746 17470 32780 17504
rect 32836 17470 32870 17504
rect 32926 17470 32960 17504
rect 33016 17470 33050 17504
rect 33106 17470 33140 17504
rect 33196 17470 33230 17504
rect 33286 17470 33320 17504
rect 33940 18360 33974 18394
rect 34030 18360 34064 18394
rect 34120 18360 34154 18394
rect 34210 18360 34244 18394
rect 34300 18360 34334 18394
rect 34390 18360 34424 18394
rect 34480 18360 34514 18394
rect 34570 18360 34604 18394
rect 34660 18360 34694 18394
rect 33828 18303 33862 18337
rect 34718 18284 34752 18318
rect 33828 18213 33862 18247
rect 33828 18123 33862 18157
rect 33828 18033 33862 18067
rect 33828 17943 33862 17977
rect 33828 17853 33862 17887
rect 33828 17763 33862 17797
rect 33828 17673 33862 17707
rect 33828 17583 33862 17617
rect 34718 18194 34752 18228
rect 34718 18104 34752 18138
rect 34718 18014 34752 18048
rect 34718 17924 34752 17958
rect 34718 17834 34752 17868
rect 34718 17744 34752 17778
rect 34718 17654 34752 17688
rect 34718 17564 34752 17598
rect 33906 17470 33940 17504
rect 33996 17470 34030 17504
rect 34086 17470 34120 17504
rect 34176 17470 34210 17504
rect 34266 17470 34300 17504
rect 34356 17470 34390 17504
rect 34446 17470 34480 17504
rect 34536 17470 34570 17504
rect 34626 17470 34660 17504
rect 35280 18360 35314 18394
rect 35370 18360 35404 18394
rect 35460 18360 35494 18394
rect 35550 18360 35584 18394
rect 35640 18360 35674 18394
rect 35730 18360 35764 18394
rect 35820 18360 35854 18394
rect 35910 18360 35944 18394
rect 36000 18360 36034 18394
rect 35168 18303 35202 18337
rect 36058 18284 36092 18318
rect 35168 18213 35202 18247
rect 35168 18123 35202 18157
rect 35168 18033 35202 18067
rect 35168 17943 35202 17977
rect 35168 17853 35202 17887
rect 35168 17763 35202 17797
rect 35168 17673 35202 17707
rect 35168 17583 35202 17617
rect 36058 18194 36092 18228
rect 36058 18104 36092 18138
rect 36058 18014 36092 18048
rect 36058 17924 36092 17958
rect 36058 17834 36092 17868
rect 36058 17744 36092 17778
rect 36058 17654 36092 17688
rect 36058 17564 36092 17598
rect 35246 17470 35280 17504
rect 35336 17470 35370 17504
rect 35426 17470 35460 17504
rect 35516 17470 35550 17504
rect 35606 17470 35640 17504
rect 35696 17470 35730 17504
rect 35786 17470 35820 17504
rect 35876 17470 35910 17504
rect 35966 17470 36000 17504
rect 36620 18360 36654 18394
rect 36710 18360 36744 18394
rect 36800 18360 36834 18394
rect 36890 18360 36924 18394
rect 36980 18360 37014 18394
rect 37070 18360 37104 18394
rect 37160 18360 37194 18394
rect 37250 18360 37284 18394
rect 37340 18360 37374 18394
rect 36508 18303 36542 18337
rect 37398 18284 37432 18318
rect 36508 18213 36542 18247
rect 36508 18123 36542 18157
rect 36508 18033 36542 18067
rect 36508 17943 36542 17977
rect 36508 17853 36542 17887
rect 36508 17763 36542 17797
rect 36508 17673 36542 17707
rect 36508 17583 36542 17617
rect 37398 18194 37432 18228
rect 37398 18104 37432 18138
rect 37398 18014 37432 18048
rect 37398 17924 37432 17958
rect 37398 17834 37432 17868
rect 37398 17744 37432 17778
rect 37398 17654 37432 17688
rect 37398 17564 37432 17598
rect 36586 17470 36620 17504
rect 36676 17470 36710 17504
rect 36766 17470 36800 17504
rect 36856 17470 36890 17504
rect 36946 17470 36980 17504
rect 37036 17470 37070 17504
rect 37126 17470 37160 17504
rect 37216 17470 37250 17504
rect 37306 17470 37340 17504
rect 37960 18360 37994 18394
rect 38050 18360 38084 18394
rect 38140 18360 38174 18394
rect 38230 18360 38264 18394
rect 38320 18360 38354 18394
rect 38410 18360 38444 18394
rect 38500 18360 38534 18394
rect 38590 18360 38624 18394
rect 38680 18360 38714 18394
rect 37848 18303 37882 18337
rect 38738 18284 38772 18318
rect 37848 18213 37882 18247
rect 37848 18123 37882 18157
rect 37848 18033 37882 18067
rect 37848 17943 37882 17977
rect 37848 17853 37882 17887
rect 37848 17763 37882 17797
rect 37848 17673 37882 17707
rect 37848 17583 37882 17617
rect 38738 18194 38772 18228
rect 38738 18104 38772 18138
rect 38738 18014 38772 18048
rect 38738 17924 38772 17958
rect 38738 17834 38772 17868
rect 38738 17744 38772 17778
rect 38738 17654 38772 17688
rect 38738 17564 38772 17598
rect 37926 17470 37960 17504
rect 38016 17470 38050 17504
rect 38106 17470 38140 17504
rect 38196 17470 38230 17504
rect 38286 17470 38320 17504
rect 38376 17470 38410 17504
rect 38466 17470 38500 17504
rect 38556 17470 38590 17504
rect 38646 17470 38680 17504
rect 28580 14600 28614 14634
rect 28670 14600 28704 14634
rect 28760 14600 28794 14634
rect 28850 14600 28884 14634
rect 28940 14600 28974 14634
rect 29030 14600 29064 14634
rect 29120 14600 29154 14634
rect 29210 14600 29244 14634
rect 29300 14600 29334 14634
rect 28468 14543 28502 14577
rect 29358 14524 29392 14558
rect 28468 14453 28502 14487
rect 28468 14363 28502 14397
rect 28468 14273 28502 14307
rect 28468 14183 28502 14217
rect 28468 14093 28502 14127
rect 28468 14003 28502 14037
rect 28468 13913 28502 13947
rect 28468 13823 28502 13857
rect 29358 14434 29392 14468
rect 29358 14344 29392 14378
rect 29358 14254 29392 14288
rect 29358 14164 29392 14198
rect 29358 14074 29392 14108
rect 29358 13984 29392 14018
rect 29358 13894 29392 13928
rect 29358 13804 29392 13838
rect 28546 13710 28580 13744
rect 28636 13710 28670 13744
rect 28726 13710 28760 13744
rect 28816 13710 28850 13744
rect 28906 13710 28940 13744
rect 28996 13710 29030 13744
rect 29086 13710 29120 13744
rect 29176 13710 29210 13744
rect 29266 13710 29300 13744
rect 29920 14600 29954 14634
rect 30010 14600 30044 14634
rect 30100 14600 30134 14634
rect 30190 14600 30224 14634
rect 30280 14600 30314 14634
rect 30370 14600 30404 14634
rect 30460 14600 30494 14634
rect 30550 14600 30584 14634
rect 30640 14600 30674 14634
rect 29808 14543 29842 14577
rect 30698 14524 30732 14558
rect 29808 14453 29842 14487
rect 29808 14363 29842 14397
rect 29808 14273 29842 14307
rect 29808 14183 29842 14217
rect 29808 14093 29842 14127
rect 29808 14003 29842 14037
rect 29808 13913 29842 13947
rect 29808 13823 29842 13857
rect 30698 14434 30732 14468
rect 30698 14344 30732 14378
rect 30698 14254 30732 14288
rect 30698 14164 30732 14198
rect 30698 14074 30732 14108
rect 30698 13984 30732 14018
rect 30698 13894 30732 13928
rect 30698 13804 30732 13838
rect 29886 13710 29920 13744
rect 29976 13710 30010 13744
rect 30066 13710 30100 13744
rect 30156 13710 30190 13744
rect 30246 13710 30280 13744
rect 30336 13710 30370 13744
rect 30426 13710 30460 13744
rect 30516 13710 30550 13744
rect 30606 13710 30640 13744
rect 31260 14600 31294 14634
rect 31350 14600 31384 14634
rect 31440 14600 31474 14634
rect 31530 14600 31564 14634
rect 31620 14600 31654 14634
rect 31710 14600 31744 14634
rect 31800 14600 31834 14634
rect 31890 14600 31924 14634
rect 31980 14600 32014 14634
rect 31148 14543 31182 14577
rect 32038 14524 32072 14558
rect 31148 14453 31182 14487
rect 31148 14363 31182 14397
rect 31148 14273 31182 14307
rect 31148 14183 31182 14217
rect 31148 14093 31182 14127
rect 31148 14003 31182 14037
rect 31148 13913 31182 13947
rect 31148 13823 31182 13857
rect 32038 14434 32072 14468
rect 32038 14344 32072 14378
rect 32038 14254 32072 14288
rect 32038 14164 32072 14198
rect 32038 14074 32072 14108
rect 32038 13984 32072 14018
rect 32038 13894 32072 13928
rect 32038 13804 32072 13838
rect 31226 13710 31260 13744
rect 31316 13710 31350 13744
rect 31406 13710 31440 13744
rect 31496 13710 31530 13744
rect 31586 13710 31620 13744
rect 31676 13710 31710 13744
rect 31766 13710 31800 13744
rect 31856 13710 31890 13744
rect 31946 13710 31980 13744
rect 32600 14600 32634 14634
rect 32690 14600 32724 14634
rect 32780 14600 32814 14634
rect 32870 14600 32904 14634
rect 32960 14600 32994 14634
rect 33050 14600 33084 14634
rect 33140 14600 33174 14634
rect 33230 14600 33264 14634
rect 33320 14600 33354 14634
rect 32488 14543 32522 14577
rect 33378 14524 33412 14558
rect 32488 14453 32522 14487
rect 32488 14363 32522 14397
rect 32488 14273 32522 14307
rect 32488 14183 32522 14217
rect 32488 14093 32522 14127
rect 32488 14003 32522 14037
rect 32488 13913 32522 13947
rect 32488 13823 32522 13857
rect 33378 14434 33412 14468
rect 33378 14344 33412 14378
rect 33378 14254 33412 14288
rect 33378 14164 33412 14198
rect 33378 14074 33412 14108
rect 33378 13984 33412 14018
rect 33378 13894 33412 13928
rect 33378 13804 33412 13838
rect 32566 13710 32600 13744
rect 32656 13710 32690 13744
rect 32746 13710 32780 13744
rect 32836 13710 32870 13744
rect 32926 13710 32960 13744
rect 33016 13710 33050 13744
rect 33106 13710 33140 13744
rect 33196 13710 33230 13744
rect 33286 13710 33320 13744
rect 33940 14600 33974 14634
rect 34030 14600 34064 14634
rect 34120 14600 34154 14634
rect 34210 14600 34244 14634
rect 34300 14600 34334 14634
rect 34390 14600 34424 14634
rect 34480 14600 34514 14634
rect 34570 14600 34604 14634
rect 34660 14600 34694 14634
rect 33828 14543 33862 14577
rect 34718 14524 34752 14558
rect 33828 14453 33862 14487
rect 33828 14363 33862 14397
rect 33828 14273 33862 14307
rect 33828 14183 33862 14217
rect 33828 14093 33862 14127
rect 33828 14003 33862 14037
rect 33828 13913 33862 13947
rect 33828 13823 33862 13857
rect 34718 14434 34752 14468
rect 34718 14344 34752 14378
rect 34718 14254 34752 14288
rect 34718 14164 34752 14198
rect 34718 14074 34752 14108
rect 34718 13984 34752 14018
rect 34718 13894 34752 13928
rect 34718 13804 34752 13838
rect 33906 13710 33940 13744
rect 33996 13710 34030 13744
rect 34086 13710 34120 13744
rect 34176 13710 34210 13744
rect 34266 13710 34300 13744
rect 34356 13710 34390 13744
rect 34446 13710 34480 13744
rect 34536 13710 34570 13744
rect 34626 13710 34660 13744
rect 35280 14600 35314 14634
rect 35370 14600 35404 14634
rect 35460 14600 35494 14634
rect 35550 14600 35584 14634
rect 35640 14600 35674 14634
rect 35730 14600 35764 14634
rect 35820 14600 35854 14634
rect 35910 14600 35944 14634
rect 36000 14600 36034 14634
rect 35168 14543 35202 14577
rect 36058 14524 36092 14558
rect 35168 14453 35202 14487
rect 35168 14363 35202 14397
rect 35168 14273 35202 14307
rect 35168 14183 35202 14217
rect 35168 14093 35202 14127
rect 35168 14003 35202 14037
rect 35168 13913 35202 13947
rect 35168 13823 35202 13857
rect 36058 14434 36092 14468
rect 36058 14344 36092 14378
rect 36058 14254 36092 14288
rect 36058 14164 36092 14198
rect 36058 14074 36092 14108
rect 36058 13984 36092 14018
rect 36058 13894 36092 13928
rect 36058 13804 36092 13838
rect 35246 13710 35280 13744
rect 35336 13710 35370 13744
rect 35426 13710 35460 13744
rect 35516 13710 35550 13744
rect 35606 13710 35640 13744
rect 35696 13710 35730 13744
rect 35786 13710 35820 13744
rect 35876 13710 35910 13744
rect 35966 13710 36000 13744
rect 36620 14600 36654 14634
rect 36710 14600 36744 14634
rect 36800 14600 36834 14634
rect 36890 14600 36924 14634
rect 36980 14600 37014 14634
rect 37070 14600 37104 14634
rect 37160 14600 37194 14634
rect 37250 14600 37284 14634
rect 37340 14600 37374 14634
rect 36508 14543 36542 14577
rect 37398 14524 37432 14558
rect 36508 14453 36542 14487
rect 36508 14363 36542 14397
rect 36508 14273 36542 14307
rect 36508 14183 36542 14217
rect 36508 14093 36542 14127
rect 36508 14003 36542 14037
rect 36508 13913 36542 13947
rect 36508 13823 36542 13857
rect 37398 14434 37432 14468
rect 37398 14344 37432 14378
rect 37398 14254 37432 14288
rect 37398 14164 37432 14198
rect 37398 14074 37432 14108
rect 37398 13984 37432 14018
rect 37398 13894 37432 13928
rect 37398 13804 37432 13838
rect 36586 13710 36620 13744
rect 36676 13710 36710 13744
rect 36766 13710 36800 13744
rect 36856 13710 36890 13744
rect 36946 13710 36980 13744
rect 37036 13710 37070 13744
rect 37126 13710 37160 13744
rect 37216 13710 37250 13744
rect 37306 13710 37340 13744
rect 37960 14600 37994 14634
rect 38050 14600 38084 14634
rect 38140 14600 38174 14634
rect 38230 14600 38264 14634
rect 38320 14600 38354 14634
rect 38410 14600 38444 14634
rect 38500 14600 38534 14634
rect 38590 14600 38624 14634
rect 38680 14600 38714 14634
rect 37848 14543 37882 14577
rect 38738 14524 38772 14558
rect 37848 14453 37882 14487
rect 37848 14363 37882 14397
rect 37848 14273 37882 14307
rect 37848 14183 37882 14217
rect 37848 14093 37882 14127
rect 37848 14003 37882 14037
rect 37848 13913 37882 13947
rect 37848 13823 37882 13857
rect 38738 14434 38772 14468
rect 38738 14344 38772 14378
rect 38738 14254 38772 14288
rect 38738 14164 38772 14198
rect 38738 14074 38772 14108
rect 38738 13984 38772 14018
rect 38738 13894 38772 13928
rect 38738 13804 38772 13838
rect 37926 13710 37960 13744
rect 38016 13710 38050 13744
rect 38106 13710 38140 13744
rect 38196 13710 38230 13744
rect 38286 13710 38320 13744
rect 38376 13710 38410 13744
rect 38466 13710 38500 13744
rect 38556 13710 38590 13744
rect 38646 13710 38680 13744
<< poly >>
rect 15123 41197 15523 41223
rect 15581 41197 15981 41223
rect 16039 41197 16439 41223
rect 16497 41197 16897 41223
rect 16955 41197 17355 41223
rect 17413 41197 17813 41223
rect 17871 41197 18271 41223
rect 18329 41197 18729 41223
rect 18787 41197 19187 41223
rect 19245 41197 19645 41223
rect 19703 41197 20103 41223
rect 20161 41197 20561 41223
rect 20619 41197 21019 41223
rect 21077 41197 21477 41223
rect 21535 41197 21935 41223
rect 21993 41197 22393 41223
rect 22451 41197 22851 41223
rect 22909 41197 23309 41223
rect 23367 41197 23767 41223
rect 23825 41197 24225 41223
rect 24283 41197 24683 41223
rect 24741 41197 25141 41223
rect 25199 41197 25599 41223
rect 25657 41197 26057 41223
rect 26115 41197 26515 41223
rect 26573 41197 26973 41223
rect 27031 41197 27431 41223
rect 27489 41197 27889 41223
rect 27947 41197 28347 41223
rect 28405 41197 28805 41223
rect 28863 41197 29263 41223
rect 29321 41197 29721 41223
rect 29779 41197 30179 41223
rect 30237 41197 30637 41223
rect 30695 41197 31095 41223
rect 31153 41197 31553 41223
rect 31611 41197 32011 41223
rect 32069 41197 32469 41223
rect 32527 41197 32927 41223
rect 32985 41197 33385 41223
rect 33443 41197 33843 41223
rect 33901 41197 34301 41223
rect 34359 41197 34759 41223
rect 34817 41197 35217 41223
rect 35275 41197 35675 41223
rect 35733 41197 36133 41223
rect 36191 41197 36591 41223
rect 36649 41197 37049 41223
rect 37107 41197 37507 41223
rect 37565 41197 37965 41223
rect 38023 41197 38423 41223
rect 38481 41197 38881 41223
rect 38939 41197 39339 41223
rect 39397 41197 39797 41223
rect 39855 41197 40255 41223
rect 40313 41197 40713 41223
rect 40771 41197 41171 41223
rect 41229 41197 41629 41223
rect 41687 41197 42087 41223
rect 42145 41197 42545 41223
rect 6042 40952 6442 40978
rect 6042 40126 6442 40152
rect 6190 39776 6310 40126
rect 15123 39881 15523 39907
rect 15581 39881 15981 39907
rect 16039 39881 16439 39907
rect 16497 39881 16897 39907
rect 16955 39881 17355 39907
rect 17413 39881 17813 39907
rect 17871 39881 18271 39907
rect 18329 39881 18729 39907
rect 18787 39881 19187 39907
rect 19245 39881 19645 39907
rect 19703 39881 20103 39907
rect 20161 39881 20561 39907
rect 20619 39881 21019 39907
rect 21077 39881 21477 39907
rect 21535 39881 21935 39907
rect 21993 39881 22393 39907
rect 22451 39881 22851 39907
rect 22909 39881 23309 39907
rect 23367 39881 23767 39907
rect 23825 39881 24225 39907
rect 24283 39881 24683 39907
rect 24741 39881 25141 39907
rect 25199 39881 25599 39907
rect 25657 39881 26057 39907
rect 26115 39881 26515 39907
rect 26573 39881 26973 39907
rect 27031 39881 27431 39907
rect 27489 39881 27889 39907
rect 27947 39881 28347 39907
rect 28405 39881 28805 39907
rect 28863 39881 29263 39907
rect 29321 39881 29721 39907
rect 29779 39881 30179 39907
rect 30237 39881 30637 39907
rect 30695 39881 31095 39907
rect 31153 39881 31553 39907
rect 31611 39881 32011 39907
rect 32069 39881 32469 39907
rect 32527 39881 32927 39907
rect 32985 39881 33385 39907
rect 33443 39881 33843 39907
rect 33901 39881 34301 39907
rect 34359 39881 34759 39907
rect 34817 39881 35217 39907
rect 35275 39881 35675 39907
rect 35733 39881 36133 39907
rect 36191 39881 36591 39907
rect 36649 39881 37049 39907
rect 37107 39881 37507 39907
rect 37565 39881 37965 39907
rect 38023 39881 38423 39907
rect 38481 39881 38881 39907
rect 38939 39881 39339 39907
rect 39397 39881 39797 39907
rect 39855 39881 40255 39907
rect 40313 39881 40713 39907
rect 40771 39881 41171 39907
rect 41229 39881 41629 39907
rect 41687 39881 42087 39907
rect 42145 39881 42545 39907
rect 6064 39743 6500 39776
rect 6064 39709 6167 39743
rect 6201 39709 6500 39743
rect 15270 39736 15390 39881
rect 15726 39736 15846 39881
rect 16182 39736 16302 39881
rect 16638 39736 16758 39881
rect 17094 39736 17214 39881
rect 17550 39736 17670 39881
rect 18006 39736 18126 39881
rect 18462 39736 18582 39881
rect 18918 39736 19038 39881
rect 19374 39736 19494 39881
rect 19830 39736 19950 39881
rect 20286 39736 20406 39881
rect 20742 39736 20862 39881
rect 21198 39736 21318 39881
rect 21654 39736 21774 39881
rect 22110 39736 22230 39881
rect 22566 39736 22686 39881
rect 23022 39736 23142 39881
rect 23478 39736 23598 39881
rect 23934 39736 24054 39881
rect 24390 39736 24510 39881
rect 24846 39736 24966 39881
rect 25302 39736 25422 39881
rect 25758 39736 25878 39881
rect 26214 39736 26334 39881
rect 26670 39736 26790 39881
rect 27126 39736 27246 39881
rect 27582 39736 27702 39881
rect 28038 39736 28158 39881
rect 28494 39736 28614 39881
rect 28950 39736 29070 39881
rect 29406 39736 29526 39881
rect 29862 39736 29982 39881
rect 30318 39736 30438 39881
rect 30774 39736 30894 39881
rect 31230 39736 31350 39881
rect 31686 39736 31806 39881
rect 32142 39736 32262 39881
rect 32598 39736 32718 39881
rect 33054 39736 33174 39881
rect 33510 39736 33630 39881
rect 33966 39736 34086 39881
rect 34422 39736 34542 39881
rect 34878 39736 34998 39881
rect 35334 39736 35454 39881
rect 35790 39736 35910 39881
rect 36246 39736 36366 39881
rect 36702 39736 36822 39881
rect 37158 39736 37278 39881
rect 37614 39736 37734 39881
rect 38070 39736 38190 39881
rect 38526 39736 38646 39881
rect 38982 39736 39102 39881
rect 39438 39736 39558 39881
rect 39894 39736 40014 39881
rect 40350 39736 40470 39881
rect 40806 39736 40926 39881
rect 41262 39736 41382 39881
rect 41718 39736 41838 39881
rect 42174 39736 42294 39881
rect 6064 39676 6500 39709
rect 15030 39703 42638 39736
rect 15030 39669 15213 39703
rect 15247 39669 15613 39703
rect 15647 39669 16013 39703
rect 16047 39669 16413 39703
rect 16447 39669 16813 39703
rect 16847 39669 17213 39703
rect 17247 39669 17613 39703
rect 17647 39669 18013 39703
rect 18047 39669 18413 39703
rect 18447 39669 18813 39703
rect 18847 39669 19213 39703
rect 19247 39669 19613 39703
rect 19647 39669 20013 39703
rect 20047 39669 20413 39703
rect 20447 39669 20813 39703
rect 20847 39669 21213 39703
rect 21247 39669 21613 39703
rect 21647 39669 22013 39703
rect 22047 39669 22413 39703
rect 22447 39669 22813 39703
rect 22847 39669 23213 39703
rect 23247 39669 23613 39703
rect 23647 39669 24013 39703
rect 24047 39669 24413 39703
rect 24447 39669 24813 39703
rect 24847 39669 25213 39703
rect 25247 39669 25613 39703
rect 25647 39669 26013 39703
rect 26047 39669 26413 39703
rect 26447 39669 26813 39703
rect 26847 39669 27213 39703
rect 27247 39669 27613 39703
rect 27647 39669 28013 39703
rect 28047 39669 28413 39703
rect 28447 39669 28813 39703
rect 28847 39669 29213 39703
rect 29247 39669 29613 39703
rect 29647 39669 30013 39703
rect 30047 39669 30413 39703
rect 30447 39669 30813 39703
rect 30847 39669 31213 39703
rect 31247 39669 31613 39703
rect 31647 39669 32013 39703
rect 32047 39669 32413 39703
rect 32447 39669 32813 39703
rect 32847 39669 33213 39703
rect 33247 39669 33613 39703
rect 33647 39669 34013 39703
rect 34047 39669 34413 39703
rect 34447 39669 34813 39703
rect 34847 39669 35213 39703
rect 35247 39669 35613 39703
rect 35647 39669 36013 39703
rect 36047 39669 36413 39703
rect 36447 39669 36813 39703
rect 36847 39669 37213 39703
rect 37247 39669 37613 39703
rect 37647 39669 38013 39703
rect 38047 39669 38413 39703
rect 38447 39669 38813 39703
rect 38847 39669 39213 39703
rect 39247 39669 39613 39703
rect 39647 39669 40013 39703
rect 40047 39669 40413 39703
rect 40447 39669 40813 39703
rect 40847 39669 41213 39703
rect 41247 39669 41613 39703
rect 41647 39669 42013 39703
rect 42047 39669 42413 39703
rect 42447 39669 42638 39703
rect 15030 39636 42638 39669
rect 28386 37192 28786 37218
rect 28386 36366 28786 36392
rect 28534 36016 28654 36366
rect 28408 35983 28844 36016
rect 28408 35949 28511 35983
rect 28545 35949 28844 35983
rect 28408 35916 28844 35949
rect 14241 33677 14641 33703
rect 14699 33677 15099 33703
rect 15157 33677 15557 33703
rect 15615 33677 16015 33703
rect 16073 33677 16473 33703
rect 16531 33677 16931 33703
rect 16989 33677 17389 33703
rect 17447 33677 17847 33703
rect 17905 33677 18305 33703
rect 18363 33677 18763 33703
rect 18821 33677 19221 33703
rect 19279 33677 19679 33703
rect 19737 33677 20137 33703
rect 20195 33677 20595 33703
rect 20653 33677 21053 33703
rect 21111 33677 21511 33703
rect 21569 33677 21969 33703
rect 22027 33677 22427 33703
rect 22485 33677 22885 33703
rect 22943 33677 23343 33703
rect 23401 33677 23801 33703
rect 23859 33677 24259 33703
rect 24317 33677 24717 33703
rect 24775 33677 25175 33703
rect 25233 33677 25633 33703
rect 25691 33677 26091 33703
rect 26149 33677 26549 33703
rect 26607 33677 27007 33703
rect 27065 33677 27465 33703
rect 27523 33677 27923 33703
rect 27981 33677 28381 33703
rect 28439 33677 28839 33703
rect 28897 33677 29297 33703
rect 29355 33677 29755 33703
rect 29813 33677 30213 33703
rect 30271 33677 30671 33703
rect 30729 33677 31129 33703
rect 31187 33677 31587 33703
rect 31645 33677 32045 33703
rect 32103 33677 32503 33703
rect 32561 33677 32961 33703
rect 33019 33677 33419 33703
rect 33477 33677 33877 33703
rect 33935 33677 34335 33703
rect 34393 33677 34793 33703
rect 34851 33677 35251 33703
rect 35309 33677 35709 33703
rect 35767 33677 36167 33703
rect 36225 33677 36625 33703
rect 36683 33677 37083 33703
rect 37141 33677 37541 33703
rect 37599 33677 37999 33703
rect 38057 33677 38457 33703
rect 38515 33677 38915 33703
rect 38973 33677 39373 33703
rect 39431 33677 39831 33703
rect 39889 33677 40289 33703
rect 40347 33677 40747 33703
rect 40805 33677 41205 33703
rect 41263 33677 41663 33703
rect 14241 32361 14641 32387
rect 14699 32361 15099 32387
rect 15157 32361 15557 32387
rect 15615 32361 16015 32387
rect 16073 32361 16473 32387
rect 16531 32361 16931 32387
rect 16989 32361 17389 32387
rect 17447 32361 17847 32387
rect 17905 32361 18305 32387
rect 18363 32361 18763 32387
rect 18821 32361 19221 32387
rect 19279 32361 19679 32387
rect 19737 32361 20137 32387
rect 20195 32361 20595 32387
rect 20653 32361 21053 32387
rect 21111 32361 21511 32387
rect 21569 32361 21969 32387
rect 22027 32361 22427 32387
rect 22485 32361 22885 32387
rect 22943 32361 23343 32387
rect 23401 32361 23801 32387
rect 23859 32361 24259 32387
rect 24317 32361 24717 32387
rect 24775 32361 25175 32387
rect 25233 32361 25633 32387
rect 25691 32361 26091 32387
rect 26149 32361 26549 32387
rect 26607 32361 27007 32387
rect 27065 32361 27465 32387
rect 27523 32361 27923 32387
rect 27981 32361 28381 32387
rect 28439 32361 28839 32387
rect 28897 32361 29297 32387
rect 29355 32361 29755 32387
rect 29813 32361 30213 32387
rect 30271 32361 30671 32387
rect 30729 32361 31129 32387
rect 31187 32361 31587 32387
rect 31645 32361 32045 32387
rect 32103 32361 32503 32387
rect 32561 32361 32961 32387
rect 33019 32361 33419 32387
rect 33477 32361 33877 32387
rect 33935 32361 34335 32387
rect 34393 32361 34793 32387
rect 34851 32361 35251 32387
rect 35309 32361 35709 32387
rect 35767 32361 36167 32387
rect 36225 32361 36625 32387
rect 36683 32361 37083 32387
rect 37141 32361 37541 32387
rect 37599 32361 37999 32387
rect 38057 32361 38457 32387
rect 38515 32361 38915 32387
rect 38973 32361 39373 32387
rect 39431 32361 39831 32387
rect 39889 32361 40289 32387
rect 40347 32361 40747 32387
rect 40805 32361 41205 32387
rect 41263 32361 41663 32387
rect 14388 32216 14508 32361
rect 14844 32216 14964 32361
rect 15300 32216 15420 32361
rect 15756 32216 15876 32361
rect 16212 32216 16332 32361
rect 16668 32216 16788 32361
rect 17124 32216 17244 32361
rect 17580 32216 17700 32361
rect 18036 32216 18156 32361
rect 18492 32216 18612 32361
rect 18948 32216 19068 32361
rect 19404 32216 19524 32361
rect 19860 32216 19980 32361
rect 20316 32216 20436 32361
rect 20772 32216 20892 32361
rect 21228 32216 21348 32361
rect 21684 32216 21804 32361
rect 22140 32216 22260 32361
rect 22596 32216 22716 32361
rect 23052 32216 23172 32361
rect 23508 32216 23628 32361
rect 23964 32216 24084 32361
rect 24420 32216 24540 32361
rect 24876 32216 24996 32361
rect 25332 32216 25452 32361
rect 25788 32216 25908 32361
rect 26244 32216 26364 32361
rect 26700 32216 26820 32361
rect 27156 32216 27276 32361
rect 27612 32216 27732 32361
rect 28068 32216 28188 32361
rect 28524 32216 28644 32361
rect 28980 32216 29100 32361
rect 29436 32216 29556 32361
rect 29892 32216 30012 32361
rect 30348 32216 30468 32361
rect 30804 32216 30924 32361
rect 31260 32216 31380 32361
rect 31716 32216 31836 32361
rect 32172 32216 32292 32361
rect 32628 32216 32748 32361
rect 33084 32216 33204 32361
rect 33540 32216 33660 32361
rect 33996 32216 34116 32361
rect 34452 32216 34572 32361
rect 34908 32216 35028 32361
rect 35364 32216 35484 32361
rect 35820 32216 35940 32361
rect 36276 32216 36396 32361
rect 36732 32216 36852 32361
rect 37188 32216 37308 32361
rect 37644 32216 37764 32361
rect 38100 32216 38220 32361
rect 38556 32216 38676 32361
rect 39012 32216 39132 32361
rect 39468 32216 39588 32361
rect 39924 32216 40044 32361
rect 40380 32216 40500 32361
rect 40836 32216 40956 32361
rect 41292 32216 41412 32361
rect 14148 32183 41756 32216
rect 14148 32149 14331 32183
rect 14365 32149 14731 32183
rect 14765 32149 15131 32183
rect 15165 32149 15531 32183
rect 15565 32149 15931 32183
rect 15965 32149 16331 32183
rect 16365 32149 16731 32183
rect 16765 32149 17131 32183
rect 17165 32149 17531 32183
rect 17565 32149 17931 32183
rect 17965 32149 18331 32183
rect 18365 32149 18731 32183
rect 18765 32149 19131 32183
rect 19165 32149 19531 32183
rect 19565 32149 19931 32183
rect 19965 32149 20331 32183
rect 20365 32149 20731 32183
rect 20765 32149 21131 32183
rect 21165 32149 21531 32183
rect 21565 32149 21931 32183
rect 21965 32149 22331 32183
rect 22365 32149 22731 32183
rect 22765 32149 23131 32183
rect 23165 32149 23531 32183
rect 23565 32149 23931 32183
rect 23965 32149 24331 32183
rect 24365 32149 24731 32183
rect 24765 32149 25131 32183
rect 25165 32149 25531 32183
rect 25565 32149 25931 32183
rect 25965 32149 26331 32183
rect 26365 32149 26731 32183
rect 26765 32149 27131 32183
rect 27165 32149 27531 32183
rect 27565 32149 27931 32183
rect 27965 32149 28331 32183
rect 28365 32149 28731 32183
rect 28765 32149 29131 32183
rect 29165 32149 29531 32183
rect 29565 32149 29931 32183
rect 29965 32149 30331 32183
rect 30365 32149 30731 32183
rect 30765 32149 31131 32183
rect 31165 32149 31531 32183
rect 31565 32149 31931 32183
rect 31965 32149 32331 32183
rect 32365 32149 32731 32183
rect 32765 32149 33131 32183
rect 33165 32149 33531 32183
rect 33565 32149 33931 32183
rect 33965 32149 34331 32183
rect 34365 32149 34731 32183
rect 34765 32149 35131 32183
rect 35165 32149 35531 32183
rect 35565 32149 35931 32183
rect 35965 32149 36331 32183
rect 36365 32149 36731 32183
rect 36765 32149 37131 32183
rect 37165 32149 37531 32183
rect 37565 32149 37931 32183
rect 37965 32149 38331 32183
rect 38365 32149 38731 32183
rect 38765 32149 39131 32183
rect 39165 32149 39531 32183
rect 39565 32149 39931 32183
rect 39965 32149 40331 32183
rect 40365 32149 40731 32183
rect 40765 32149 41131 32183
rect 41165 32149 41531 32183
rect 41565 32149 41756 32183
rect 14148 32116 41756 32149
rect 6107 29917 6507 29943
rect 6565 29917 6965 29943
rect 7023 29917 7423 29943
rect 7481 29917 7881 29943
rect 7939 29917 8339 29943
rect 8397 29917 8797 29943
rect 8855 29917 9255 29943
rect 9313 29917 9713 29943
rect 9771 29917 10171 29943
rect 10229 29917 10629 29943
rect 10687 29917 11087 29943
rect 11145 29917 11545 29943
rect 11603 29917 12003 29943
rect 12061 29917 12461 29943
rect 12519 29917 12919 29943
rect 12977 29917 13377 29943
rect 13435 29917 13835 29943
rect 13893 29917 14293 29943
rect 14351 29917 14751 29943
rect 14809 29917 15209 29943
rect 15267 29917 15667 29943
rect 15725 29917 16125 29943
rect 16183 29917 16583 29943
rect 16641 29917 17041 29943
rect 17099 29917 17499 29943
rect 17557 29917 17957 29943
rect 18015 29917 18415 29943
rect 18473 29917 18873 29943
rect 18931 29917 19331 29943
rect 19389 29917 19789 29943
rect 19847 29917 20247 29943
rect 20305 29917 20705 29943
rect 20763 29917 21163 29943
rect 21221 29917 21621 29943
rect 21679 29917 22079 29943
rect 22137 29917 22537 29943
rect 22595 29917 22995 29943
rect 23053 29917 23453 29943
rect 23511 29917 23911 29943
rect 23969 29917 24369 29943
rect 24427 29917 24827 29943
rect 24885 29917 25285 29943
rect 25343 29917 25743 29943
rect 25801 29917 26201 29943
rect 26259 29917 26659 29943
rect 26717 29917 27117 29943
rect 27175 29917 27575 29943
rect 27633 29917 28033 29943
rect 28091 29917 28491 29943
rect 28549 29917 28949 29943
rect 29007 29917 29407 29943
rect 29465 29917 29865 29943
rect 29923 29917 30323 29943
rect 30381 29917 30781 29943
rect 30839 29917 31239 29943
rect 31297 29917 31697 29943
rect 31755 29917 32155 29943
rect 32213 29917 32613 29943
rect 32671 29917 33071 29943
rect 33129 29917 33529 29943
rect 34135 29917 34535 29943
rect 34593 29917 34993 29943
rect 35051 29917 35451 29943
rect 35509 29917 35909 29943
rect 35967 29917 36367 29943
rect 36425 29917 36825 29943
rect 6107 28601 6507 28627
rect 6565 28601 6965 28627
rect 7023 28601 7423 28627
rect 7481 28601 7881 28627
rect 7939 28601 8339 28627
rect 8397 28601 8797 28627
rect 8855 28601 9255 28627
rect 9313 28601 9713 28627
rect 9771 28601 10171 28627
rect 10229 28601 10629 28627
rect 10687 28601 11087 28627
rect 11145 28601 11545 28627
rect 11603 28601 12003 28627
rect 12061 28601 12461 28627
rect 12519 28601 12919 28627
rect 12977 28601 13377 28627
rect 13435 28601 13835 28627
rect 13893 28601 14293 28627
rect 14351 28601 14751 28627
rect 14809 28601 15209 28627
rect 15267 28601 15667 28627
rect 15725 28601 16125 28627
rect 16183 28601 16583 28627
rect 16641 28601 17041 28627
rect 17099 28601 17499 28627
rect 17557 28601 17957 28627
rect 18015 28601 18415 28627
rect 18473 28601 18873 28627
rect 18931 28601 19331 28627
rect 19389 28601 19789 28627
rect 19847 28601 20247 28627
rect 20305 28601 20705 28627
rect 20763 28601 21163 28627
rect 21221 28601 21621 28627
rect 21679 28601 22079 28627
rect 22137 28601 22537 28627
rect 22595 28601 22995 28627
rect 23053 28601 23453 28627
rect 23511 28601 23911 28627
rect 23969 28601 24369 28627
rect 24427 28601 24827 28627
rect 24885 28601 25285 28627
rect 25343 28601 25743 28627
rect 25801 28601 26201 28627
rect 26259 28601 26659 28627
rect 26717 28601 27117 28627
rect 27175 28601 27575 28627
rect 27633 28601 28033 28627
rect 28091 28601 28491 28627
rect 28549 28601 28949 28627
rect 29007 28601 29407 28627
rect 29465 28601 29865 28627
rect 29923 28601 30323 28627
rect 30381 28601 30781 28627
rect 30839 28601 31239 28627
rect 31297 28601 31697 28627
rect 31755 28601 32155 28627
rect 32213 28601 32613 28627
rect 32671 28601 33071 28627
rect 33129 28601 33529 28627
rect 34135 28601 34535 28627
rect 34593 28601 34993 28627
rect 35051 28601 35451 28627
rect 35509 28601 35909 28627
rect 35967 28601 36367 28627
rect 36425 28601 36825 28627
rect 6254 28456 6374 28601
rect 6710 28456 6830 28601
rect 7166 28456 7286 28601
rect 7622 28456 7742 28601
rect 8078 28456 8198 28601
rect 8534 28456 8654 28601
rect 8990 28456 9110 28601
rect 9446 28456 9566 28601
rect 9902 28456 10022 28601
rect 10358 28456 10478 28601
rect 10814 28456 10934 28601
rect 11270 28456 11390 28601
rect 11726 28456 11846 28601
rect 12182 28456 12302 28601
rect 12638 28456 12758 28601
rect 13094 28456 13214 28601
rect 13550 28456 13670 28601
rect 14006 28456 14126 28601
rect 14462 28456 14582 28601
rect 14918 28456 15038 28601
rect 15374 28456 15494 28601
rect 15830 28456 15950 28601
rect 16286 28456 16406 28601
rect 16742 28456 16862 28601
rect 17198 28456 17318 28601
rect 17654 28456 17774 28601
rect 18110 28456 18230 28601
rect 18566 28456 18686 28601
rect 19022 28456 19142 28601
rect 19478 28456 19598 28601
rect 19934 28456 20054 28601
rect 20390 28456 20510 28601
rect 20846 28456 20966 28601
rect 21302 28456 21422 28601
rect 21758 28456 21878 28601
rect 22214 28456 22334 28601
rect 22670 28456 22790 28601
rect 23126 28456 23246 28601
rect 23582 28456 23702 28601
rect 24038 28456 24158 28601
rect 24494 28456 24614 28601
rect 24950 28456 25070 28601
rect 25406 28456 25526 28601
rect 25862 28456 25982 28601
rect 26318 28456 26438 28601
rect 26774 28456 26894 28601
rect 27230 28456 27350 28601
rect 27686 28456 27806 28601
rect 28142 28456 28262 28601
rect 28598 28456 28718 28601
rect 29054 28456 29174 28601
rect 29510 28456 29630 28601
rect 29966 28456 30086 28601
rect 30422 28456 30542 28601
rect 30878 28456 30998 28601
rect 31334 28456 31454 28601
rect 31790 28456 31910 28601
rect 32246 28456 32366 28601
rect 32702 28456 32822 28601
rect 33158 28456 33278 28601
rect 34282 28456 34402 28601
rect 34738 28456 34858 28601
rect 35194 28456 35314 28601
rect 35650 28456 35770 28601
rect 36106 28456 36226 28601
rect 36562 28456 36682 28601
rect 6014 28423 33622 28456
rect 6014 28389 6197 28423
rect 6231 28389 6597 28423
rect 6631 28389 6997 28423
rect 7031 28389 7397 28423
rect 7431 28389 7797 28423
rect 7831 28389 8197 28423
rect 8231 28389 8597 28423
rect 8631 28389 8997 28423
rect 9031 28389 9397 28423
rect 9431 28389 9797 28423
rect 9831 28389 10197 28423
rect 10231 28389 10597 28423
rect 10631 28389 10997 28423
rect 11031 28389 11397 28423
rect 11431 28389 11797 28423
rect 11831 28389 12197 28423
rect 12231 28389 12597 28423
rect 12631 28389 12997 28423
rect 13031 28389 13397 28423
rect 13431 28389 13797 28423
rect 13831 28389 14197 28423
rect 14231 28389 14597 28423
rect 14631 28389 14997 28423
rect 15031 28389 15397 28423
rect 15431 28389 15797 28423
rect 15831 28389 16197 28423
rect 16231 28389 16597 28423
rect 16631 28389 16997 28423
rect 17031 28389 17397 28423
rect 17431 28389 17797 28423
rect 17831 28389 18197 28423
rect 18231 28389 18597 28423
rect 18631 28389 18997 28423
rect 19031 28389 19397 28423
rect 19431 28389 19797 28423
rect 19831 28389 20197 28423
rect 20231 28389 20597 28423
rect 20631 28389 20997 28423
rect 21031 28389 21397 28423
rect 21431 28389 21797 28423
rect 21831 28389 22197 28423
rect 22231 28389 22597 28423
rect 22631 28389 22997 28423
rect 23031 28389 23397 28423
rect 23431 28389 23797 28423
rect 23831 28389 24197 28423
rect 24231 28389 24597 28423
rect 24631 28389 24997 28423
rect 25031 28389 25397 28423
rect 25431 28389 25797 28423
rect 25831 28389 26197 28423
rect 26231 28389 26597 28423
rect 26631 28389 26997 28423
rect 27031 28389 27397 28423
rect 27431 28389 27797 28423
rect 27831 28389 28197 28423
rect 28231 28389 28597 28423
rect 28631 28389 28997 28423
rect 29031 28389 29397 28423
rect 29431 28389 29797 28423
rect 29831 28389 30197 28423
rect 30231 28389 30597 28423
rect 30631 28389 30997 28423
rect 31031 28389 31397 28423
rect 31431 28389 31797 28423
rect 31831 28389 32197 28423
rect 32231 28389 32597 28423
rect 32631 28389 32997 28423
rect 33031 28389 33397 28423
rect 33431 28389 33622 28423
rect 6014 28356 33622 28389
rect 34042 28423 36918 28456
rect 34042 28389 34225 28423
rect 34259 28389 34625 28423
rect 34659 28389 35025 28423
rect 35059 28389 35425 28423
rect 35459 28389 35825 28423
rect 35859 28389 36225 28423
rect 36259 28389 36625 28423
rect 36659 28389 36918 28423
rect 34042 28356 36918 28389
rect 9635 26157 10035 26183
rect 10093 26157 10493 26183
rect 10551 26157 10951 26183
rect 11009 26157 11409 26183
rect 11467 26157 11867 26183
rect 11925 26157 12325 26183
rect 12383 26157 12783 26183
rect 12841 26157 13241 26183
rect 13299 26157 13699 26183
rect 13757 26157 14157 26183
rect 14215 26157 14615 26183
rect 14673 26157 15073 26183
rect 23026 25912 23426 25938
rect 23484 25912 23884 25938
rect 23942 25912 24342 25938
rect 24400 25912 24800 25938
rect 24858 25912 25258 25938
rect 25316 25912 25716 25938
rect 25774 25912 26174 25938
rect 26232 25912 26632 25938
rect 26690 25912 27090 25938
rect 23026 25086 23426 25112
rect 23484 25086 23884 25112
rect 23942 25086 24342 25112
rect 24400 25086 24800 25112
rect 24858 25086 25258 25112
rect 25316 25086 25716 25112
rect 25774 25086 26174 25112
rect 26232 25086 26632 25112
rect 26690 25086 27090 25112
rect 23174 24896 23294 25086
rect 23630 24896 23750 25086
rect 24086 24896 24206 25086
rect 24542 24896 24662 25086
rect 24998 24896 25118 25086
rect 25454 24896 25574 25086
rect 25910 24896 26030 25086
rect 26366 24896 26486 25086
rect 26822 24896 26942 25086
rect 9635 24841 10035 24867
rect 10093 24841 10493 24867
rect 10551 24841 10951 24867
rect 11009 24841 11409 24867
rect 11467 24841 11867 24867
rect 11925 24841 12325 24867
rect 12383 24841 12783 24867
rect 12841 24841 13241 24867
rect 13299 24841 13699 24867
rect 13757 24841 14157 24867
rect 14215 24841 14615 24867
rect 14673 24841 15073 24867
rect 23048 24863 27148 24896
rect 9782 24696 9902 24841
rect 10238 24696 10358 24841
rect 10694 24696 10814 24841
rect 11150 24696 11270 24841
rect 11606 24696 11726 24841
rect 12062 24696 12182 24841
rect 12518 24696 12638 24841
rect 12974 24696 13094 24841
rect 13430 24696 13550 24841
rect 13886 24696 14006 24841
rect 14342 24696 14462 24841
rect 14798 24696 14918 24841
rect 23048 24829 23151 24863
rect 23185 24829 23551 24863
rect 23585 24829 23951 24863
rect 23985 24829 24351 24863
rect 24385 24829 24751 24863
rect 24785 24829 25151 24863
rect 25185 24829 25551 24863
rect 25585 24829 25951 24863
rect 25985 24829 26351 24863
rect 26385 24829 26751 24863
rect 26785 24829 27148 24863
rect 23048 24796 27148 24829
rect 9542 24663 15166 24696
rect 9542 24629 9725 24663
rect 9759 24629 10125 24663
rect 10159 24629 10525 24663
rect 10559 24629 10925 24663
rect 10959 24629 11325 24663
rect 11359 24629 11725 24663
rect 11759 24629 12125 24663
rect 12159 24629 12525 24663
rect 12559 24629 12925 24663
rect 12959 24629 13325 24663
rect 13359 24629 13725 24663
rect 13759 24629 14125 24663
rect 14159 24629 14525 24663
rect 14559 24629 14925 24663
rect 14959 24629 15166 24663
rect 9542 24596 15166 24629
rect 7773 22397 8173 22423
rect 8231 22397 8631 22423
rect 8689 22397 9089 22423
rect 9147 22397 9547 22423
rect 9605 22397 10005 22423
rect 10063 22397 10463 22423
rect 10521 22397 10921 22423
rect 10979 22397 11379 22423
rect 11437 22397 11837 22423
rect 11895 22397 12295 22423
rect 12353 22397 12753 22423
rect 12811 22397 13211 22423
rect 23026 22152 23426 22178
rect 23484 22152 23884 22178
rect 23942 22152 24342 22178
rect 24400 22152 24800 22178
rect 24858 22152 25258 22178
rect 25316 22152 25716 22178
rect 25774 22152 26174 22178
rect 26232 22152 26632 22178
rect 26690 22152 27090 22178
rect 23026 21326 23426 21352
rect 23484 21326 23884 21352
rect 23942 21326 24342 21352
rect 24400 21326 24800 21352
rect 24858 21326 25258 21352
rect 25316 21326 25716 21352
rect 25774 21326 26174 21352
rect 26232 21326 26632 21352
rect 26690 21326 27090 21352
rect 23174 21136 23294 21326
rect 23630 21136 23750 21326
rect 24086 21136 24206 21326
rect 24542 21136 24662 21326
rect 24998 21136 25118 21326
rect 25454 21136 25574 21326
rect 25910 21136 26030 21326
rect 26366 21136 26486 21326
rect 26822 21136 26942 21326
rect 7773 21081 8173 21107
rect 8231 21081 8631 21107
rect 8689 21081 9089 21107
rect 9147 21081 9547 21107
rect 9605 21081 10005 21107
rect 10063 21081 10463 21107
rect 10521 21081 10921 21107
rect 10979 21081 11379 21107
rect 11437 21081 11837 21107
rect 11895 21081 12295 21107
rect 12353 21081 12753 21107
rect 12811 21081 13211 21107
rect 7920 20936 8040 21081
rect 8376 20936 8496 21081
rect 8832 20936 8952 21081
rect 9288 20936 9408 21081
rect 9744 20936 9864 21081
rect 10200 20936 10320 21081
rect 10656 20936 10776 21081
rect 11112 20936 11232 21081
rect 11568 20936 11688 21081
rect 12024 20936 12144 21081
rect 12480 20936 12600 21081
rect 12936 20936 13056 21081
rect 23048 21103 27148 21136
rect 23048 21069 23151 21103
rect 23185 21069 23551 21103
rect 23585 21069 23951 21103
rect 23985 21069 24351 21103
rect 24385 21069 24751 21103
rect 24785 21069 25151 21103
rect 25185 21069 25551 21103
rect 25585 21069 25951 21103
rect 25985 21069 26351 21103
rect 26385 21069 26751 21103
rect 26785 21069 27148 21103
rect 23048 21036 27148 21069
rect 7680 20903 13304 20936
rect 7680 20869 7863 20903
rect 7897 20869 8263 20903
rect 8297 20869 8663 20903
rect 8697 20869 9063 20903
rect 9097 20869 9463 20903
rect 9497 20869 9863 20903
rect 9897 20869 10263 20903
rect 10297 20869 10663 20903
rect 10697 20869 11063 20903
rect 11097 20869 11463 20903
rect 11497 20869 11863 20903
rect 11897 20869 12263 20903
rect 12297 20869 12663 20903
rect 12697 20869 13063 20903
rect 13097 20869 13304 20903
rect 7680 20836 13304 20869
rect 24041 18637 24441 18663
rect 24499 18637 24899 18663
rect 24957 18637 25357 18663
rect 25415 18637 25815 18663
rect 25873 18637 26273 18663
rect 26331 18637 26731 18663
rect 6072 18392 6472 18418
rect 6530 18392 6930 18418
rect 6988 18392 7388 18418
rect 7446 18392 7846 18418
rect 7904 18392 8304 18418
rect 8362 18392 8762 18418
rect 8820 18392 9220 18418
rect 9278 18392 9678 18418
rect 9736 18392 10136 18418
rect 6072 17566 6472 17592
rect 6530 17566 6930 17592
rect 6988 17566 7388 17592
rect 7446 17566 7846 17592
rect 7904 17566 8304 17592
rect 8362 17566 8762 17592
rect 8820 17566 9220 17592
rect 9278 17566 9678 17592
rect 9736 17566 10136 17592
rect 6220 17376 6340 17566
rect 6676 17376 6796 17566
rect 7132 17376 7252 17566
rect 7588 17376 7708 17566
rect 8044 17376 8164 17566
rect 8500 17376 8620 17566
rect 8956 17376 9076 17566
rect 9412 17376 9532 17566
rect 9868 17376 9988 17566
rect 6094 17343 10194 17376
rect 6094 17309 6197 17343
rect 6231 17309 6597 17343
rect 6631 17309 6997 17343
rect 7031 17309 7397 17343
rect 7431 17309 7797 17343
rect 7831 17309 8197 17343
rect 8231 17309 8597 17343
rect 8631 17309 8997 17343
rect 9031 17309 9397 17343
rect 9431 17309 9797 17343
rect 9831 17309 10194 17343
rect 6094 17276 10194 17309
rect 24041 17321 24441 17347
rect 24499 17321 24899 17347
rect 24957 17321 25357 17347
rect 25415 17321 25815 17347
rect 25873 17321 26273 17347
rect 26331 17321 26731 17347
rect 24188 17176 24308 17321
rect 24644 17176 24764 17321
rect 25100 17176 25220 17321
rect 25556 17176 25676 17321
rect 26012 17176 26132 17321
rect 26468 17176 26588 17321
rect 23948 17143 26824 17176
rect 23948 17109 24131 17143
rect 24165 17109 24531 17143
rect 24565 17109 24931 17143
rect 24965 17109 25331 17143
rect 25365 17109 25731 17143
rect 25765 17109 26131 17143
rect 26165 17109 26531 17143
rect 26565 17109 26824 17143
rect 23948 17076 26824 17109
<< polycont >>
rect 6167 39709 6201 39743
rect 15213 39669 15247 39703
rect 15613 39669 15647 39703
rect 16013 39669 16047 39703
rect 16413 39669 16447 39703
rect 16813 39669 16847 39703
rect 17213 39669 17247 39703
rect 17613 39669 17647 39703
rect 18013 39669 18047 39703
rect 18413 39669 18447 39703
rect 18813 39669 18847 39703
rect 19213 39669 19247 39703
rect 19613 39669 19647 39703
rect 20013 39669 20047 39703
rect 20413 39669 20447 39703
rect 20813 39669 20847 39703
rect 21213 39669 21247 39703
rect 21613 39669 21647 39703
rect 22013 39669 22047 39703
rect 22413 39669 22447 39703
rect 22813 39669 22847 39703
rect 23213 39669 23247 39703
rect 23613 39669 23647 39703
rect 24013 39669 24047 39703
rect 24413 39669 24447 39703
rect 24813 39669 24847 39703
rect 25213 39669 25247 39703
rect 25613 39669 25647 39703
rect 26013 39669 26047 39703
rect 26413 39669 26447 39703
rect 26813 39669 26847 39703
rect 27213 39669 27247 39703
rect 27613 39669 27647 39703
rect 28013 39669 28047 39703
rect 28413 39669 28447 39703
rect 28813 39669 28847 39703
rect 29213 39669 29247 39703
rect 29613 39669 29647 39703
rect 30013 39669 30047 39703
rect 30413 39669 30447 39703
rect 30813 39669 30847 39703
rect 31213 39669 31247 39703
rect 31613 39669 31647 39703
rect 32013 39669 32047 39703
rect 32413 39669 32447 39703
rect 32813 39669 32847 39703
rect 33213 39669 33247 39703
rect 33613 39669 33647 39703
rect 34013 39669 34047 39703
rect 34413 39669 34447 39703
rect 34813 39669 34847 39703
rect 35213 39669 35247 39703
rect 35613 39669 35647 39703
rect 36013 39669 36047 39703
rect 36413 39669 36447 39703
rect 36813 39669 36847 39703
rect 37213 39669 37247 39703
rect 37613 39669 37647 39703
rect 38013 39669 38047 39703
rect 38413 39669 38447 39703
rect 38813 39669 38847 39703
rect 39213 39669 39247 39703
rect 39613 39669 39647 39703
rect 40013 39669 40047 39703
rect 40413 39669 40447 39703
rect 40813 39669 40847 39703
rect 41213 39669 41247 39703
rect 41613 39669 41647 39703
rect 42013 39669 42047 39703
rect 42413 39669 42447 39703
rect 28511 35949 28545 35983
rect 14331 32149 14365 32183
rect 14731 32149 14765 32183
rect 15131 32149 15165 32183
rect 15531 32149 15565 32183
rect 15931 32149 15965 32183
rect 16331 32149 16365 32183
rect 16731 32149 16765 32183
rect 17131 32149 17165 32183
rect 17531 32149 17565 32183
rect 17931 32149 17965 32183
rect 18331 32149 18365 32183
rect 18731 32149 18765 32183
rect 19131 32149 19165 32183
rect 19531 32149 19565 32183
rect 19931 32149 19965 32183
rect 20331 32149 20365 32183
rect 20731 32149 20765 32183
rect 21131 32149 21165 32183
rect 21531 32149 21565 32183
rect 21931 32149 21965 32183
rect 22331 32149 22365 32183
rect 22731 32149 22765 32183
rect 23131 32149 23165 32183
rect 23531 32149 23565 32183
rect 23931 32149 23965 32183
rect 24331 32149 24365 32183
rect 24731 32149 24765 32183
rect 25131 32149 25165 32183
rect 25531 32149 25565 32183
rect 25931 32149 25965 32183
rect 26331 32149 26365 32183
rect 26731 32149 26765 32183
rect 27131 32149 27165 32183
rect 27531 32149 27565 32183
rect 27931 32149 27965 32183
rect 28331 32149 28365 32183
rect 28731 32149 28765 32183
rect 29131 32149 29165 32183
rect 29531 32149 29565 32183
rect 29931 32149 29965 32183
rect 30331 32149 30365 32183
rect 30731 32149 30765 32183
rect 31131 32149 31165 32183
rect 31531 32149 31565 32183
rect 31931 32149 31965 32183
rect 32331 32149 32365 32183
rect 32731 32149 32765 32183
rect 33131 32149 33165 32183
rect 33531 32149 33565 32183
rect 33931 32149 33965 32183
rect 34331 32149 34365 32183
rect 34731 32149 34765 32183
rect 35131 32149 35165 32183
rect 35531 32149 35565 32183
rect 35931 32149 35965 32183
rect 36331 32149 36365 32183
rect 36731 32149 36765 32183
rect 37131 32149 37165 32183
rect 37531 32149 37565 32183
rect 37931 32149 37965 32183
rect 38331 32149 38365 32183
rect 38731 32149 38765 32183
rect 39131 32149 39165 32183
rect 39531 32149 39565 32183
rect 39931 32149 39965 32183
rect 40331 32149 40365 32183
rect 40731 32149 40765 32183
rect 41131 32149 41165 32183
rect 41531 32149 41565 32183
rect 6197 28389 6231 28423
rect 6597 28389 6631 28423
rect 6997 28389 7031 28423
rect 7397 28389 7431 28423
rect 7797 28389 7831 28423
rect 8197 28389 8231 28423
rect 8597 28389 8631 28423
rect 8997 28389 9031 28423
rect 9397 28389 9431 28423
rect 9797 28389 9831 28423
rect 10197 28389 10231 28423
rect 10597 28389 10631 28423
rect 10997 28389 11031 28423
rect 11397 28389 11431 28423
rect 11797 28389 11831 28423
rect 12197 28389 12231 28423
rect 12597 28389 12631 28423
rect 12997 28389 13031 28423
rect 13397 28389 13431 28423
rect 13797 28389 13831 28423
rect 14197 28389 14231 28423
rect 14597 28389 14631 28423
rect 14997 28389 15031 28423
rect 15397 28389 15431 28423
rect 15797 28389 15831 28423
rect 16197 28389 16231 28423
rect 16597 28389 16631 28423
rect 16997 28389 17031 28423
rect 17397 28389 17431 28423
rect 17797 28389 17831 28423
rect 18197 28389 18231 28423
rect 18597 28389 18631 28423
rect 18997 28389 19031 28423
rect 19397 28389 19431 28423
rect 19797 28389 19831 28423
rect 20197 28389 20231 28423
rect 20597 28389 20631 28423
rect 20997 28389 21031 28423
rect 21397 28389 21431 28423
rect 21797 28389 21831 28423
rect 22197 28389 22231 28423
rect 22597 28389 22631 28423
rect 22997 28389 23031 28423
rect 23397 28389 23431 28423
rect 23797 28389 23831 28423
rect 24197 28389 24231 28423
rect 24597 28389 24631 28423
rect 24997 28389 25031 28423
rect 25397 28389 25431 28423
rect 25797 28389 25831 28423
rect 26197 28389 26231 28423
rect 26597 28389 26631 28423
rect 26997 28389 27031 28423
rect 27397 28389 27431 28423
rect 27797 28389 27831 28423
rect 28197 28389 28231 28423
rect 28597 28389 28631 28423
rect 28997 28389 29031 28423
rect 29397 28389 29431 28423
rect 29797 28389 29831 28423
rect 30197 28389 30231 28423
rect 30597 28389 30631 28423
rect 30997 28389 31031 28423
rect 31397 28389 31431 28423
rect 31797 28389 31831 28423
rect 32197 28389 32231 28423
rect 32597 28389 32631 28423
rect 32997 28389 33031 28423
rect 33397 28389 33431 28423
rect 34225 28389 34259 28423
rect 34625 28389 34659 28423
rect 35025 28389 35059 28423
rect 35425 28389 35459 28423
rect 35825 28389 35859 28423
rect 36225 28389 36259 28423
rect 36625 28389 36659 28423
rect 23151 24829 23185 24863
rect 23551 24829 23585 24863
rect 23951 24829 23985 24863
rect 24351 24829 24385 24863
rect 24751 24829 24785 24863
rect 25151 24829 25185 24863
rect 25551 24829 25585 24863
rect 25951 24829 25985 24863
rect 26351 24829 26385 24863
rect 26751 24829 26785 24863
rect 9725 24629 9759 24663
rect 10125 24629 10159 24663
rect 10525 24629 10559 24663
rect 10925 24629 10959 24663
rect 11325 24629 11359 24663
rect 11725 24629 11759 24663
rect 12125 24629 12159 24663
rect 12525 24629 12559 24663
rect 12925 24629 12959 24663
rect 13325 24629 13359 24663
rect 13725 24629 13759 24663
rect 14125 24629 14159 24663
rect 14525 24629 14559 24663
rect 14925 24629 14959 24663
rect 23151 21069 23185 21103
rect 23551 21069 23585 21103
rect 23951 21069 23985 21103
rect 24351 21069 24385 21103
rect 24751 21069 24785 21103
rect 25151 21069 25185 21103
rect 25551 21069 25585 21103
rect 25951 21069 25985 21103
rect 26351 21069 26385 21103
rect 26751 21069 26785 21103
rect 7863 20869 7897 20903
rect 8263 20869 8297 20903
rect 8663 20869 8697 20903
rect 9063 20869 9097 20903
rect 9463 20869 9497 20903
rect 9863 20869 9897 20903
rect 10263 20869 10297 20903
rect 10663 20869 10697 20903
rect 11063 20869 11097 20903
rect 11463 20869 11497 20903
rect 11863 20869 11897 20903
rect 12263 20869 12297 20903
rect 12663 20869 12697 20903
rect 13063 20869 13097 20903
rect 6197 17309 6231 17343
rect 6597 17309 6631 17343
rect 6997 17309 7031 17343
rect 7397 17309 7431 17343
rect 7797 17309 7831 17343
rect 8197 17309 8231 17343
rect 8597 17309 8631 17343
rect 8997 17309 9031 17343
rect 9397 17309 9431 17343
rect 9797 17309 9831 17343
rect 24131 17109 24165 17143
rect 24531 17109 24565 17143
rect 24931 17109 24965 17143
rect 25331 17109 25365 17143
rect 25731 17109 25765 17143
rect 26131 17109 26165 17143
rect 26531 17109 26565 17143
<< xpolycontact >>
rect 39746 36867 40178 37437
rect 41754 36867 42186 37437
rect 39746 35907 40178 36477
rect 41754 35907 42186 36477
rect 37394 29347 37826 29917
rect 39402 29347 39834 29917
rect 40138 29347 40570 29917
rect 42146 29347 42578 29917
rect 37394 28387 37826 28957
rect 39402 28387 39834 28957
rect 40138 28387 40570 28957
rect 42146 28387 42578 28957
rect 6720 25587 7152 26157
rect 8728 25587 9160 26157
rect 6720 24627 7152 25197
rect 8728 24627 9160 25197
rect 39746 25587 40178 26157
rect 41754 25587 42186 26157
rect 39746 24627 40178 25197
rect 41754 24627 42186 25197
rect 39746 21827 40178 22397
rect 41754 21827 42186 22397
rect 39746 20867 40178 21437
rect 41754 20867 42186 21437
rect 10640 18067 11072 18637
rect 12648 18067 13080 18637
rect 13384 18067 13816 18637
rect 15392 18067 15824 18637
rect 10640 17107 11072 17677
rect 12648 17107 13080 17677
rect 13384 17107 13816 17677
rect 15392 17107 15824 17677
rect 39256 18067 39688 18637
rect 41264 18067 41696 18637
rect 39256 17107 39688 17677
rect 41264 17107 41696 17677
rect 7896 14307 8328 14877
rect 9904 14307 10336 14877
rect 10640 14307 11072 14877
rect 12648 14307 13080 14877
rect 13384 14307 13816 14877
rect 15392 14307 15824 14877
rect 23576 14307 24008 14877
rect 25584 14307 26016 14877
rect 7896 13347 8328 13917
rect 9904 13347 10336 13917
rect 10640 13347 11072 13917
rect 12648 13347 13080 13917
rect 13384 13347 13816 13917
rect 15392 13347 15824 13917
rect 23576 13347 24008 13917
rect 25584 13347 26016 13917
rect 39256 14307 39688 14877
rect 41264 14307 41696 14877
rect 39256 13347 39688 13917
rect 41264 13347 41696 13917
rect 7896 10547 8328 11117
rect 9904 10547 10336 11117
rect 10640 10547 11072 11117
rect 12648 10547 13080 11117
rect 13384 10547 13816 11117
rect 15392 10547 15824 11117
rect 23577 10547 24009 11117
rect 26159 10547 26591 11117
rect 26908 10547 27340 11117
rect 28916 10547 29348 11117
rect 29652 10547 30084 11117
rect 31660 10547 32092 11117
rect 32396 10547 32828 11117
rect 34404 10547 34836 11117
rect 35140 10547 35572 11117
rect 37148 10547 37580 11117
rect 37884 10547 38316 11117
rect 39892 10547 40324 11117
rect 7896 9587 8328 10157
rect 9904 9587 10336 10157
rect 10640 9587 11072 10157
rect 12648 9587 13080 10157
rect 13384 9587 13816 10157
rect 15392 9587 15824 10157
rect 23577 9587 24009 10157
rect 26159 9587 26591 10157
rect 26908 9587 27340 10157
rect 28916 9587 29348 10157
rect 29652 9587 30084 10157
rect 31660 9587 32092 10157
rect 32396 9587 32828 10157
rect 34404 9587 34836 10157
rect 35140 9587 35572 10157
rect 37148 9587 37580 10157
rect 37884 9587 38316 10157
rect 39892 9587 40324 10157
rect 7896 6787 8328 7357
rect 9904 6787 10336 7357
rect 14267 6787 14699 7357
rect 16849 6787 17281 7357
rect 17598 6787 18030 7357
rect 19606 6787 20038 7357
rect 20342 6787 20774 7357
rect 22350 6787 22782 7357
rect 23086 6787 23518 7357
rect 25094 6787 25526 7357
rect 25830 6787 26262 7357
rect 27838 6787 28270 7357
rect 28574 6787 29006 7357
rect 30582 6787 31014 7357
rect 31318 6787 31750 7357
rect 33326 6787 33758 7357
rect 35140 6787 35572 7357
rect 37148 6787 37580 7357
rect 37884 6787 38316 7357
rect 39892 6787 40324 7357
rect 7896 5827 8328 6397
rect 9904 5827 10336 6397
rect 14267 5827 14699 6397
rect 16849 5827 17281 6397
rect 17598 5827 18030 6397
rect 19606 5827 20038 6397
rect 20342 5827 20774 6397
rect 22350 5827 22782 6397
rect 23086 5827 23518 6397
rect 25094 5827 25526 6397
rect 25830 5827 26262 6397
rect 27838 5827 28270 6397
rect 28574 5827 29006 6397
rect 30582 5827 31014 6397
rect 31318 5827 31750 6397
rect 33326 5827 33758 6397
rect 35140 5827 35572 6397
rect 37148 5827 37580 6397
rect 37884 5827 38316 6397
rect 39892 5827 40324 6397
<< xpolyres >>
rect 40178 36867 41754 37437
rect 40178 35907 41754 36477
rect 37826 29347 39402 29917
rect 40570 29347 42146 29917
rect 37826 28387 39402 28957
rect 40570 28387 42146 28957
rect 7152 25587 8728 26157
rect 7152 24627 8728 25197
rect 40178 25587 41754 26157
rect 40178 24627 41754 25197
rect 40178 21827 41754 22397
rect 40178 20867 41754 21437
rect 11072 18067 12648 18637
rect 13816 18067 15392 18637
rect 11072 17107 12648 17677
rect 13816 17107 15392 17677
rect 39688 18067 41264 18637
rect 39688 17107 41264 17677
rect 8328 14307 9904 14877
rect 11072 14307 12648 14877
rect 13816 14307 15392 14877
rect 24008 14307 25584 14877
rect 8328 13347 9904 13917
rect 11072 13347 12648 13917
rect 13816 13347 15392 13917
rect 24008 13347 25584 13917
rect 39688 14307 41264 14877
rect 39688 13347 41264 13917
rect 8328 10547 9904 11117
rect 11072 10547 12648 11117
rect 13816 10547 15392 11117
rect 24009 10547 26159 11117
rect 27340 10547 28916 11117
rect 30084 10547 31660 11117
rect 32828 10547 34404 11117
rect 35572 10547 37148 11117
rect 38316 10547 39892 11117
rect 8328 9587 9904 10157
rect 11072 9587 12648 10157
rect 13816 9587 15392 10157
rect 24009 9587 26159 10157
rect 27340 9587 28916 10157
rect 30084 9587 31660 10157
rect 32828 9587 34404 10157
rect 35572 9587 37148 10157
rect 38316 9587 39892 10157
rect 8328 6787 9904 7357
rect 14699 6787 16849 7357
rect 18030 6787 19606 7357
rect 20774 6787 22350 7357
rect 23518 6787 25094 7357
rect 26262 6787 27838 7357
rect 29006 6787 30582 7357
rect 31750 6787 33326 7357
rect 35572 6787 37148 7357
rect 38316 6787 39892 7357
rect 8328 5827 9904 6397
rect 14699 5827 16849 6397
rect 18030 5827 19606 6397
rect 20774 5827 22350 6397
rect 23518 5827 25094 6397
rect 26262 5827 27838 6397
rect 29006 5827 30582 6397
rect 31750 5827 33326 6397
rect 35572 5827 37148 6397
rect 38316 5827 39892 6397
<< locali >>
rect 5886 41449 6500 41462
rect 5886 41415 6167 41449
rect 6201 41415 6500 41449
rect 5886 41402 6500 41415
rect 6800 41449 13968 41462
rect 6800 41415 6983 41449
rect 7017 41415 7383 41449
rect 7417 41415 7783 41449
rect 7817 41415 8183 41449
rect 8217 41415 8583 41449
rect 8617 41415 8983 41449
rect 9017 41415 9383 41449
rect 9417 41415 9783 41449
rect 9817 41415 10183 41449
rect 10217 41415 10583 41449
rect 10617 41415 10983 41449
rect 11017 41415 11383 41449
rect 11417 41415 11783 41449
rect 11817 41415 12183 41449
rect 12217 41415 12583 41449
rect 12617 41415 12983 41449
rect 13017 41415 13383 41449
rect 13417 41415 13783 41449
rect 13817 41415 13968 41449
rect 6800 41402 13968 41415
rect 14932 41449 42638 41462
rect 14932 41415 15213 41449
rect 15247 41415 15613 41449
rect 15647 41415 16013 41449
rect 16047 41415 16413 41449
rect 16447 41415 16813 41449
rect 16847 41415 17213 41449
rect 17247 41415 17613 41449
rect 17647 41415 18013 41449
rect 18047 41415 18413 41449
rect 18447 41415 18813 41449
rect 18847 41415 19213 41449
rect 19247 41415 19613 41449
rect 19647 41415 20013 41449
rect 20047 41415 20413 41449
rect 20447 41415 20813 41449
rect 20847 41415 21213 41449
rect 21247 41415 21613 41449
rect 21647 41415 22013 41449
rect 22047 41415 22413 41449
rect 22447 41415 22813 41449
rect 22847 41415 23213 41449
rect 23247 41415 23613 41449
rect 23647 41415 24013 41449
rect 24047 41415 24413 41449
rect 24447 41415 24813 41449
rect 24847 41415 25213 41449
rect 25247 41415 25613 41449
rect 25647 41415 26013 41449
rect 26047 41415 26413 41449
rect 26447 41415 26813 41449
rect 26847 41415 27213 41449
rect 27247 41415 27613 41449
rect 27647 41415 28013 41449
rect 28047 41415 28413 41449
rect 28447 41415 28813 41449
rect 28847 41415 29213 41449
rect 29247 41415 29613 41449
rect 29647 41415 30013 41449
rect 30047 41415 30413 41449
rect 30447 41415 30813 41449
rect 30847 41415 31213 41449
rect 31247 41415 31613 41449
rect 31647 41415 32013 41449
rect 32047 41415 32413 41449
rect 32447 41415 32813 41449
rect 32847 41415 33213 41449
rect 33247 41415 33613 41449
rect 33647 41415 34013 41449
rect 34047 41415 34413 41449
rect 34447 41415 34813 41449
rect 34847 41415 35213 41449
rect 35247 41415 35613 41449
rect 35647 41415 36013 41449
rect 36047 41415 36413 41449
rect 36447 41415 36813 41449
rect 36847 41415 37213 41449
rect 37247 41415 37613 41449
rect 37647 41415 38013 41449
rect 38047 41415 38413 41449
rect 38447 41415 38813 41449
rect 38847 41415 39213 41449
rect 39247 41415 39613 41449
rect 39647 41415 40013 41449
rect 40047 41415 40413 41449
rect 40447 41415 40813 41449
rect 40847 41415 41213 41449
rect 41247 41415 41613 41449
rect 41647 41415 42013 41449
rect 42047 41415 42413 41449
rect 42447 41415 42638 41449
rect 14932 41402 42638 41415
rect 14960 41309 15020 41402
rect 16008 41359 16168 41402
rect 16008 41325 16073 41359
rect 16107 41325 16168 41359
rect 16008 41322 16168 41325
rect 17308 41359 17468 41402
rect 17308 41325 17373 41359
rect 17407 41325 17468 41359
rect 17308 41322 17468 41325
rect 18608 41359 18768 41402
rect 18608 41325 18673 41359
rect 18707 41325 18768 41359
rect 18608 41322 18768 41325
rect 19908 41359 20068 41402
rect 19908 41325 19973 41359
rect 20007 41325 20068 41359
rect 19908 41322 20068 41325
rect 21208 41359 21368 41402
rect 21208 41325 21273 41359
rect 21307 41325 21368 41359
rect 21208 41322 21368 41325
rect 22508 41359 22668 41402
rect 22508 41325 22573 41359
rect 22607 41325 22668 41359
rect 22508 41322 22668 41325
rect 23808 41359 23968 41402
rect 23808 41325 23873 41359
rect 23907 41325 23968 41359
rect 23808 41322 23968 41325
rect 25108 41359 25268 41402
rect 25108 41325 25173 41359
rect 25207 41325 25268 41359
rect 25108 41322 25268 41325
rect 26408 41359 26568 41402
rect 26408 41325 26473 41359
rect 26507 41325 26568 41359
rect 26408 41322 26568 41325
rect 27708 41359 27868 41402
rect 27708 41325 27773 41359
rect 27807 41325 27868 41359
rect 27708 41322 27868 41325
rect 29008 41359 29168 41402
rect 29008 41325 29073 41359
rect 29107 41325 29168 41359
rect 29008 41322 29168 41325
rect 30308 41359 30468 41402
rect 30308 41325 30373 41359
rect 30407 41325 30468 41359
rect 30308 41322 30468 41325
rect 31608 41359 31768 41402
rect 31608 41325 31673 41359
rect 31707 41325 31768 41359
rect 31608 41322 31768 41325
rect 32908 41359 33068 41402
rect 32908 41325 32973 41359
rect 33007 41325 33068 41359
rect 32908 41322 33068 41325
rect 34208 41359 34368 41402
rect 34208 41325 34273 41359
rect 34307 41325 34368 41359
rect 34208 41322 34368 41325
rect 35508 41359 35668 41402
rect 35508 41325 35573 41359
rect 35607 41325 35668 41359
rect 35508 41322 35668 41325
rect 36808 41359 36968 41402
rect 36808 41325 36873 41359
rect 36907 41325 36968 41359
rect 36808 41322 36968 41325
rect 38108 41359 38268 41402
rect 38108 41325 38173 41359
rect 38207 41325 38268 41359
rect 38108 41322 38268 41325
rect 39408 41359 39568 41402
rect 39408 41325 39473 41359
rect 39507 41325 39568 41359
rect 39408 41322 39568 41325
rect 40708 41359 40868 41402
rect 40708 41325 40773 41359
rect 40807 41325 40868 41359
rect 40708 41322 40868 41325
rect 5984 41242 6500 41302
rect 14960 41275 14973 41309
rect 15007 41275 15020 41309
rect 6453 40956 6487 41242
rect 14960 41192 15020 41275
rect 15090 41242 42638 41282
rect 15077 41181 15111 41201
rect 15077 41113 15111 41147
rect 15077 41045 15111 41075
rect 15077 40977 15111 41003
rect 5996 40929 6030 40956
rect 6453 40938 6488 40956
rect 5996 40857 6030 40875
rect 5996 40785 6030 40807
rect 5996 40713 6030 40739
rect 5996 40641 6030 40671
rect 5996 40569 6030 40603
rect 5996 40501 6030 40535
rect 5996 40433 6030 40463
rect 5996 40365 6030 40391
rect 5996 40297 6030 40319
rect 5996 40229 6030 40247
rect 5995 40175 5996 40206
rect 5995 40148 6030 40175
rect 6454 40929 6488 40938
rect 6454 40857 6488 40875
rect 6454 40785 6488 40807
rect 6454 40713 6488 40739
rect 6454 40641 6488 40671
rect 6454 40569 6488 40603
rect 6454 40501 6488 40535
rect 6454 40433 6488 40463
rect 6454 40365 6488 40391
rect 6454 40297 6488 40319
rect 6454 40229 6488 40247
rect 6454 40148 6488 40175
rect 15077 40909 15111 40931
rect 15077 40841 15111 40859
rect 15077 40773 15111 40787
rect 15077 40705 15111 40715
rect 15077 40637 15111 40643
rect 15077 40569 15111 40571
rect 15077 40533 15111 40535
rect 15077 40461 15111 40467
rect 15077 40389 15111 40399
rect 15077 40317 15111 40331
rect 15077 40245 15111 40263
rect 15077 40173 15111 40195
rect 5995 39982 6029 40148
rect 15077 40101 15111 40127
rect 15077 40029 15111 40059
rect 5984 39967 6500 39982
rect 5984 39933 6469 39967
rect 15077 39957 15111 39991
rect 5984 39922 6500 39933
rect 15077 39822 15111 39923
rect 15535 41181 15569 41242
rect 15535 41113 15569 41147
rect 15535 41045 15569 41075
rect 15535 40977 15569 41003
rect 15535 40909 15569 40931
rect 15535 40841 15569 40859
rect 15535 40773 15569 40787
rect 15535 40705 15569 40715
rect 15535 40637 15569 40643
rect 15535 40569 15569 40571
rect 15535 40533 15569 40535
rect 15535 40461 15569 40467
rect 15535 40389 15569 40399
rect 15535 40317 15569 40331
rect 15535 40245 15569 40263
rect 15535 40173 15569 40195
rect 15535 40101 15569 40127
rect 15535 40029 15569 40059
rect 15535 39957 15569 39991
rect 15535 39903 15569 39923
rect 15993 41181 16027 41201
rect 15993 41113 16027 41147
rect 15993 41045 16027 41075
rect 15993 40977 16027 41003
rect 15993 40909 16027 40931
rect 15993 40841 16027 40859
rect 15993 40773 16027 40787
rect 15993 40705 16027 40715
rect 15993 40637 16027 40643
rect 15993 40569 16027 40571
rect 15993 40533 16027 40535
rect 15993 40461 16027 40467
rect 15993 40389 16027 40399
rect 15993 40317 16027 40331
rect 15993 40245 16027 40263
rect 15993 40173 16027 40195
rect 15993 40101 16027 40127
rect 15993 40029 16027 40059
rect 15993 39957 16027 39991
rect 15993 39822 16027 39923
rect 16451 41181 16485 41242
rect 16451 41113 16485 41147
rect 16451 41045 16485 41075
rect 16451 40977 16485 41003
rect 16451 40909 16485 40931
rect 16451 40841 16485 40859
rect 16451 40773 16485 40787
rect 16451 40705 16485 40715
rect 16451 40637 16485 40643
rect 16451 40569 16485 40571
rect 16451 40533 16485 40535
rect 16451 40461 16485 40467
rect 16451 40389 16485 40399
rect 16451 40317 16485 40331
rect 16451 40245 16485 40263
rect 16451 40173 16485 40195
rect 16451 40101 16485 40127
rect 16451 40029 16485 40059
rect 16451 39957 16485 39991
rect 16451 39903 16485 39923
rect 16909 41181 16943 41201
rect 16909 41113 16943 41147
rect 16909 41045 16943 41075
rect 16909 40977 16943 41003
rect 16909 40909 16943 40931
rect 16909 40841 16943 40859
rect 16909 40773 16943 40787
rect 16909 40705 16943 40715
rect 16909 40637 16943 40643
rect 16909 40569 16943 40571
rect 16909 40533 16943 40535
rect 16909 40461 16943 40467
rect 16909 40389 16943 40399
rect 16909 40317 16943 40331
rect 16909 40245 16943 40263
rect 16909 40173 16943 40195
rect 16909 40101 16943 40127
rect 16909 40029 16943 40059
rect 16909 39957 16943 39991
rect 16909 39822 16943 39923
rect 17367 41181 17401 41242
rect 17367 41113 17401 41147
rect 17367 41045 17401 41075
rect 17367 40977 17401 41003
rect 17367 40909 17401 40931
rect 17367 40841 17401 40859
rect 17367 40773 17401 40787
rect 17367 40705 17401 40715
rect 17367 40637 17401 40643
rect 17367 40569 17401 40571
rect 17367 40533 17401 40535
rect 17367 40461 17401 40467
rect 17367 40389 17401 40399
rect 17367 40317 17401 40331
rect 17367 40245 17401 40263
rect 17367 40173 17401 40195
rect 17367 40101 17401 40127
rect 17367 40029 17401 40059
rect 17367 39957 17401 39991
rect 17367 39903 17401 39923
rect 17825 41181 17859 41201
rect 17825 41113 17859 41147
rect 17825 41045 17859 41075
rect 17825 40977 17859 41003
rect 17825 40909 17859 40931
rect 17825 40841 17859 40859
rect 17825 40773 17859 40787
rect 17825 40705 17859 40715
rect 17825 40637 17859 40643
rect 17825 40569 17859 40571
rect 17825 40533 17859 40535
rect 17825 40461 17859 40467
rect 17825 40389 17859 40399
rect 17825 40317 17859 40331
rect 17825 40245 17859 40263
rect 17825 40173 17859 40195
rect 17825 40101 17859 40127
rect 17825 40029 17859 40059
rect 17825 39957 17859 39991
rect 17825 39822 17859 39923
rect 18283 41181 18317 41242
rect 18283 41113 18317 41147
rect 18283 41045 18317 41075
rect 18283 40977 18317 41003
rect 18283 40909 18317 40931
rect 18283 40841 18317 40859
rect 18283 40773 18317 40787
rect 18283 40705 18317 40715
rect 18283 40637 18317 40643
rect 18283 40569 18317 40571
rect 18283 40533 18317 40535
rect 18283 40461 18317 40467
rect 18283 40389 18317 40399
rect 18283 40317 18317 40331
rect 18283 40245 18317 40263
rect 18283 40173 18317 40195
rect 18283 40101 18317 40127
rect 18283 40029 18317 40059
rect 18283 39957 18317 39991
rect 18283 39903 18317 39923
rect 18741 41181 18775 41201
rect 18741 41113 18775 41147
rect 18741 41045 18775 41075
rect 18741 40977 18775 41003
rect 18741 40909 18775 40931
rect 18741 40841 18775 40859
rect 18741 40773 18775 40787
rect 18741 40705 18775 40715
rect 18741 40637 18775 40643
rect 18741 40569 18775 40571
rect 18741 40533 18775 40535
rect 18741 40461 18775 40467
rect 18741 40389 18775 40399
rect 18741 40317 18775 40331
rect 18741 40245 18775 40263
rect 18741 40173 18775 40195
rect 18741 40101 18775 40127
rect 18741 40029 18775 40059
rect 18741 39957 18775 39991
rect 18741 39822 18775 39923
rect 19199 41181 19233 41242
rect 19199 41113 19233 41147
rect 19199 41045 19233 41075
rect 19199 40977 19233 41003
rect 19199 40909 19233 40931
rect 19199 40841 19233 40859
rect 19199 40773 19233 40787
rect 19199 40705 19233 40715
rect 19199 40637 19233 40643
rect 19199 40569 19233 40571
rect 19199 40533 19233 40535
rect 19199 40461 19233 40467
rect 19199 40389 19233 40399
rect 19199 40317 19233 40331
rect 19199 40245 19233 40263
rect 19199 40173 19233 40195
rect 19199 40101 19233 40127
rect 19199 40029 19233 40059
rect 19199 39957 19233 39991
rect 19199 39903 19233 39923
rect 19657 41181 19691 41201
rect 19657 41113 19691 41147
rect 19657 41045 19691 41075
rect 19657 40977 19691 41003
rect 19657 40909 19691 40931
rect 19657 40841 19691 40859
rect 19657 40773 19691 40787
rect 19657 40705 19691 40715
rect 19657 40637 19691 40643
rect 19657 40569 19691 40571
rect 19657 40533 19691 40535
rect 19657 40461 19691 40467
rect 19657 40389 19691 40399
rect 19657 40317 19691 40331
rect 19657 40245 19691 40263
rect 19657 40173 19691 40195
rect 19657 40101 19691 40127
rect 19657 40029 19691 40059
rect 19657 39957 19691 39991
rect 19657 39822 19691 39923
rect 20115 41181 20149 41242
rect 20115 41113 20149 41147
rect 20115 41045 20149 41075
rect 20115 40977 20149 41003
rect 20115 40909 20149 40931
rect 20115 40841 20149 40859
rect 20115 40773 20149 40787
rect 20115 40705 20149 40715
rect 20115 40637 20149 40643
rect 20115 40569 20149 40571
rect 20115 40533 20149 40535
rect 20115 40461 20149 40467
rect 20115 40389 20149 40399
rect 20115 40317 20149 40331
rect 20115 40245 20149 40263
rect 20115 40173 20149 40195
rect 20115 40101 20149 40127
rect 20115 40029 20149 40059
rect 20115 39957 20149 39991
rect 20115 39903 20149 39923
rect 20573 41181 20607 41201
rect 20573 41113 20607 41147
rect 20573 41045 20607 41075
rect 20573 40977 20607 41003
rect 20573 40909 20607 40931
rect 20573 40841 20607 40859
rect 20573 40773 20607 40787
rect 20573 40705 20607 40715
rect 20573 40637 20607 40643
rect 20573 40569 20607 40571
rect 20573 40533 20607 40535
rect 20573 40461 20607 40467
rect 20573 40389 20607 40399
rect 20573 40317 20607 40331
rect 20573 40245 20607 40263
rect 20573 40173 20607 40195
rect 20573 40101 20607 40127
rect 20573 40029 20607 40059
rect 20573 39957 20607 39991
rect 20573 39822 20607 39923
rect 21031 41181 21065 41242
rect 21031 41113 21065 41147
rect 21031 41045 21065 41075
rect 21031 40977 21065 41003
rect 21031 40909 21065 40931
rect 21031 40841 21065 40859
rect 21031 40773 21065 40787
rect 21031 40705 21065 40715
rect 21031 40637 21065 40643
rect 21031 40569 21065 40571
rect 21031 40533 21065 40535
rect 21031 40461 21065 40467
rect 21031 40389 21065 40399
rect 21031 40317 21065 40331
rect 21031 40245 21065 40263
rect 21031 40173 21065 40195
rect 21031 40101 21065 40127
rect 21031 40029 21065 40059
rect 21031 39957 21065 39991
rect 21031 39903 21065 39923
rect 21489 41181 21523 41201
rect 21489 41113 21523 41147
rect 21489 41045 21523 41075
rect 21489 40977 21523 41003
rect 21489 40909 21523 40931
rect 21489 40841 21523 40859
rect 21489 40773 21523 40787
rect 21489 40705 21523 40715
rect 21489 40637 21523 40643
rect 21489 40569 21523 40571
rect 21489 40533 21523 40535
rect 21489 40461 21523 40467
rect 21489 40389 21523 40399
rect 21489 40317 21523 40331
rect 21489 40245 21523 40263
rect 21489 40173 21523 40195
rect 21489 40101 21523 40127
rect 21489 40029 21523 40059
rect 21489 39957 21523 39991
rect 21489 39822 21523 39923
rect 21947 41181 21981 41242
rect 21947 41113 21981 41147
rect 21947 41045 21981 41075
rect 21947 40977 21981 41003
rect 21947 40909 21981 40931
rect 21947 40841 21981 40859
rect 21947 40773 21981 40787
rect 21947 40705 21981 40715
rect 21947 40637 21981 40643
rect 21947 40569 21981 40571
rect 21947 40533 21981 40535
rect 21947 40461 21981 40467
rect 21947 40389 21981 40399
rect 21947 40317 21981 40331
rect 21947 40245 21981 40263
rect 21947 40173 21981 40195
rect 21947 40101 21981 40127
rect 21947 40029 21981 40059
rect 21947 39957 21981 39991
rect 21947 39903 21981 39923
rect 22405 41181 22439 41201
rect 22405 41113 22439 41147
rect 22405 41045 22439 41075
rect 22405 40977 22439 41003
rect 22405 40909 22439 40931
rect 22405 40841 22439 40859
rect 22405 40773 22439 40787
rect 22405 40705 22439 40715
rect 22405 40637 22439 40643
rect 22405 40569 22439 40571
rect 22405 40533 22439 40535
rect 22405 40461 22439 40467
rect 22405 40389 22439 40399
rect 22405 40317 22439 40331
rect 22405 40245 22439 40263
rect 22405 40173 22439 40195
rect 22405 40101 22439 40127
rect 22405 40029 22439 40059
rect 22405 39957 22439 39991
rect 22405 39822 22439 39923
rect 22863 41181 22897 41242
rect 22863 41113 22897 41147
rect 22863 41045 22897 41075
rect 22863 40977 22897 41003
rect 22863 40909 22897 40931
rect 22863 40841 22897 40859
rect 22863 40773 22897 40787
rect 22863 40705 22897 40715
rect 22863 40637 22897 40643
rect 22863 40569 22897 40571
rect 22863 40533 22897 40535
rect 22863 40461 22897 40467
rect 22863 40389 22897 40399
rect 22863 40317 22897 40331
rect 22863 40245 22897 40263
rect 22863 40173 22897 40195
rect 22863 40101 22897 40127
rect 22863 40029 22897 40059
rect 22863 39957 22897 39991
rect 22863 39903 22897 39923
rect 23321 41181 23355 41201
rect 23321 41113 23355 41147
rect 23321 41045 23355 41075
rect 23321 40977 23355 41003
rect 23321 40909 23355 40931
rect 23321 40841 23355 40859
rect 23321 40773 23355 40787
rect 23321 40705 23355 40715
rect 23321 40637 23355 40643
rect 23321 40569 23355 40571
rect 23321 40533 23355 40535
rect 23321 40461 23355 40467
rect 23321 40389 23355 40399
rect 23321 40317 23355 40331
rect 23321 40245 23355 40263
rect 23321 40173 23355 40195
rect 23321 40101 23355 40127
rect 23321 40029 23355 40059
rect 23321 39957 23355 39991
rect 23321 39822 23355 39923
rect 23779 41181 23813 41242
rect 23779 41113 23813 41147
rect 23779 41045 23813 41075
rect 23779 40977 23813 41003
rect 23779 40909 23813 40931
rect 23779 40841 23813 40859
rect 23779 40773 23813 40787
rect 23779 40705 23813 40715
rect 23779 40637 23813 40643
rect 23779 40569 23813 40571
rect 23779 40533 23813 40535
rect 23779 40461 23813 40467
rect 23779 40389 23813 40399
rect 23779 40317 23813 40331
rect 23779 40245 23813 40263
rect 23779 40173 23813 40195
rect 23779 40101 23813 40127
rect 23779 40029 23813 40059
rect 23779 39957 23813 39991
rect 23779 39903 23813 39923
rect 24237 41181 24271 41201
rect 24237 41113 24271 41147
rect 24237 41045 24271 41075
rect 24237 40977 24271 41003
rect 24237 40909 24271 40931
rect 24237 40841 24271 40859
rect 24237 40773 24271 40787
rect 24237 40705 24271 40715
rect 24237 40637 24271 40643
rect 24237 40569 24271 40571
rect 24237 40533 24271 40535
rect 24237 40461 24271 40467
rect 24237 40389 24271 40399
rect 24237 40317 24271 40331
rect 24237 40245 24271 40263
rect 24237 40173 24271 40195
rect 24237 40101 24271 40127
rect 24237 40029 24271 40059
rect 24237 39957 24271 39991
rect 24237 39822 24271 39923
rect 24695 41181 24729 41242
rect 24695 41113 24729 41147
rect 24695 41045 24729 41075
rect 24695 40977 24729 41003
rect 24695 40909 24729 40931
rect 24695 40841 24729 40859
rect 24695 40773 24729 40787
rect 24695 40705 24729 40715
rect 24695 40637 24729 40643
rect 24695 40569 24729 40571
rect 24695 40533 24729 40535
rect 24695 40461 24729 40467
rect 24695 40389 24729 40399
rect 24695 40317 24729 40331
rect 24695 40245 24729 40263
rect 24695 40173 24729 40195
rect 24695 40101 24729 40127
rect 24695 40029 24729 40059
rect 24695 39957 24729 39991
rect 24695 39903 24729 39923
rect 25153 41181 25187 41201
rect 25153 41113 25187 41147
rect 25153 41045 25187 41075
rect 25153 40977 25187 41003
rect 25153 40909 25187 40931
rect 25153 40841 25187 40859
rect 25153 40773 25187 40787
rect 25153 40705 25187 40715
rect 25153 40637 25187 40643
rect 25153 40569 25187 40571
rect 25153 40533 25187 40535
rect 25153 40461 25187 40467
rect 25153 40389 25187 40399
rect 25153 40317 25187 40331
rect 25153 40245 25187 40263
rect 25153 40173 25187 40195
rect 25153 40101 25187 40127
rect 25153 40029 25187 40059
rect 25153 39957 25187 39991
rect 25153 39822 25187 39923
rect 25611 41181 25645 41242
rect 25611 41113 25645 41147
rect 25611 41045 25645 41075
rect 25611 40977 25645 41003
rect 25611 40909 25645 40931
rect 25611 40841 25645 40859
rect 25611 40773 25645 40787
rect 25611 40705 25645 40715
rect 25611 40637 25645 40643
rect 25611 40569 25645 40571
rect 25611 40533 25645 40535
rect 25611 40461 25645 40467
rect 25611 40389 25645 40399
rect 25611 40317 25645 40331
rect 25611 40245 25645 40263
rect 25611 40173 25645 40195
rect 25611 40101 25645 40127
rect 25611 40029 25645 40059
rect 25611 39957 25645 39991
rect 25611 39903 25645 39923
rect 26069 41181 26103 41201
rect 26069 41113 26103 41147
rect 26069 41045 26103 41075
rect 26069 40977 26103 41003
rect 26069 40909 26103 40931
rect 26069 40841 26103 40859
rect 26069 40773 26103 40787
rect 26069 40705 26103 40715
rect 26069 40637 26103 40643
rect 26069 40569 26103 40571
rect 26069 40533 26103 40535
rect 26069 40461 26103 40467
rect 26069 40389 26103 40399
rect 26069 40317 26103 40331
rect 26069 40245 26103 40263
rect 26069 40173 26103 40195
rect 26069 40101 26103 40127
rect 26069 40029 26103 40059
rect 26069 39957 26103 39991
rect 26069 39822 26103 39923
rect 26527 41181 26561 41242
rect 26527 41113 26561 41147
rect 26527 41045 26561 41075
rect 26527 40977 26561 41003
rect 26527 40909 26561 40931
rect 26527 40841 26561 40859
rect 26527 40773 26561 40787
rect 26527 40705 26561 40715
rect 26527 40637 26561 40643
rect 26527 40569 26561 40571
rect 26527 40533 26561 40535
rect 26527 40461 26561 40467
rect 26527 40389 26561 40399
rect 26527 40317 26561 40331
rect 26527 40245 26561 40263
rect 26527 40173 26561 40195
rect 26527 40101 26561 40127
rect 26527 40029 26561 40059
rect 26527 39957 26561 39991
rect 26527 39903 26561 39923
rect 26985 41181 27019 41201
rect 26985 41113 27019 41147
rect 26985 41045 27019 41075
rect 26985 40977 27019 41003
rect 26985 40909 27019 40931
rect 26985 40841 27019 40859
rect 26985 40773 27019 40787
rect 26985 40705 27019 40715
rect 26985 40637 27019 40643
rect 26985 40569 27019 40571
rect 26985 40533 27019 40535
rect 26985 40461 27019 40467
rect 26985 40389 27019 40399
rect 26985 40317 27019 40331
rect 26985 40245 27019 40263
rect 26985 40173 27019 40195
rect 26985 40101 27019 40127
rect 26985 40029 27019 40059
rect 26985 39957 27019 39991
rect 26985 39822 27019 39923
rect 27443 41181 27477 41242
rect 27443 41113 27477 41147
rect 27443 41045 27477 41075
rect 27443 40977 27477 41003
rect 27443 40909 27477 40931
rect 27443 40841 27477 40859
rect 27443 40773 27477 40787
rect 27443 40705 27477 40715
rect 27443 40637 27477 40643
rect 27443 40569 27477 40571
rect 27443 40533 27477 40535
rect 27443 40461 27477 40467
rect 27443 40389 27477 40399
rect 27443 40317 27477 40331
rect 27443 40245 27477 40263
rect 27443 40173 27477 40195
rect 27443 40101 27477 40127
rect 27443 40029 27477 40059
rect 27443 39957 27477 39991
rect 27443 39903 27477 39923
rect 27901 41181 27935 41201
rect 27901 41113 27935 41147
rect 27901 41045 27935 41075
rect 27901 40977 27935 41003
rect 27901 40909 27935 40931
rect 27901 40841 27935 40859
rect 27901 40773 27935 40787
rect 27901 40705 27935 40715
rect 27901 40637 27935 40643
rect 27901 40569 27935 40571
rect 27901 40533 27935 40535
rect 27901 40461 27935 40467
rect 27901 40389 27935 40399
rect 27901 40317 27935 40331
rect 27901 40245 27935 40263
rect 27901 40173 27935 40195
rect 27901 40101 27935 40127
rect 27901 40029 27935 40059
rect 27901 39957 27935 39991
rect 27901 39822 27935 39923
rect 28359 41181 28393 41242
rect 28359 41113 28393 41147
rect 28359 41045 28393 41075
rect 28359 40977 28393 41003
rect 28359 40909 28393 40931
rect 28359 40841 28393 40859
rect 28359 40773 28393 40787
rect 28359 40705 28393 40715
rect 28359 40637 28393 40643
rect 28359 40569 28393 40571
rect 28359 40533 28393 40535
rect 28359 40461 28393 40467
rect 28359 40389 28393 40399
rect 28359 40317 28393 40331
rect 28359 40245 28393 40263
rect 28359 40173 28393 40195
rect 28359 40101 28393 40127
rect 28359 40029 28393 40059
rect 28359 39957 28393 39991
rect 28359 39903 28393 39923
rect 28817 41181 28851 41201
rect 28817 41113 28851 41147
rect 28817 41045 28851 41075
rect 28817 40977 28851 41003
rect 28817 40909 28851 40931
rect 28817 40841 28851 40859
rect 28817 40773 28851 40787
rect 28817 40705 28851 40715
rect 28817 40637 28851 40643
rect 28817 40569 28851 40571
rect 28817 40533 28851 40535
rect 28817 40461 28851 40467
rect 28817 40389 28851 40399
rect 28817 40317 28851 40331
rect 28817 40245 28851 40263
rect 28817 40173 28851 40195
rect 28817 40101 28851 40127
rect 28817 40029 28851 40059
rect 28817 39957 28851 39991
rect 28817 39822 28851 39923
rect 29275 41181 29309 41242
rect 29275 41113 29309 41147
rect 29275 41045 29309 41075
rect 29275 40977 29309 41003
rect 29275 40909 29309 40931
rect 29275 40841 29309 40859
rect 29275 40773 29309 40787
rect 29275 40705 29309 40715
rect 29275 40637 29309 40643
rect 29275 40569 29309 40571
rect 29275 40533 29309 40535
rect 29275 40461 29309 40467
rect 29275 40389 29309 40399
rect 29275 40317 29309 40331
rect 29275 40245 29309 40263
rect 29275 40173 29309 40195
rect 29275 40101 29309 40127
rect 29275 40029 29309 40059
rect 29275 39957 29309 39991
rect 29275 39903 29309 39923
rect 29733 41181 29767 41201
rect 29733 41113 29767 41147
rect 29733 41045 29767 41075
rect 29733 40977 29767 41003
rect 29733 40909 29767 40931
rect 29733 40841 29767 40859
rect 29733 40773 29767 40787
rect 29733 40705 29767 40715
rect 29733 40637 29767 40643
rect 29733 40569 29767 40571
rect 29733 40533 29767 40535
rect 29733 40461 29767 40467
rect 29733 40389 29767 40399
rect 29733 40317 29767 40331
rect 29733 40245 29767 40263
rect 29733 40173 29767 40195
rect 29733 40101 29767 40127
rect 29733 40029 29767 40059
rect 29733 39957 29767 39991
rect 29733 39822 29767 39923
rect 30191 41181 30225 41242
rect 30191 41113 30225 41147
rect 30191 41045 30225 41075
rect 30191 40977 30225 41003
rect 30191 40909 30225 40931
rect 30191 40841 30225 40859
rect 30191 40773 30225 40787
rect 30191 40705 30225 40715
rect 30191 40637 30225 40643
rect 30191 40569 30225 40571
rect 30191 40533 30225 40535
rect 30191 40461 30225 40467
rect 30191 40389 30225 40399
rect 30191 40317 30225 40331
rect 30191 40245 30225 40263
rect 30191 40173 30225 40195
rect 30191 40101 30225 40127
rect 30191 40029 30225 40059
rect 30191 39957 30225 39991
rect 30191 39903 30225 39923
rect 30649 41181 30683 41201
rect 30649 41113 30683 41147
rect 30649 41045 30683 41075
rect 30649 40977 30683 41003
rect 30649 40909 30683 40931
rect 30649 40841 30683 40859
rect 30649 40773 30683 40787
rect 30649 40705 30683 40715
rect 30649 40637 30683 40643
rect 30649 40569 30683 40571
rect 30649 40533 30683 40535
rect 30649 40461 30683 40467
rect 30649 40389 30683 40399
rect 30649 40317 30683 40331
rect 30649 40245 30683 40263
rect 30649 40173 30683 40195
rect 30649 40101 30683 40127
rect 30649 40029 30683 40059
rect 30649 39957 30683 39991
rect 30649 39822 30683 39923
rect 31107 41181 31141 41242
rect 31107 41113 31141 41147
rect 31107 41045 31141 41075
rect 31107 40977 31141 41003
rect 31107 40909 31141 40931
rect 31107 40841 31141 40859
rect 31107 40773 31141 40787
rect 31107 40705 31141 40715
rect 31107 40637 31141 40643
rect 31107 40569 31141 40571
rect 31107 40533 31141 40535
rect 31107 40461 31141 40467
rect 31107 40389 31141 40399
rect 31107 40317 31141 40331
rect 31107 40245 31141 40263
rect 31107 40173 31141 40195
rect 31107 40101 31141 40127
rect 31107 40029 31141 40059
rect 31107 39957 31141 39991
rect 31107 39903 31141 39923
rect 31565 41181 31599 41201
rect 31565 41113 31599 41147
rect 31565 41045 31599 41075
rect 31565 40977 31599 41003
rect 31565 40909 31599 40931
rect 31565 40841 31599 40859
rect 31565 40773 31599 40787
rect 31565 40705 31599 40715
rect 31565 40637 31599 40643
rect 31565 40569 31599 40571
rect 31565 40533 31599 40535
rect 31565 40461 31599 40467
rect 31565 40389 31599 40399
rect 31565 40317 31599 40331
rect 31565 40245 31599 40263
rect 31565 40173 31599 40195
rect 31565 40101 31599 40127
rect 31565 40029 31599 40059
rect 31565 39957 31599 39991
rect 31565 39822 31599 39923
rect 32023 41181 32057 41242
rect 32023 41113 32057 41147
rect 32023 41045 32057 41075
rect 32023 40977 32057 41003
rect 32023 40909 32057 40931
rect 32023 40841 32057 40859
rect 32023 40773 32057 40787
rect 32023 40705 32057 40715
rect 32023 40637 32057 40643
rect 32023 40569 32057 40571
rect 32023 40533 32057 40535
rect 32023 40461 32057 40467
rect 32023 40389 32057 40399
rect 32023 40317 32057 40331
rect 32023 40245 32057 40263
rect 32023 40173 32057 40195
rect 32023 40101 32057 40127
rect 32023 40029 32057 40059
rect 32023 39957 32057 39991
rect 32023 39903 32057 39923
rect 32481 41181 32515 41201
rect 32481 41113 32515 41147
rect 32481 41045 32515 41075
rect 32481 40977 32515 41003
rect 32481 40909 32515 40931
rect 32481 40841 32515 40859
rect 32481 40773 32515 40787
rect 32481 40705 32515 40715
rect 32481 40637 32515 40643
rect 32481 40569 32515 40571
rect 32481 40533 32515 40535
rect 32481 40461 32515 40467
rect 32481 40389 32515 40399
rect 32481 40317 32515 40331
rect 32481 40245 32515 40263
rect 32481 40173 32515 40195
rect 32481 40101 32515 40127
rect 32481 40029 32515 40059
rect 32481 39957 32515 39991
rect 32481 39822 32515 39923
rect 32939 41181 32973 41242
rect 32939 41113 32973 41147
rect 32939 41045 32973 41075
rect 32939 40977 32973 41003
rect 32939 40909 32973 40931
rect 32939 40841 32973 40859
rect 32939 40773 32973 40787
rect 32939 40705 32973 40715
rect 32939 40637 32973 40643
rect 32939 40569 32973 40571
rect 32939 40533 32973 40535
rect 32939 40461 32973 40467
rect 32939 40389 32973 40399
rect 32939 40317 32973 40331
rect 32939 40245 32973 40263
rect 32939 40173 32973 40195
rect 32939 40101 32973 40127
rect 32939 40029 32973 40059
rect 32939 39957 32973 39991
rect 32939 39903 32973 39923
rect 33397 41181 33431 41201
rect 33397 41113 33431 41147
rect 33397 41045 33431 41075
rect 33397 40977 33431 41003
rect 33397 40909 33431 40931
rect 33397 40841 33431 40859
rect 33397 40773 33431 40787
rect 33397 40705 33431 40715
rect 33397 40637 33431 40643
rect 33397 40569 33431 40571
rect 33397 40533 33431 40535
rect 33397 40461 33431 40467
rect 33397 40389 33431 40399
rect 33397 40317 33431 40331
rect 33397 40245 33431 40263
rect 33397 40173 33431 40195
rect 33397 40101 33431 40127
rect 33397 40029 33431 40059
rect 33397 39957 33431 39991
rect 33397 39822 33431 39923
rect 33855 41181 33889 41242
rect 33855 41113 33889 41147
rect 33855 41045 33889 41075
rect 33855 40977 33889 41003
rect 33855 40909 33889 40931
rect 33855 40841 33889 40859
rect 33855 40773 33889 40787
rect 33855 40705 33889 40715
rect 33855 40637 33889 40643
rect 33855 40569 33889 40571
rect 33855 40533 33889 40535
rect 33855 40461 33889 40467
rect 33855 40389 33889 40399
rect 33855 40317 33889 40331
rect 33855 40245 33889 40263
rect 33855 40173 33889 40195
rect 33855 40101 33889 40127
rect 33855 40029 33889 40059
rect 33855 39957 33889 39991
rect 33855 39903 33889 39923
rect 34313 41181 34347 41201
rect 34313 41113 34347 41147
rect 34313 41045 34347 41075
rect 34313 40977 34347 41003
rect 34313 40909 34347 40931
rect 34313 40841 34347 40859
rect 34313 40773 34347 40787
rect 34313 40705 34347 40715
rect 34313 40637 34347 40643
rect 34313 40569 34347 40571
rect 34313 40533 34347 40535
rect 34313 40461 34347 40467
rect 34313 40389 34347 40399
rect 34313 40317 34347 40331
rect 34313 40245 34347 40263
rect 34313 40173 34347 40195
rect 34313 40101 34347 40127
rect 34313 40029 34347 40059
rect 34313 39957 34347 39991
rect 34313 39822 34347 39923
rect 34771 41181 34805 41242
rect 34771 41113 34805 41147
rect 34771 41045 34805 41075
rect 34771 40977 34805 41003
rect 34771 40909 34805 40931
rect 34771 40841 34805 40859
rect 34771 40773 34805 40787
rect 34771 40705 34805 40715
rect 34771 40637 34805 40643
rect 34771 40569 34805 40571
rect 34771 40533 34805 40535
rect 34771 40461 34805 40467
rect 34771 40389 34805 40399
rect 34771 40317 34805 40331
rect 34771 40245 34805 40263
rect 34771 40173 34805 40195
rect 34771 40101 34805 40127
rect 34771 40029 34805 40059
rect 34771 39957 34805 39991
rect 34771 39903 34805 39923
rect 35229 41181 35263 41201
rect 35229 41113 35263 41147
rect 35229 41045 35263 41075
rect 35229 40977 35263 41003
rect 35229 40909 35263 40931
rect 35229 40841 35263 40859
rect 35229 40773 35263 40787
rect 35229 40705 35263 40715
rect 35229 40637 35263 40643
rect 35229 40569 35263 40571
rect 35229 40533 35263 40535
rect 35229 40461 35263 40467
rect 35229 40389 35263 40399
rect 35229 40317 35263 40331
rect 35229 40245 35263 40263
rect 35229 40173 35263 40195
rect 35229 40101 35263 40127
rect 35229 40029 35263 40059
rect 35229 39957 35263 39991
rect 35229 39822 35263 39923
rect 35687 41181 35721 41242
rect 35687 41113 35721 41147
rect 35687 41045 35721 41075
rect 35687 40977 35721 41003
rect 35687 40909 35721 40931
rect 35687 40841 35721 40859
rect 35687 40773 35721 40787
rect 35687 40705 35721 40715
rect 35687 40637 35721 40643
rect 35687 40569 35721 40571
rect 35687 40533 35721 40535
rect 35687 40461 35721 40467
rect 35687 40389 35721 40399
rect 35687 40317 35721 40331
rect 35687 40245 35721 40263
rect 35687 40173 35721 40195
rect 35687 40101 35721 40127
rect 35687 40029 35721 40059
rect 35687 39957 35721 39991
rect 35687 39903 35721 39923
rect 36145 41181 36179 41201
rect 36145 41113 36179 41147
rect 36145 41045 36179 41075
rect 36145 40977 36179 41003
rect 36145 40909 36179 40931
rect 36145 40841 36179 40859
rect 36145 40773 36179 40787
rect 36145 40705 36179 40715
rect 36145 40637 36179 40643
rect 36145 40569 36179 40571
rect 36145 40533 36179 40535
rect 36145 40461 36179 40467
rect 36145 40389 36179 40399
rect 36145 40317 36179 40331
rect 36145 40245 36179 40263
rect 36145 40173 36179 40195
rect 36145 40101 36179 40127
rect 36145 40029 36179 40059
rect 36145 39957 36179 39991
rect 36145 39822 36179 39923
rect 36603 41181 36637 41242
rect 36603 41113 36637 41147
rect 36603 41045 36637 41075
rect 36603 40977 36637 41003
rect 36603 40909 36637 40931
rect 36603 40841 36637 40859
rect 36603 40773 36637 40787
rect 36603 40705 36637 40715
rect 36603 40637 36637 40643
rect 36603 40569 36637 40571
rect 36603 40533 36637 40535
rect 36603 40461 36637 40467
rect 36603 40389 36637 40399
rect 36603 40317 36637 40331
rect 36603 40245 36637 40263
rect 36603 40173 36637 40195
rect 36603 40101 36637 40127
rect 36603 40029 36637 40059
rect 36603 39957 36637 39991
rect 36603 39903 36637 39923
rect 37061 41181 37095 41201
rect 37061 41113 37095 41147
rect 37061 41045 37095 41075
rect 37061 40977 37095 41003
rect 37061 40909 37095 40931
rect 37061 40841 37095 40859
rect 37061 40773 37095 40787
rect 37061 40705 37095 40715
rect 37061 40637 37095 40643
rect 37061 40569 37095 40571
rect 37061 40533 37095 40535
rect 37061 40461 37095 40467
rect 37061 40389 37095 40399
rect 37061 40317 37095 40331
rect 37061 40245 37095 40263
rect 37061 40173 37095 40195
rect 37061 40101 37095 40127
rect 37061 40029 37095 40059
rect 37061 39957 37095 39991
rect 37061 39822 37095 39923
rect 37519 41181 37553 41242
rect 37519 41113 37553 41147
rect 37519 41045 37553 41075
rect 37519 40977 37553 41003
rect 37519 40909 37553 40931
rect 37519 40841 37553 40859
rect 37519 40773 37553 40787
rect 37519 40705 37553 40715
rect 37519 40637 37553 40643
rect 37519 40569 37553 40571
rect 37519 40533 37553 40535
rect 37519 40461 37553 40467
rect 37519 40389 37553 40399
rect 37519 40317 37553 40331
rect 37519 40245 37553 40263
rect 37519 40173 37553 40195
rect 37519 40101 37553 40127
rect 37519 40029 37553 40059
rect 37519 39957 37553 39991
rect 37519 39903 37553 39923
rect 37977 41181 38011 41201
rect 37977 41113 38011 41147
rect 37977 41045 38011 41075
rect 37977 40977 38011 41003
rect 37977 40909 38011 40931
rect 37977 40841 38011 40859
rect 37977 40773 38011 40787
rect 37977 40705 38011 40715
rect 37977 40637 38011 40643
rect 37977 40569 38011 40571
rect 37977 40533 38011 40535
rect 37977 40461 38011 40467
rect 37977 40389 38011 40399
rect 37977 40317 38011 40331
rect 37977 40245 38011 40263
rect 37977 40173 38011 40195
rect 37977 40101 38011 40127
rect 37977 40029 38011 40059
rect 37977 39957 38011 39991
rect 37977 39822 38011 39923
rect 38435 41181 38469 41242
rect 38435 41113 38469 41147
rect 38435 41045 38469 41075
rect 38435 40977 38469 41003
rect 38435 40909 38469 40931
rect 38435 40841 38469 40859
rect 38435 40773 38469 40787
rect 38435 40705 38469 40715
rect 38435 40637 38469 40643
rect 38435 40569 38469 40571
rect 38435 40533 38469 40535
rect 38435 40461 38469 40467
rect 38435 40389 38469 40399
rect 38435 40317 38469 40331
rect 38435 40245 38469 40263
rect 38435 40173 38469 40195
rect 38435 40101 38469 40127
rect 38435 40029 38469 40059
rect 38435 39957 38469 39991
rect 38435 39903 38469 39923
rect 38893 41181 38927 41201
rect 38893 41113 38927 41147
rect 38893 41045 38927 41075
rect 38893 40977 38927 41003
rect 38893 40909 38927 40931
rect 38893 40841 38927 40859
rect 38893 40773 38927 40787
rect 38893 40705 38927 40715
rect 38893 40637 38927 40643
rect 38893 40569 38927 40571
rect 38893 40533 38927 40535
rect 38893 40461 38927 40467
rect 38893 40389 38927 40399
rect 38893 40317 38927 40331
rect 38893 40245 38927 40263
rect 38893 40173 38927 40195
rect 38893 40101 38927 40127
rect 38893 40029 38927 40059
rect 38893 39957 38927 39991
rect 15030 39797 38669 39822
rect 38893 39822 38927 39923
rect 39351 41181 39385 41242
rect 39351 41113 39385 41147
rect 39351 41045 39385 41075
rect 39351 40977 39385 41003
rect 39351 40909 39385 40931
rect 39351 40841 39385 40859
rect 39351 40773 39385 40787
rect 39351 40705 39385 40715
rect 39351 40637 39385 40643
rect 39351 40569 39385 40571
rect 39351 40533 39385 40535
rect 39351 40461 39385 40467
rect 39351 40389 39385 40399
rect 39351 40317 39385 40331
rect 39351 40245 39385 40263
rect 39351 40173 39385 40195
rect 39351 40101 39385 40127
rect 39351 40029 39385 40059
rect 39351 39957 39385 39991
rect 39351 39903 39385 39923
rect 39809 41181 39843 41201
rect 39809 41113 39843 41147
rect 39809 41045 39843 41075
rect 39809 40977 39843 41003
rect 39809 40909 39843 40931
rect 39809 40841 39843 40859
rect 39809 40773 39843 40787
rect 39809 40705 39843 40715
rect 39809 40637 39843 40643
rect 39809 40569 39843 40571
rect 39809 40533 39843 40535
rect 39809 40461 39843 40467
rect 39809 40389 39843 40399
rect 39809 40317 39843 40331
rect 39809 40245 39843 40263
rect 39809 40173 39843 40195
rect 39809 40101 39843 40127
rect 39809 40029 39843 40059
rect 39809 39957 39843 39991
rect 39809 39822 39843 39923
rect 40267 41181 40301 41242
rect 40267 41113 40301 41147
rect 40267 41045 40301 41075
rect 40267 40977 40301 41003
rect 40267 40909 40301 40931
rect 40267 40841 40301 40859
rect 40267 40773 40301 40787
rect 40267 40705 40301 40715
rect 40267 40637 40301 40643
rect 40267 40569 40301 40571
rect 40267 40533 40301 40535
rect 40267 40461 40301 40467
rect 40267 40389 40301 40399
rect 40267 40317 40301 40331
rect 40267 40245 40301 40263
rect 40267 40173 40301 40195
rect 40267 40101 40301 40127
rect 40267 40029 40301 40059
rect 40267 39957 40301 39991
rect 40267 39903 40301 39923
rect 40725 41181 40759 41201
rect 40725 41113 40759 41147
rect 40725 41045 40759 41075
rect 40725 40977 40759 41003
rect 40725 40909 40759 40931
rect 40725 40841 40759 40859
rect 40725 40773 40759 40787
rect 40725 40705 40759 40715
rect 40725 40637 40759 40643
rect 40725 40569 40759 40571
rect 40725 40533 40759 40535
rect 40725 40461 40759 40467
rect 40725 40389 40759 40399
rect 40725 40317 40759 40331
rect 40725 40245 40759 40263
rect 40725 40173 40759 40195
rect 40725 40101 40759 40127
rect 40725 40029 40759 40059
rect 40725 39957 40759 39991
rect 40725 39822 40759 39923
rect 41183 41181 41217 41242
rect 41183 41113 41217 41147
rect 41183 41045 41217 41075
rect 41183 40977 41217 41003
rect 41183 40909 41217 40931
rect 41183 40841 41217 40859
rect 41183 40773 41217 40787
rect 41183 40705 41217 40715
rect 41183 40637 41217 40643
rect 41183 40569 41217 40571
rect 41183 40533 41217 40535
rect 41183 40461 41217 40467
rect 41183 40389 41217 40399
rect 41183 40317 41217 40331
rect 41183 40245 41217 40263
rect 41183 40173 41217 40195
rect 41183 40101 41217 40127
rect 41183 40029 41217 40059
rect 41183 39957 41217 39991
rect 41183 39903 41217 39923
rect 41641 41181 41675 41201
rect 41641 41113 41675 41147
rect 41641 41045 41675 41075
rect 41641 40977 41675 41003
rect 41641 40909 41675 40931
rect 41641 40841 41675 40859
rect 41641 40773 41675 40787
rect 41641 40705 41675 40715
rect 41641 40637 41675 40643
rect 41641 40569 41675 40571
rect 41641 40533 41675 40535
rect 41641 40461 41675 40467
rect 41641 40389 41675 40399
rect 41641 40317 41675 40331
rect 41641 40245 41675 40263
rect 41641 40173 41675 40195
rect 41641 40101 41675 40127
rect 41641 40029 41675 40059
rect 41641 39957 41675 39991
rect 41641 39822 41675 39923
rect 42099 41181 42133 41242
rect 42099 41113 42133 41147
rect 42099 41045 42133 41075
rect 42099 40977 42133 41003
rect 42099 40909 42133 40931
rect 42099 40841 42133 40859
rect 42099 40773 42133 40787
rect 42099 40705 42133 40715
rect 42099 40637 42133 40643
rect 42099 40569 42133 40571
rect 42099 40533 42133 40535
rect 42099 40461 42133 40467
rect 42099 40389 42133 40399
rect 42099 40317 42133 40331
rect 42099 40245 42133 40263
rect 42099 40173 42133 40195
rect 42099 40101 42133 40127
rect 42099 40029 42133 40059
rect 42099 39957 42133 39991
rect 42099 39903 42133 39923
rect 42557 41181 42591 41201
rect 42557 41113 42591 41147
rect 42557 41045 42591 41075
rect 42557 40977 42591 41003
rect 42557 40909 42591 40931
rect 42557 40841 42591 40859
rect 42557 40773 42591 40787
rect 42557 40705 42591 40715
rect 42557 40637 42591 40643
rect 42557 40569 42591 40571
rect 42557 40533 42591 40535
rect 42557 40461 42591 40467
rect 42557 40389 42591 40399
rect 42557 40317 42591 40331
rect 42557 40245 42591 40263
rect 42557 40173 42591 40195
rect 42557 40101 42591 40127
rect 42557 40029 42591 40059
rect 42557 39957 42591 39991
rect 42557 39822 42591 39923
rect 38703 39797 42638 39822
rect 5914 39709 5974 39792
rect 5914 39675 5927 39709
rect 5961 39675 5974 39709
rect 6064 39743 6469 39756
rect 6064 39709 6167 39743
rect 6201 39729 6469 39743
rect 15030 39762 42638 39797
rect 6201 39709 6500 39729
rect 6064 39696 6500 39709
rect 15030 39703 42638 39716
rect 15030 39695 15213 39703
rect 5914 39582 5974 39675
rect 15059 39669 15213 39695
rect 15247 39669 15613 39703
rect 15647 39669 16013 39703
rect 16047 39669 16413 39703
rect 16447 39669 16813 39703
rect 16847 39669 17213 39703
rect 17247 39669 17613 39703
rect 17647 39669 18013 39703
rect 18047 39669 18413 39703
rect 18447 39669 18813 39703
rect 18847 39669 19213 39703
rect 19247 39669 19613 39703
rect 19647 39669 20013 39703
rect 20047 39669 20413 39703
rect 20447 39669 20813 39703
rect 20847 39669 21213 39703
rect 21247 39669 21613 39703
rect 21647 39669 22013 39703
rect 22047 39669 22413 39703
rect 22447 39669 22813 39703
rect 22847 39669 23213 39703
rect 23247 39669 23613 39703
rect 23647 39669 24013 39703
rect 24047 39669 24413 39703
rect 24447 39669 24813 39703
rect 24847 39669 25213 39703
rect 25247 39669 25613 39703
rect 25647 39669 26013 39703
rect 26047 39669 26413 39703
rect 26447 39669 26813 39703
rect 26847 39669 27213 39703
rect 27247 39669 27613 39703
rect 27647 39695 28013 39703
rect 27663 39669 28013 39695
rect 28047 39669 28413 39703
rect 28447 39669 28813 39703
rect 28847 39669 29213 39703
rect 29247 39669 29613 39703
rect 29647 39669 30013 39703
rect 30047 39669 30413 39703
rect 30447 39669 30813 39703
rect 30847 39669 31213 39703
rect 31247 39669 31613 39703
rect 31647 39669 32013 39703
rect 32047 39669 32413 39703
rect 32447 39669 32813 39703
rect 32847 39669 33213 39703
rect 33247 39669 33613 39703
rect 33647 39669 34013 39703
rect 34047 39669 34413 39703
rect 34447 39669 34813 39703
rect 34847 39669 35213 39703
rect 35247 39669 35613 39703
rect 35647 39669 36013 39703
rect 36047 39669 36413 39703
rect 36447 39669 36813 39703
rect 36847 39669 37213 39703
rect 37247 39669 37613 39703
rect 37647 39669 38013 39703
rect 38047 39669 38413 39703
rect 38447 39669 38813 39703
rect 38847 39669 39213 39703
rect 39247 39669 39613 39703
rect 39647 39669 40013 39703
rect 40047 39669 40413 39703
rect 40447 39669 40813 39703
rect 40847 39669 41213 39703
rect 41247 39669 41613 39703
rect 41647 39669 42013 39703
rect 42047 39669 42413 39703
rect 42447 39669 42638 39703
rect 15059 39661 27629 39669
rect 27663 39661 42638 39669
rect 15030 39656 42638 39661
rect 5886 39569 6500 39582
rect 5886 39535 6167 39569
rect 6201 39535 6500 39569
rect 5886 39522 6500 39535
rect 6800 39569 13968 39582
rect 6800 39535 6983 39569
rect 7017 39535 7383 39569
rect 7417 39535 7783 39569
rect 7817 39535 8183 39569
rect 8217 39535 8583 39569
rect 8617 39535 8983 39569
rect 9017 39535 9383 39569
rect 9417 39535 9783 39569
rect 9817 39535 10183 39569
rect 10217 39535 10583 39569
rect 10617 39535 10983 39569
rect 11017 39535 11383 39569
rect 11417 39535 11783 39569
rect 11817 39535 12183 39569
rect 12217 39535 12583 39569
rect 12617 39535 12983 39569
rect 13017 39535 13383 39569
rect 13417 39535 13783 39569
rect 13817 39535 13968 39569
rect 6800 39522 13968 39535
rect 14932 39569 42638 39582
rect 14932 39535 15213 39569
rect 15247 39535 15613 39569
rect 15647 39535 16013 39569
rect 16047 39535 16413 39569
rect 16447 39535 16813 39569
rect 16847 39535 17213 39569
rect 17247 39535 17613 39569
rect 17647 39535 18013 39569
rect 18047 39535 18413 39569
rect 18447 39535 18813 39569
rect 18847 39535 19213 39569
rect 19247 39535 19613 39569
rect 19647 39535 20013 39569
rect 20047 39535 20413 39569
rect 20447 39535 20813 39569
rect 20847 39535 21213 39569
rect 21247 39535 21613 39569
rect 21647 39535 22013 39569
rect 22047 39535 22413 39569
rect 22447 39535 22813 39569
rect 22847 39535 23213 39569
rect 23247 39535 23613 39569
rect 23647 39535 24013 39569
rect 24047 39535 24413 39569
rect 24447 39535 24813 39569
rect 24847 39535 25213 39569
rect 25247 39535 25613 39569
rect 25647 39535 26013 39569
rect 26047 39535 26413 39569
rect 26447 39535 26813 39569
rect 26847 39535 27213 39569
rect 27247 39535 27613 39569
rect 27647 39535 28013 39569
rect 28047 39535 28413 39569
rect 28447 39535 28813 39569
rect 28847 39535 29213 39569
rect 29247 39535 29613 39569
rect 29647 39535 30013 39569
rect 30047 39535 30413 39569
rect 30447 39535 30813 39569
rect 30847 39535 31213 39569
rect 31247 39535 31613 39569
rect 31647 39535 32013 39569
rect 32047 39535 32413 39569
rect 32447 39535 32813 39569
rect 32847 39535 33213 39569
rect 33247 39535 33613 39569
rect 33647 39535 34013 39569
rect 34047 39535 34413 39569
rect 34447 39535 34813 39569
rect 34847 39535 35213 39569
rect 35247 39535 35613 39569
rect 35647 39535 36013 39569
rect 36047 39535 36413 39569
rect 36447 39535 36813 39569
rect 36847 39535 37213 39569
rect 37247 39535 37613 39569
rect 37647 39535 38013 39569
rect 38047 39535 38413 39569
rect 38447 39535 38813 39569
rect 38847 39535 39213 39569
rect 39247 39535 39613 39569
rect 39647 39535 40013 39569
rect 40047 39535 40413 39569
rect 40447 39535 40813 39569
rect 40847 39535 41213 39569
rect 41247 39535 41613 39569
rect 41647 39535 42013 39569
rect 42047 39535 42413 39569
rect 42447 39535 42638 39569
rect 14932 39522 42638 39535
rect 5918 37689 13086 37702
rect 5918 37655 6101 37689
rect 6135 37655 6501 37689
rect 6535 37655 6901 37689
rect 6935 37655 7301 37689
rect 7335 37655 7701 37689
rect 7735 37655 8101 37689
rect 8135 37655 8501 37689
rect 8535 37655 8901 37689
rect 8935 37655 9301 37689
rect 9335 37655 9701 37689
rect 9735 37655 10101 37689
rect 10135 37655 10501 37689
rect 10535 37655 10901 37689
rect 10935 37655 11301 37689
rect 11335 37655 11701 37689
rect 11735 37655 12101 37689
rect 12135 37655 12501 37689
rect 12535 37655 12901 37689
rect 12935 37655 13086 37689
rect 5918 37642 13086 37655
rect 13366 37689 20534 37702
rect 13366 37655 13549 37689
rect 13583 37655 13949 37689
rect 13983 37655 14349 37689
rect 14383 37655 14749 37689
rect 14783 37655 15149 37689
rect 15183 37655 15549 37689
rect 15583 37655 15949 37689
rect 15983 37655 16349 37689
rect 16383 37655 16749 37689
rect 16783 37655 17149 37689
rect 17183 37655 17549 37689
rect 17583 37655 17949 37689
rect 17983 37655 18349 37689
rect 18383 37655 18749 37689
rect 18783 37655 19149 37689
rect 19183 37655 19549 37689
rect 19583 37655 19949 37689
rect 19983 37655 20349 37689
rect 20383 37655 20534 37689
rect 13366 37642 20534 37655
rect 20814 37689 27982 37702
rect 20814 37655 20997 37689
rect 21031 37655 21397 37689
rect 21431 37655 21797 37689
rect 21831 37655 22197 37689
rect 22231 37655 22597 37689
rect 22631 37655 22997 37689
rect 23031 37655 23397 37689
rect 23431 37655 23797 37689
rect 23831 37655 24197 37689
rect 24231 37655 24597 37689
rect 24631 37655 24997 37689
rect 25031 37655 25397 37689
rect 25431 37655 25797 37689
rect 25831 37655 26197 37689
rect 26231 37655 26597 37689
rect 26631 37655 26997 37689
rect 27031 37655 27397 37689
rect 27431 37655 27797 37689
rect 27831 37655 27982 37689
rect 20814 37642 27982 37655
rect 28230 37689 28844 37702
rect 28230 37655 28511 37689
rect 28545 37655 28844 37689
rect 28230 37642 28844 37655
rect 30024 37689 39404 37702
rect 30024 37655 30207 37689
rect 30241 37655 30407 37689
rect 30441 37655 30607 37689
rect 30641 37655 30807 37689
rect 30841 37655 31007 37689
rect 31041 37655 31207 37689
rect 31241 37655 31407 37689
rect 31441 37655 31607 37689
rect 31641 37655 31807 37689
rect 31841 37655 32007 37689
rect 32041 37655 32207 37689
rect 32241 37655 32407 37689
rect 32441 37655 32607 37689
rect 32641 37655 32807 37689
rect 32841 37655 33007 37689
rect 33041 37655 33207 37689
rect 33241 37655 33407 37689
rect 33441 37655 33607 37689
rect 33641 37655 33807 37689
rect 33841 37655 34007 37689
rect 34041 37655 34207 37689
rect 34241 37655 34407 37689
rect 34441 37655 34607 37689
rect 34641 37655 34807 37689
rect 34841 37655 35007 37689
rect 35041 37655 35207 37689
rect 35241 37655 35407 37689
rect 35441 37655 35607 37689
rect 35641 37655 35807 37689
rect 35841 37655 36007 37689
rect 36041 37655 36207 37689
rect 36241 37655 36407 37689
rect 36441 37655 36607 37689
rect 36641 37655 36807 37689
rect 36841 37655 37007 37689
rect 37041 37655 37207 37689
rect 37241 37655 37407 37689
rect 37441 37655 37607 37689
rect 37641 37655 37807 37689
rect 37841 37655 38007 37689
rect 38041 37655 38207 37689
rect 38241 37655 38407 37689
rect 38441 37655 38607 37689
rect 38641 37655 38807 37689
rect 38841 37655 39007 37689
rect 39041 37655 39207 37689
rect 39241 37655 39404 37689
rect 30024 37642 39404 37655
rect 39746 37689 42186 37702
rect 39746 37655 39929 37689
rect 39963 37655 40129 37689
rect 40163 37655 40329 37689
rect 40363 37655 40529 37689
rect 40563 37655 40729 37689
rect 40763 37655 40929 37689
rect 40963 37655 41129 37689
rect 41163 37655 41329 37689
rect 41363 37655 41529 37689
rect 41563 37655 41729 37689
rect 41763 37655 41929 37689
rect 41963 37655 42186 37689
rect 39746 37642 42186 37655
rect 28328 37519 28844 37542
rect 28328 37485 28825 37519
rect 28328 37482 28844 37485
rect 28797 37196 28831 37482
rect 30050 37356 39378 37376
rect 30050 37322 30070 37356
rect 30104 37322 30160 37356
rect 30194 37341 30250 37356
rect 30284 37341 30340 37356
rect 30374 37341 30430 37356
rect 30464 37341 30520 37356
rect 30554 37341 30610 37356
rect 30644 37341 30700 37356
rect 30734 37341 30790 37356
rect 30824 37341 30880 37356
rect 30914 37341 30970 37356
rect 31004 37341 31060 37356
rect 31094 37341 31150 37356
rect 31184 37341 31240 37356
rect 30214 37322 30250 37341
rect 30304 37322 30340 37341
rect 30394 37322 30430 37341
rect 30484 37322 30520 37341
rect 30574 37322 30610 37341
rect 30664 37322 30700 37341
rect 30754 37322 30790 37341
rect 30844 37322 30880 37341
rect 30934 37322 30970 37341
rect 31024 37322 31060 37341
rect 31114 37322 31150 37341
rect 31204 37322 31240 37341
rect 31274 37322 31410 37356
rect 31444 37322 31500 37356
rect 31534 37341 31590 37356
rect 31624 37341 31680 37356
rect 31714 37341 31770 37356
rect 31804 37341 31860 37356
rect 31894 37341 31950 37356
rect 31984 37341 32040 37356
rect 32074 37341 32130 37356
rect 32164 37341 32220 37356
rect 32254 37341 32310 37356
rect 32344 37341 32400 37356
rect 32434 37341 32490 37356
rect 32524 37341 32580 37356
rect 31554 37322 31590 37341
rect 31644 37322 31680 37341
rect 31734 37322 31770 37341
rect 31824 37322 31860 37341
rect 31914 37322 31950 37341
rect 32004 37322 32040 37341
rect 32094 37322 32130 37341
rect 32184 37322 32220 37341
rect 32274 37322 32310 37341
rect 32364 37322 32400 37341
rect 32454 37322 32490 37341
rect 32544 37322 32580 37341
rect 32614 37322 32750 37356
rect 32784 37322 32840 37356
rect 32874 37341 32930 37356
rect 32964 37341 33020 37356
rect 33054 37341 33110 37356
rect 33144 37341 33200 37356
rect 33234 37341 33290 37356
rect 33324 37341 33380 37356
rect 33414 37341 33470 37356
rect 33504 37341 33560 37356
rect 33594 37341 33650 37356
rect 33684 37341 33740 37356
rect 33774 37341 33830 37356
rect 33864 37341 33920 37356
rect 32894 37322 32930 37341
rect 32984 37322 33020 37341
rect 33074 37322 33110 37341
rect 33164 37322 33200 37341
rect 33254 37322 33290 37341
rect 33344 37322 33380 37341
rect 33434 37322 33470 37341
rect 33524 37322 33560 37341
rect 33614 37322 33650 37341
rect 33704 37322 33740 37341
rect 33794 37322 33830 37341
rect 33884 37322 33920 37341
rect 33954 37322 34090 37356
rect 34124 37322 34180 37356
rect 34214 37341 34270 37356
rect 34304 37341 34360 37356
rect 34394 37341 34450 37356
rect 34484 37341 34540 37356
rect 34574 37341 34630 37356
rect 34664 37341 34720 37356
rect 34754 37341 34810 37356
rect 34844 37341 34900 37356
rect 34934 37341 34990 37356
rect 35024 37341 35080 37356
rect 35114 37341 35170 37356
rect 35204 37341 35260 37356
rect 34234 37322 34270 37341
rect 34324 37322 34360 37341
rect 34414 37322 34450 37341
rect 34504 37322 34540 37341
rect 34594 37322 34630 37341
rect 34684 37322 34720 37341
rect 34774 37322 34810 37341
rect 34864 37322 34900 37341
rect 34954 37322 34990 37341
rect 35044 37322 35080 37341
rect 35134 37322 35170 37341
rect 35224 37322 35260 37341
rect 35294 37322 35430 37356
rect 35464 37322 35520 37356
rect 35554 37341 35610 37356
rect 35644 37341 35700 37356
rect 35734 37341 35790 37356
rect 35824 37341 35880 37356
rect 35914 37341 35970 37356
rect 36004 37341 36060 37356
rect 36094 37341 36150 37356
rect 36184 37341 36240 37356
rect 36274 37341 36330 37356
rect 36364 37341 36420 37356
rect 36454 37341 36510 37356
rect 36544 37341 36600 37356
rect 35574 37322 35610 37341
rect 35664 37322 35700 37341
rect 35754 37322 35790 37341
rect 35844 37322 35880 37341
rect 35934 37322 35970 37341
rect 36024 37322 36060 37341
rect 36114 37322 36150 37341
rect 36204 37322 36240 37341
rect 36294 37322 36330 37341
rect 36384 37322 36420 37341
rect 36474 37322 36510 37341
rect 36564 37322 36600 37341
rect 36634 37322 36770 37356
rect 36804 37322 36860 37356
rect 36894 37341 36950 37356
rect 36984 37341 37040 37356
rect 37074 37341 37130 37356
rect 37164 37341 37220 37356
rect 37254 37341 37310 37356
rect 37344 37341 37400 37356
rect 37434 37341 37490 37356
rect 37524 37341 37580 37356
rect 37614 37341 37670 37356
rect 37704 37341 37760 37356
rect 37794 37341 37850 37356
rect 37884 37341 37940 37356
rect 36914 37322 36950 37341
rect 37004 37322 37040 37341
rect 37094 37322 37130 37341
rect 37184 37322 37220 37341
rect 37274 37322 37310 37341
rect 37364 37322 37400 37341
rect 37454 37322 37490 37341
rect 37544 37322 37580 37341
rect 37634 37322 37670 37341
rect 37724 37322 37760 37341
rect 37814 37322 37850 37341
rect 37904 37322 37940 37341
rect 37974 37322 38110 37356
rect 38144 37322 38200 37356
rect 38234 37341 38290 37356
rect 38324 37341 38380 37356
rect 38414 37341 38470 37356
rect 38504 37341 38560 37356
rect 38594 37341 38650 37356
rect 38684 37341 38740 37356
rect 38774 37341 38830 37356
rect 38864 37341 38920 37356
rect 38954 37341 39010 37356
rect 39044 37341 39100 37356
rect 39134 37341 39190 37356
rect 39224 37341 39280 37356
rect 38254 37322 38290 37341
rect 38344 37322 38380 37341
rect 38434 37322 38470 37341
rect 38524 37322 38560 37341
rect 38614 37322 38650 37341
rect 38704 37322 38740 37341
rect 38794 37322 38830 37341
rect 38884 37322 38920 37341
rect 38974 37322 39010 37341
rect 39064 37322 39100 37341
rect 39154 37322 39190 37341
rect 39244 37322 39280 37341
rect 39314 37322 39378 37356
rect 30050 37318 30180 37322
rect 30050 37284 30084 37318
rect 30118 37307 30180 37318
rect 30214 37307 30270 37322
rect 30304 37307 30360 37322
rect 30394 37307 30450 37322
rect 30484 37307 30540 37322
rect 30574 37307 30630 37322
rect 30664 37307 30720 37322
rect 30754 37307 30810 37322
rect 30844 37307 30900 37322
rect 30934 37307 30990 37322
rect 31024 37307 31080 37322
rect 31114 37307 31170 37322
rect 31204 37318 31520 37322
rect 31204 37307 31271 37318
rect 30118 37284 31271 37307
rect 31305 37284 31424 37318
rect 31458 37307 31520 37318
rect 31554 37307 31610 37322
rect 31644 37307 31700 37322
rect 31734 37307 31790 37322
rect 31824 37307 31880 37322
rect 31914 37307 31970 37322
rect 32004 37307 32060 37322
rect 32094 37307 32150 37322
rect 32184 37307 32240 37322
rect 32274 37307 32330 37322
rect 32364 37307 32420 37322
rect 32454 37307 32510 37322
rect 32544 37318 32860 37322
rect 32544 37307 32611 37318
rect 31458 37284 32611 37307
rect 32645 37284 32764 37318
rect 32798 37307 32860 37318
rect 32894 37307 32950 37322
rect 32984 37307 33040 37322
rect 33074 37307 33130 37322
rect 33164 37307 33220 37322
rect 33254 37307 33310 37322
rect 33344 37307 33400 37322
rect 33434 37307 33490 37322
rect 33524 37307 33580 37322
rect 33614 37307 33670 37322
rect 33704 37307 33760 37322
rect 33794 37307 33850 37322
rect 33884 37318 34200 37322
rect 33884 37307 33951 37318
rect 32798 37284 33951 37307
rect 33985 37284 34104 37318
rect 34138 37307 34200 37318
rect 34234 37307 34290 37322
rect 34324 37307 34380 37322
rect 34414 37307 34470 37322
rect 34504 37307 34560 37322
rect 34594 37307 34650 37322
rect 34684 37307 34740 37322
rect 34774 37307 34830 37322
rect 34864 37307 34920 37322
rect 34954 37307 35010 37322
rect 35044 37307 35100 37322
rect 35134 37307 35190 37322
rect 35224 37318 35540 37322
rect 35224 37307 35291 37318
rect 34138 37284 35291 37307
rect 35325 37284 35444 37318
rect 35478 37307 35540 37318
rect 35574 37307 35630 37322
rect 35664 37307 35720 37322
rect 35754 37307 35810 37322
rect 35844 37307 35900 37322
rect 35934 37307 35990 37322
rect 36024 37307 36080 37322
rect 36114 37307 36170 37322
rect 36204 37307 36260 37322
rect 36294 37307 36350 37322
rect 36384 37307 36440 37322
rect 36474 37307 36530 37322
rect 36564 37318 36880 37322
rect 36564 37307 36631 37318
rect 35478 37284 36631 37307
rect 36665 37284 36784 37318
rect 36818 37307 36880 37318
rect 36914 37307 36970 37322
rect 37004 37307 37060 37322
rect 37094 37307 37150 37322
rect 37184 37307 37240 37322
rect 37274 37307 37330 37322
rect 37364 37307 37420 37322
rect 37454 37307 37510 37322
rect 37544 37307 37600 37322
rect 37634 37307 37690 37322
rect 37724 37307 37780 37322
rect 37814 37307 37870 37322
rect 37904 37318 38220 37322
rect 37904 37307 37971 37318
rect 36818 37284 37971 37307
rect 38005 37284 38124 37318
rect 38158 37307 38220 37318
rect 38254 37307 38310 37322
rect 38344 37307 38400 37322
rect 38434 37307 38490 37322
rect 38524 37307 38580 37322
rect 38614 37307 38670 37322
rect 38704 37307 38760 37322
rect 38794 37307 38850 37322
rect 38884 37307 38940 37322
rect 38974 37307 39030 37322
rect 39064 37307 39120 37322
rect 39154 37307 39210 37322
rect 39244 37318 39378 37322
rect 39244 37307 39311 37318
rect 38158 37284 39311 37307
rect 39345 37284 39378 37318
rect 30050 37277 39378 37284
rect 30050 37228 30149 37277
rect 28340 37169 28374 37196
rect 28797 37178 28832 37196
rect 28340 37097 28374 37115
rect 28340 37025 28374 37047
rect 28340 36953 28374 36979
rect 28340 36881 28374 36911
rect 28340 36809 28374 36843
rect 28340 36741 28374 36775
rect 28340 36673 28374 36703
rect 28340 36605 28374 36631
rect 28340 36537 28374 36559
rect 28340 36469 28374 36487
rect 28339 36415 28340 36446
rect 28339 36388 28374 36415
rect 28798 37169 28832 37178
rect 28798 37097 28832 37115
rect 28798 37025 28832 37047
rect 28798 36953 28832 36979
rect 28798 36881 28832 36911
rect 28798 36809 28832 36843
rect 28798 36741 28832 36775
rect 28798 36673 28832 36703
rect 28798 36605 28832 36631
rect 28798 36537 28832 36559
rect 28798 36469 28832 36487
rect 28798 36388 28832 36415
rect 30050 37194 30084 37228
rect 30118 37194 30149 37228
rect 31239 37228 31489 37277
rect 30050 37138 30149 37194
rect 30050 37104 30084 37138
rect 30118 37104 30149 37138
rect 30050 37048 30149 37104
rect 30050 37014 30084 37048
rect 30118 37014 30149 37048
rect 30050 36958 30149 37014
rect 30050 36924 30084 36958
rect 30118 36924 30149 36958
rect 30050 36868 30149 36924
rect 30050 36834 30084 36868
rect 30118 36834 30149 36868
rect 30050 36778 30149 36834
rect 30050 36744 30084 36778
rect 30118 36744 30149 36778
rect 30050 36688 30149 36744
rect 30050 36654 30084 36688
rect 30118 36654 30149 36688
rect 30050 36598 30149 36654
rect 30050 36564 30084 36598
rect 30118 36564 30149 36598
rect 30050 36508 30149 36564
rect 30050 36474 30084 36508
rect 30118 36474 30149 36508
rect 30050 36418 30149 36474
rect 28339 36227 28373 36388
rect 30050 36384 30084 36418
rect 30118 36384 30149 36418
rect 30050 36328 30149 36384
rect 30050 36294 30084 36328
rect 30118 36294 30149 36328
rect 30050 36238 30149 36294
rect 30213 37196 31175 37213
rect 30213 37162 30234 37196
rect 30268 37162 30324 37196
rect 30358 37194 30414 37196
rect 30448 37194 30504 37196
rect 30538 37194 30594 37196
rect 30628 37194 30684 37196
rect 30718 37194 30774 37196
rect 30808 37194 30864 37196
rect 30898 37194 30954 37196
rect 30988 37194 31044 37196
rect 31078 37194 31134 37196
rect 30378 37162 30414 37194
rect 30468 37162 30504 37194
rect 30558 37162 30594 37194
rect 30648 37162 30684 37194
rect 30738 37162 30774 37194
rect 30828 37162 30864 37194
rect 30918 37162 30954 37194
rect 31008 37162 31044 37194
rect 31098 37162 31134 37194
rect 31168 37162 31175 37196
rect 30213 37160 30344 37162
rect 30378 37160 30434 37162
rect 30468 37160 30524 37162
rect 30558 37160 30614 37162
rect 30648 37160 30704 37162
rect 30738 37160 30794 37162
rect 30828 37160 30884 37162
rect 30918 37160 30974 37162
rect 31008 37160 31064 37162
rect 31098 37160 31175 37162
rect 30213 37141 31175 37160
rect 30213 37137 30285 37141
rect 30213 37103 30232 37137
rect 30266 37103 30285 37137
rect 30213 37047 30285 37103
rect 31103 37118 31175 37141
rect 31103 37084 31122 37118
rect 31156 37084 31175 37118
rect 30213 37013 30232 37047
rect 30266 37013 30285 37047
rect 30213 36957 30285 37013
rect 30213 36923 30232 36957
rect 30266 36923 30285 36957
rect 30213 36867 30285 36923
rect 30213 36833 30232 36867
rect 30266 36833 30285 36867
rect 30213 36777 30285 36833
rect 30213 36743 30232 36777
rect 30266 36743 30285 36777
rect 30213 36687 30285 36743
rect 30213 36653 30232 36687
rect 30266 36653 30285 36687
rect 30213 36597 30285 36653
rect 30213 36563 30232 36597
rect 30266 36563 30285 36597
rect 30213 36507 30285 36563
rect 30213 36473 30232 36507
rect 30266 36473 30285 36507
rect 30213 36417 30285 36473
rect 30213 36383 30232 36417
rect 30266 36383 30285 36417
rect 30347 37020 31041 37079
rect 30347 36986 30408 37020
rect 30442 36992 30498 37020
rect 30532 36992 30588 37020
rect 30622 36992 30678 37020
rect 30454 36986 30498 36992
rect 30554 36986 30588 36992
rect 30654 36986 30678 36992
rect 30712 36992 30768 37020
rect 30712 36986 30720 36992
rect 30347 36958 30420 36986
rect 30454 36958 30520 36986
rect 30554 36958 30620 36986
rect 30654 36958 30720 36986
rect 30754 36986 30768 36992
rect 30802 36992 30858 37020
rect 30802 36986 30820 36992
rect 30754 36958 30820 36986
rect 30854 36986 30858 36992
rect 30892 36992 30948 37020
rect 30892 36986 30920 36992
rect 30982 36986 31041 37020
rect 30854 36958 30920 36986
rect 30954 36958 31041 36986
rect 30347 36930 31041 36958
rect 30347 36896 30408 36930
rect 30442 36896 30498 36930
rect 30532 36896 30588 36930
rect 30622 36896 30678 36930
rect 30712 36896 30768 36930
rect 30802 36896 30858 36930
rect 30892 36896 30948 36930
rect 30982 36896 31041 36930
rect 30347 36892 31041 36896
rect 30347 36858 30420 36892
rect 30454 36858 30520 36892
rect 30554 36858 30620 36892
rect 30654 36858 30720 36892
rect 30754 36858 30820 36892
rect 30854 36858 30920 36892
rect 30954 36858 31041 36892
rect 30347 36840 31041 36858
rect 30347 36806 30408 36840
rect 30442 36806 30498 36840
rect 30532 36806 30588 36840
rect 30622 36806 30678 36840
rect 30712 36806 30768 36840
rect 30802 36806 30858 36840
rect 30892 36806 30948 36840
rect 30982 36806 31041 36840
rect 30347 36792 31041 36806
rect 30347 36758 30420 36792
rect 30454 36758 30520 36792
rect 30554 36758 30620 36792
rect 30654 36758 30720 36792
rect 30754 36758 30820 36792
rect 30854 36758 30920 36792
rect 30954 36758 31041 36792
rect 30347 36750 31041 36758
rect 30347 36716 30408 36750
rect 30442 36716 30498 36750
rect 30532 36716 30588 36750
rect 30622 36716 30678 36750
rect 30712 36716 30768 36750
rect 30802 36716 30858 36750
rect 30892 36716 30948 36750
rect 30982 36716 31041 36750
rect 30347 36692 31041 36716
rect 30347 36660 30420 36692
rect 30454 36660 30520 36692
rect 30554 36660 30620 36692
rect 30654 36660 30720 36692
rect 30347 36626 30408 36660
rect 30454 36658 30498 36660
rect 30554 36658 30588 36660
rect 30654 36658 30678 36660
rect 30442 36626 30498 36658
rect 30532 36626 30588 36658
rect 30622 36626 30678 36658
rect 30712 36658 30720 36660
rect 30754 36660 30820 36692
rect 30754 36658 30768 36660
rect 30712 36626 30768 36658
rect 30802 36658 30820 36660
rect 30854 36660 30920 36692
rect 30954 36660 31041 36692
rect 30854 36658 30858 36660
rect 30802 36626 30858 36658
rect 30892 36658 30920 36660
rect 30892 36626 30948 36658
rect 30982 36626 31041 36660
rect 30347 36592 31041 36626
rect 30347 36570 30420 36592
rect 30454 36570 30520 36592
rect 30554 36570 30620 36592
rect 30654 36570 30720 36592
rect 30347 36536 30408 36570
rect 30454 36558 30498 36570
rect 30554 36558 30588 36570
rect 30654 36558 30678 36570
rect 30442 36536 30498 36558
rect 30532 36536 30588 36558
rect 30622 36536 30678 36558
rect 30712 36558 30720 36570
rect 30754 36570 30820 36592
rect 30754 36558 30768 36570
rect 30712 36536 30768 36558
rect 30802 36558 30820 36570
rect 30854 36570 30920 36592
rect 30954 36570 31041 36592
rect 30854 36558 30858 36570
rect 30802 36536 30858 36558
rect 30892 36558 30920 36570
rect 30892 36536 30948 36558
rect 30982 36536 31041 36570
rect 30347 36492 31041 36536
rect 30347 36480 30420 36492
rect 30454 36480 30520 36492
rect 30554 36480 30620 36492
rect 30654 36480 30720 36492
rect 30347 36446 30408 36480
rect 30454 36458 30498 36480
rect 30554 36458 30588 36480
rect 30654 36458 30678 36480
rect 30442 36446 30498 36458
rect 30532 36446 30588 36458
rect 30622 36446 30678 36458
rect 30712 36458 30720 36480
rect 30754 36480 30820 36492
rect 30754 36458 30768 36480
rect 30712 36446 30768 36458
rect 30802 36458 30820 36480
rect 30854 36480 30920 36492
rect 30954 36480 31041 36492
rect 30854 36458 30858 36480
rect 30802 36446 30858 36458
rect 30892 36458 30920 36480
rect 30892 36446 30948 36458
rect 30982 36446 31041 36480
rect 30347 36385 31041 36446
rect 31103 37028 31175 37084
rect 31103 36994 31122 37028
rect 31156 36994 31175 37028
rect 31103 36938 31175 36994
rect 31103 36904 31122 36938
rect 31156 36904 31175 36938
rect 31103 36848 31175 36904
rect 31103 36814 31122 36848
rect 31156 36814 31175 36848
rect 31103 36758 31175 36814
rect 31103 36724 31122 36758
rect 31156 36724 31175 36758
rect 31103 36668 31175 36724
rect 31103 36634 31122 36668
rect 31156 36634 31175 36668
rect 31103 36578 31175 36634
rect 31103 36544 31122 36578
rect 31156 36544 31175 36578
rect 31103 36488 31175 36544
rect 31103 36454 31122 36488
rect 31156 36454 31175 36488
rect 31103 36398 31175 36454
rect 30213 36323 30285 36383
rect 31103 36364 31122 36398
rect 31156 36364 31175 36398
rect 31103 36323 31175 36364
rect 30213 36304 31175 36323
rect 30213 36270 30310 36304
rect 30344 36270 30400 36304
rect 30434 36270 30490 36304
rect 30524 36270 30580 36304
rect 30614 36270 30670 36304
rect 30704 36270 30760 36304
rect 30794 36270 30850 36304
rect 30884 36270 30940 36304
rect 30974 36270 31030 36304
rect 31064 36270 31175 36304
rect 30213 36251 31175 36270
rect 31239 37194 31271 37228
rect 31305 37194 31424 37228
rect 31458 37194 31489 37228
rect 32579 37228 32829 37277
rect 31239 37138 31489 37194
rect 31239 37104 31271 37138
rect 31305 37104 31424 37138
rect 31458 37104 31489 37138
rect 31239 37048 31489 37104
rect 31239 37014 31271 37048
rect 31305 37014 31424 37048
rect 31458 37014 31489 37048
rect 31239 36958 31489 37014
rect 31239 36924 31271 36958
rect 31305 36924 31424 36958
rect 31458 36924 31489 36958
rect 31239 36868 31489 36924
rect 31239 36834 31271 36868
rect 31305 36834 31424 36868
rect 31458 36834 31489 36868
rect 31239 36778 31489 36834
rect 31239 36744 31271 36778
rect 31305 36744 31424 36778
rect 31458 36744 31489 36778
rect 31239 36688 31489 36744
rect 31239 36654 31271 36688
rect 31305 36654 31424 36688
rect 31458 36654 31489 36688
rect 31239 36598 31489 36654
rect 31239 36564 31271 36598
rect 31305 36564 31424 36598
rect 31458 36564 31489 36598
rect 31239 36508 31489 36564
rect 31239 36474 31271 36508
rect 31305 36474 31424 36508
rect 31458 36474 31489 36508
rect 31239 36418 31489 36474
rect 31239 36384 31271 36418
rect 31305 36384 31424 36418
rect 31458 36384 31489 36418
rect 31239 36328 31489 36384
rect 31239 36294 31271 36328
rect 31305 36294 31424 36328
rect 31458 36294 31489 36328
rect 28339 36222 28365 36227
rect 28328 36193 28365 36222
rect 28399 36193 28844 36222
rect 28328 36162 28844 36193
rect 30050 36204 30084 36238
rect 30118 36204 30149 36238
rect 30050 36187 30149 36204
rect 31239 36238 31489 36294
rect 31553 37196 32515 37213
rect 31553 37162 31574 37196
rect 31608 37162 31664 37196
rect 31698 37194 31754 37196
rect 31788 37194 31844 37196
rect 31878 37194 31934 37196
rect 31968 37194 32024 37196
rect 32058 37194 32114 37196
rect 32148 37194 32204 37196
rect 32238 37194 32294 37196
rect 32328 37194 32384 37196
rect 32418 37194 32474 37196
rect 31718 37162 31754 37194
rect 31808 37162 31844 37194
rect 31898 37162 31934 37194
rect 31988 37162 32024 37194
rect 32078 37162 32114 37194
rect 32168 37162 32204 37194
rect 32258 37162 32294 37194
rect 32348 37162 32384 37194
rect 32438 37162 32474 37194
rect 32508 37162 32515 37196
rect 31553 37160 31684 37162
rect 31718 37160 31774 37162
rect 31808 37160 31864 37162
rect 31898 37160 31954 37162
rect 31988 37160 32044 37162
rect 32078 37160 32134 37162
rect 32168 37160 32224 37162
rect 32258 37160 32314 37162
rect 32348 37160 32404 37162
rect 32438 37160 32515 37162
rect 31553 37141 32515 37160
rect 31553 37137 31625 37141
rect 31553 37103 31572 37137
rect 31606 37103 31625 37137
rect 31553 37047 31625 37103
rect 32443 37118 32515 37141
rect 32443 37084 32462 37118
rect 32496 37084 32515 37118
rect 31553 37013 31572 37047
rect 31606 37013 31625 37047
rect 31553 36957 31625 37013
rect 31553 36923 31572 36957
rect 31606 36923 31625 36957
rect 31553 36867 31625 36923
rect 31553 36833 31572 36867
rect 31606 36833 31625 36867
rect 31553 36777 31625 36833
rect 31553 36743 31572 36777
rect 31606 36743 31625 36777
rect 31553 36687 31625 36743
rect 31553 36653 31572 36687
rect 31606 36653 31625 36687
rect 31553 36597 31625 36653
rect 31553 36563 31572 36597
rect 31606 36563 31625 36597
rect 31553 36507 31625 36563
rect 31553 36473 31572 36507
rect 31606 36473 31625 36507
rect 31553 36417 31625 36473
rect 31553 36383 31572 36417
rect 31606 36383 31625 36417
rect 31687 37020 32381 37079
rect 31687 36986 31748 37020
rect 31782 36992 31838 37020
rect 31872 36992 31928 37020
rect 31962 36992 32018 37020
rect 31794 36986 31838 36992
rect 31894 36986 31928 36992
rect 31994 36986 32018 36992
rect 32052 36992 32108 37020
rect 32052 36986 32060 36992
rect 31687 36958 31760 36986
rect 31794 36958 31860 36986
rect 31894 36958 31960 36986
rect 31994 36958 32060 36986
rect 32094 36986 32108 36992
rect 32142 36992 32198 37020
rect 32142 36986 32160 36992
rect 32094 36958 32160 36986
rect 32194 36986 32198 36992
rect 32232 36992 32288 37020
rect 32232 36986 32260 36992
rect 32322 36986 32381 37020
rect 32194 36958 32260 36986
rect 32294 36958 32381 36986
rect 31687 36930 32381 36958
rect 31687 36896 31748 36930
rect 31782 36896 31838 36930
rect 31872 36896 31928 36930
rect 31962 36896 32018 36930
rect 32052 36896 32108 36930
rect 32142 36896 32198 36930
rect 32232 36896 32288 36930
rect 32322 36896 32381 36930
rect 31687 36892 32381 36896
rect 31687 36858 31760 36892
rect 31794 36858 31860 36892
rect 31894 36858 31960 36892
rect 31994 36858 32060 36892
rect 32094 36858 32160 36892
rect 32194 36858 32260 36892
rect 32294 36858 32381 36892
rect 31687 36840 32381 36858
rect 31687 36806 31748 36840
rect 31782 36806 31838 36840
rect 31872 36806 31928 36840
rect 31962 36806 32018 36840
rect 32052 36806 32108 36840
rect 32142 36806 32198 36840
rect 32232 36806 32288 36840
rect 32322 36806 32381 36840
rect 31687 36792 32381 36806
rect 31687 36758 31760 36792
rect 31794 36758 31860 36792
rect 31894 36758 31960 36792
rect 31994 36758 32060 36792
rect 32094 36758 32160 36792
rect 32194 36758 32260 36792
rect 32294 36758 32381 36792
rect 31687 36750 32381 36758
rect 31687 36716 31748 36750
rect 31782 36716 31838 36750
rect 31872 36716 31928 36750
rect 31962 36716 32018 36750
rect 32052 36716 32108 36750
rect 32142 36716 32198 36750
rect 32232 36716 32288 36750
rect 32322 36716 32381 36750
rect 31687 36692 32381 36716
rect 31687 36660 31760 36692
rect 31794 36660 31860 36692
rect 31894 36660 31960 36692
rect 31994 36660 32060 36692
rect 31687 36626 31748 36660
rect 31794 36658 31838 36660
rect 31894 36658 31928 36660
rect 31994 36658 32018 36660
rect 31782 36626 31838 36658
rect 31872 36626 31928 36658
rect 31962 36626 32018 36658
rect 32052 36658 32060 36660
rect 32094 36660 32160 36692
rect 32094 36658 32108 36660
rect 32052 36626 32108 36658
rect 32142 36658 32160 36660
rect 32194 36660 32260 36692
rect 32294 36660 32381 36692
rect 32194 36658 32198 36660
rect 32142 36626 32198 36658
rect 32232 36658 32260 36660
rect 32232 36626 32288 36658
rect 32322 36626 32381 36660
rect 31687 36592 32381 36626
rect 31687 36570 31760 36592
rect 31794 36570 31860 36592
rect 31894 36570 31960 36592
rect 31994 36570 32060 36592
rect 31687 36536 31748 36570
rect 31794 36558 31838 36570
rect 31894 36558 31928 36570
rect 31994 36558 32018 36570
rect 31782 36536 31838 36558
rect 31872 36536 31928 36558
rect 31962 36536 32018 36558
rect 32052 36558 32060 36570
rect 32094 36570 32160 36592
rect 32094 36558 32108 36570
rect 32052 36536 32108 36558
rect 32142 36558 32160 36570
rect 32194 36570 32260 36592
rect 32294 36570 32381 36592
rect 32194 36558 32198 36570
rect 32142 36536 32198 36558
rect 32232 36558 32260 36570
rect 32232 36536 32288 36558
rect 32322 36536 32381 36570
rect 31687 36492 32381 36536
rect 31687 36480 31760 36492
rect 31794 36480 31860 36492
rect 31894 36480 31960 36492
rect 31994 36480 32060 36492
rect 31687 36446 31748 36480
rect 31794 36458 31838 36480
rect 31894 36458 31928 36480
rect 31994 36458 32018 36480
rect 31782 36446 31838 36458
rect 31872 36446 31928 36458
rect 31962 36446 32018 36458
rect 32052 36458 32060 36480
rect 32094 36480 32160 36492
rect 32094 36458 32108 36480
rect 32052 36446 32108 36458
rect 32142 36458 32160 36480
rect 32194 36480 32260 36492
rect 32294 36480 32381 36492
rect 32194 36458 32198 36480
rect 32142 36446 32198 36458
rect 32232 36458 32260 36480
rect 32232 36446 32288 36458
rect 32322 36446 32381 36480
rect 31687 36385 32381 36446
rect 32443 37028 32515 37084
rect 32443 36994 32462 37028
rect 32496 36994 32515 37028
rect 32443 36938 32515 36994
rect 32443 36904 32462 36938
rect 32496 36904 32515 36938
rect 32443 36848 32515 36904
rect 32443 36814 32462 36848
rect 32496 36814 32515 36848
rect 32443 36758 32515 36814
rect 32443 36724 32462 36758
rect 32496 36724 32515 36758
rect 32443 36668 32515 36724
rect 32443 36634 32462 36668
rect 32496 36634 32515 36668
rect 32443 36578 32515 36634
rect 32443 36544 32462 36578
rect 32496 36544 32515 36578
rect 32443 36488 32515 36544
rect 32443 36454 32462 36488
rect 32496 36454 32515 36488
rect 32443 36398 32515 36454
rect 31553 36323 31625 36383
rect 32443 36364 32462 36398
rect 32496 36364 32515 36398
rect 32443 36323 32515 36364
rect 31553 36304 32515 36323
rect 31553 36270 31650 36304
rect 31684 36270 31740 36304
rect 31774 36270 31830 36304
rect 31864 36270 31920 36304
rect 31954 36270 32010 36304
rect 32044 36270 32100 36304
rect 32134 36270 32190 36304
rect 32224 36270 32280 36304
rect 32314 36270 32370 36304
rect 32404 36270 32515 36304
rect 31553 36251 32515 36270
rect 32579 37194 32611 37228
rect 32645 37194 32764 37228
rect 32798 37194 32829 37228
rect 33919 37228 34169 37277
rect 32579 37138 32829 37194
rect 32579 37104 32611 37138
rect 32645 37104 32764 37138
rect 32798 37104 32829 37138
rect 32579 37048 32829 37104
rect 32579 37014 32611 37048
rect 32645 37014 32764 37048
rect 32798 37014 32829 37048
rect 32579 36958 32829 37014
rect 32579 36924 32611 36958
rect 32645 36924 32764 36958
rect 32798 36924 32829 36958
rect 32579 36868 32829 36924
rect 32579 36834 32611 36868
rect 32645 36834 32764 36868
rect 32798 36834 32829 36868
rect 32579 36778 32829 36834
rect 32579 36744 32611 36778
rect 32645 36744 32764 36778
rect 32798 36744 32829 36778
rect 32579 36688 32829 36744
rect 32579 36654 32611 36688
rect 32645 36654 32764 36688
rect 32798 36654 32829 36688
rect 32579 36598 32829 36654
rect 32579 36564 32611 36598
rect 32645 36564 32764 36598
rect 32798 36564 32829 36598
rect 32579 36508 32829 36564
rect 32579 36474 32611 36508
rect 32645 36474 32764 36508
rect 32798 36474 32829 36508
rect 32579 36418 32829 36474
rect 32579 36384 32611 36418
rect 32645 36384 32764 36418
rect 32798 36384 32829 36418
rect 32579 36328 32829 36384
rect 32579 36294 32611 36328
rect 32645 36294 32764 36328
rect 32798 36294 32829 36328
rect 31239 36204 31271 36238
rect 31305 36204 31424 36238
rect 31458 36204 31489 36238
rect 31239 36187 31489 36204
rect 32579 36238 32829 36294
rect 32893 37196 33855 37213
rect 32893 37162 32914 37196
rect 32948 37162 33004 37196
rect 33038 37194 33094 37196
rect 33128 37194 33184 37196
rect 33218 37194 33274 37196
rect 33308 37194 33364 37196
rect 33398 37194 33454 37196
rect 33488 37194 33544 37196
rect 33578 37194 33634 37196
rect 33668 37194 33724 37196
rect 33758 37194 33814 37196
rect 33058 37162 33094 37194
rect 33148 37162 33184 37194
rect 33238 37162 33274 37194
rect 33328 37162 33364 37194
rect 33418 37162 33454 37194
rect 33508 37162 33544 37194
rect 33598 37162 33634 37194
rect 33688 37162 33724 37194
rect 33778 37162 33814 37194
rect 33848 37162 33855 37196
rect 32893 37160 33024 37162
rect 33058 37160 33114 37162
rect 33148 37160 33204 37162
rect 33238 37160 33294 37162
rect 33328 37160 33384 37162
rect 33418 37160 33474 37162
rect 33508 37160 33564 37162
rect 33598 37160 33654 37162
rect 33688 37160 33744 37162
rect 33778 37160 33855 37162
rect 32893 37141 33855 37160
rect 32893 37137 32965 37141
rect 32893 37103 32912 37137
rect 32946 37103 32965 37137
rect 32893 37047 32965 37103
rect 33783 37118 33855 37141
rect 33783 37084 33802 37118
rect 33836 37084 33855 37118
rect 32893 37013 32912 37047
rect 32946 37013 32965 37047
rect 32893 36957 32965 37013
rect 32893 36923 32912 36957
rect 32946 36923 32965 36957
rect 32893 36867 32965 36923
rect 32893 36833 32912 36867
rect 32946 36833 32965 36867
rect 32893 36777 32965 36833
rect 32893 36743 32912 36777
rect 32946 36743 32965 36777
rect 32893 36687 32965 36743
rect 32893 36653 32912 36687
rect 32946 36653 32965 36687
rect 32893 36597 32965 36653
rect 32893 36563 32912 36597
rect 32946 36563 32965 36597
rect 32893 36507 32965 36563
rect 32893 36473 32912 36507
rect 32946 36473 32965 36507
rect 32893 36417 32965 36473
rect 32893 36383 32912 36417
rect 32946 36383 32965 36417
rect 33027 37020 33721 37079
rect 33027 36986 33088 37020
rect 33122 36992 33178 37020
rect 33212 36992 33268 37020
rect 33302 36992 33358 37020
rect 33134 36986 33178 36992
rect 33234 36986 33268 36992
rect 33334 36986 33358 36992
rect 33392 36992 33448 37020
rect 33392 36986 33400 36992
rect 33027 36958 33100 36986
rect 33134 36958 33200 36986
rect 33234 36958 33300 36986
rect 33334 36958 33400 36986
rect 33434 36986 33448 36992
rect 33482 36992 33538 37020
rect 33482 36986 33500 36992
rect 33434 36958 33500 36986
rect 33534 36986 33538 36992
rect 33572 36992 33628 37020
rect 33572 36986 33600 36992
rect 33662 36986 33721 37020
rect 33534 36958 33600 36986
rect 33634 36958 33721 36986
rect 33027 36930 33721 36958
rect 33027 36896 33088 36930
rect 33122 36896 33178 36930
rect 33212 36896 33268 36930
rect 33302 36896 33358 36930
rect 33392 36896 33448 36930
rect 33482 36896 33538 36930
rect 33572 36896 33628 36930
rect 33662 36896 33721 36930
rect 33027 36892 33721 36896
rect 33027 36858 33100 36892
rect 33134 36858 33200 36892
rect 33234 36858 33300 36892
rect 33334 36858 33400 36892
rect 33434 36858 33500 36892
rect 33534 36858 33600 36892
rect 33634 36858 33721 36892
rect 33027 36840 33721 36858
rect 33027 36806 33088 36840
rect 33122 36806 33178 36840
rect 33212 36806 33268 36840
rect 33302 36806 33358 36840
rect 33392 36806 33448 36840
rect 33482 36806 33538 36840
rect 33572 36806 33628 36840
rect 33662 36806 33721 36840
rect 33027 36792 33721 36806
rect 33027 36758 33100 36792
rect 33134 36758 33200 36792
rect 33234 36758 33300 36792
rect 33334 36758 33400 36792
rect 33434 36758 33500 36792
rect 33534 36758 33600 36792
rect 33634 36758 33721 36792
rect 33027 36750 33721 36758
rect 33027 36716 33088 36750
rect 33122 36716 33178 36750
rect 33212 36716 33268 36750
rect 33302 36716 33358 36750
rect 33392 36716 33448 36750
rect 33482 36716 33538 36750
rect 33572 36716 33628 36750
rect 33662 36716 33721 36750
rect 33027 36692 33721 36716
rect 33027 36660 33100 36692
rect 33134 36660 33200 36692
rect 33234 36660 33300 36692
rect 33334 36660 33400 36692
rect 33027 36626 33088 36660
rect 33134 36658 33178 36660
rect 33234 36658 33268 36660
rect 33334 36658 33358 36660
rect 33122 36626 33178 36658
rect 33212 36626 33268 36658
rect 33302 36626 33358 36658
rect 33392 36658 33400 36660
rect 33434 36660 33500 36692
rect 33434 36658 33448 36660
rect 33392 36626 33448 36658
rect 33482 36658 33500 36660
rect 33534 36660 33600 36692
rect 33634 36660 33721 36692
rect 33534 36658 33538 36660
rect 33482 36626 33538 36658
rect 33572 36658 33600 36660
rect 33572 36626 33628 36658
rect 33662 36626 33721 36660
rect 33027 36592 33721 36626
rect 33027 36570 33100 36592
rect 33134 36570 33200 36592
rect 33234 36570 33300 36592
rect 33334 36570 33400 36592
rect 33027 36536 33088 36570
rect 33134 36558 33178 36570
rect 33234 36558 33268 36570
rect 33334 36558 33358 36570
rect 33122 36536 33178 36558
rect 33212 36536 33268 36558
rect 33302 36536 33358 36558
rect 33392 36558 33400 36570
rect 33434 36570 33500 36592
rect 33434 36558 33448 36570
rect 33392 36536 33448 36558
rect 33482 36558 33500 36570
rect 33534 36570 33600 36592
rect 33634 36570 33721 36592
rect 33534 36558 33538 36570
rect 33482 36536 33538 36558
rect 33572 36558 33600 36570
rect 33572 36536 33628 36558
rect 33662 36536 33721 36570
rect 33027 36492 33721 36536
rect 33027 36480 33100 36492
rect 33134 36480 33200 36492
rect 33234 36480 33300 36492
rect 33334 36480 33400 36492
rect 33027 36446 33088 36480
rect 33134 36458 33178 36480
rect 33234 36458 33268 36480
rect 33334 36458 33358 36480
rect 33122 36446 33178 36458
rect 33212 36446 33268 36458
rect 33302 36446 33358 36458
rect 33392 36458 33400 36480
rect 33434 36480 33500 36492
rect 33434 36458 33448 36480
rect 33392 36446 33448 36458
rect 33482 36458 33500 36480
rect 33534 36480 33600 36492
rect 33634 36480 33721 36492
rect 33534 36458 33538 36480
rect 33482 36446 33538 36458
rect 33572 36458 33600 36480
rect 33572 36446 33628 36458
rect 33662 36446 33721 36480
rect 33027 36385 33721 36446
rect 33783 37028 33855 37084
rect 33783 36994 33802 37028
rect 33836 36994 33855 37028
rect 33783 36938 33855 36994
rect 33783 36904 33802 36938
rect 33836 36904 33855 36938
rect 33783 36848 33855 36904
rect 33783 36814 33802 36848
rect 33836 36814 33855 36848
rect 33783 36758 33855 36814
rect 33783 36724 33802 36758
rect 33836 36724 33855 36758
rect 33783 36668 33855 36724
rect 33783 36634 33802 36668
rect 33836 36634 33855 36668
rect 33783 36578 33855 36634
rect 33783 36544 33802 36578
rect 33836 36544 33855 36578
rect 33783 36488 33855 36544
rect 33783 36454 33802 36488
rect 33836 36454 33855 36488
rect 33783 36398 33855 36454
rect 32893 36323 32965 36383
rect 33783 36364 33802 36398
rect 33836 36364 33855 36398
rect 33783 36323 33855 36364
rect 32893 36304 33855 36323
rect 32893 36270 32990 36304
rect 33024 36270 33080 36304
rect 33114 36270 33170 36304
rect 33204 36270 33260 36304
rect 33294 36270 33350 36304
rect 33384 36270 33440 36304
rect 33474 36270 33530 36304
rect 33564 36270 33620 36304
rect 33654 36270 33710 36304
rect 33744 36270 33855 36304
rect 32893 36251 33855 36270
rect 33919 37194 33951 37228
rect 33985 37194 34104 37228
rect 34138 37194 34169 37228
rect 35259 37228 35509 37277
rect 33919 37138 34169 37194
rect 33919 37104 33951 37138
rect 33985 37104 34104 37138
rect 34138 37104 34169 37138
rect 33919 37048 34169 37104
rect 33919 37014 33951 37048
rect 33985 37014 34104 37048
rect 34138 37014 34169 37048
rect 33919 36958 34169 37014
rect 33919 36924 33951 36958
rect 33985 36924 34104 36958
rect 34138 36924 34169 36958
rect 33919 36868 34169 36924
rect 33919 36834 33951 36868
rect 33985 36834 34104 36868
rect 34138 36834 34169 36868
rect 33919 36778 34169 36834
rect 33919 36744 33951 36778
rect 33985 36744 34104 36778
rect 34138 36744 34169 36778
rect 33919 36688 34169 36744
rect 33919 36654 33951 36688
rect 33985 36654 34104 36688
rect 34138 36654 34169 36688
rect 33919 36598 34169 36654
rect 33919 36564 33951 36598
rect 33985 36564 34104 36598
rect 34138 36564 34169 36598
rect 33919 36508 34169 36564
rect 33919 36474 33951 36508
rect 33985 36474 34104 36508
rect 34138 36474 34169 36508
rect 33919 36418 34169 36474
rect 33919 36384 33951 36418
rect 33985 36384 34104 36418
rect 34138 36384 34169 36418
rect 33919 36328 34169 36384
rect 33919 36294 33951 36328
rect 33985 36294 34104 36328
rect 34138 36294 34169 36328
rect 32579 36204 32611 36238
rect 32645 36204 32764 36238
rect 32798 36204 32829 36238
rect 32579 36187 32829 36204
rect 33919 36238 34169 36294
rect 34233 37196 35195 37213
rect 34233 37162 34254 37196
rect 34288 37162 34344 37196
rect 34378 37194 34434 37196
rect 34468 37194 34524 37196
rect 34558 37194 34614 37196
rect 34648 37194 34704 37196
rect 34738 37194 34794 37196
rect 34828 37194 34884 37196
rect 34918 37194 34974 37196
rect 35008 37194 35064 37196
rect 35098 37194 35154 37196
rect 34398 37162 34434 37194
rect 34488 37162 34524 37194
rect 34578 37162 34614 37194
rect 34668 37162 34704 37194
rect 34758 37162 34794 37194
rect 34848 37162 34884 37194
rect 34938 37162 34974 37194
rect 35028 37162 35064 37194
rect 35118 37162 35154 37194
rect 35188 37162 35195 37196
rect 34233 37160 34364 37162
rect 34398 37160 34454 37162
rect 34488 37160 34544 37162
rect 34578 37160 34634 37162
rect 34668 37160 34724 37162
rect 34758 37160 34814 37162
rect 34848 37160 34904 37162
rect 34938 37160 34994 37162
rect 35028 37160 35084 37162
rect 35118 37160 35195 37162
rect 34233 37141 35195 37160
rect 34233 37137 34305 37141
rect 34233 37103 34252 37137
rect 34286 37103 34305 37137
rect 34233 37047 34305 37103
rect 35123 37118 35195 37141
rect 35123 37084 35142 37118
rect 35176 37084 35195 37118
rect 34233 37013 34252 37047
rect 34286 37013 34305 37047
rect 34233 36957 34305 37013
rect 34233 36923 34252 36957
rect 34286 36923 34305 36957
rect 34233 36867 34305 36923
rect 34233 36833 34252 36867
rect 34286 36833 34305 36867
rect 34233 36777 34305 36833
rect 34233 36743 34252 36777
rect 34286 36743 34305 36777
rect 34233 36687 34305 36743
rect 34233 36653 34252 36687
rect 34286 36653 34305 36687
rect 34233 36597 34305 36653
rect 34233 36563 34252 36597
rect 34286 36563 34305 36597
rect 34233 36507 34305 36563
rect 34233 36473 34252 36507
rect 34286 36473 34305 36507
rect 34233 36417 34305 36473
rect 34233 36383 34252 36417
rect 34286 36383 34305 36417
rect 34367 37020 35061 37079
rect 34367 36986 34428 37020
rect 34462 36992 34518 37020
rect 34552 36992 34608 37020
rect 34642 36992 34698 37020
rect 34474 36986 34518 36992
rect 34574 36986 34608 36992
rect 34674 36986 34698 36992
rect 34732 36992 34788 37020
rect 34732 36986 34740 36992
rect 34367 36958 34440 36986
rect 34474 36958 34540 36986
rect 34574 36958 34640 36986
rect 34674 36958 34740 36986
rect 34774 36986 34788 36992
rect 34822 36992 34878 37020
rect 34822 36986 34840 36992
rect 34774 36958 34840 36986
rect 34874 36986 34878 36992
rect 34912 36992 34968 37020
rect 34912 36986 34940 36992
rect 35002 36986 35061 37020
rect 34874 36958 34940 36986
rect 34974 36958 35061 36986
rect 34367 36930 35061 36958
rect 34367 36896 34428 36930
rect 34462 36896 34518 36930
rect 34552 36896 34608 36930
rect 34642 36896 34698 36930
rect 34732 36896 34788 36930
rect 34822 36896 34878 36930
rect 34912 36896 34968 36930
rect 35002 36896 35061 36930
rect 34367 36892 35061 36896
rect 34367 36858 34440 36892
rect 34474 36858 34540 36892
rect 34574 36858 34640 36892
rect 34674 36858 34740 36892
rect 34774 36858 34840 36892
rect 34874 36858 34940 36892
rect 34974 36858 35061 36892
rect 34367 36840 35061 36858
rect 34367 36806 34428 36840
rect 34462 36806 34518 36840
rect 34552 36806 34608 36840
rect 34642 36806 34698 36840
rect 34732 36806 34788 36840
rect 34822 36806 34878 36840
rect 34912 36806 34968 36840
rect 35002 36806 35061 36840
rect 34367 36792 35061 36806
rect 34367 36758 34440 36792
rect 34474 36758 34540 36792
rect 34574 36758 34640 36792
rect 34674 36758 34740 36792
rect 34774 36758 34840 36792
rect 34874 36758 34940 36792
rect 34974 36758 35061 36792
rect 34367 36750 35061 36758
rect 34367 36716 34428 36750
rect 34462 36716 34518 36750
rect 34552 36716 34608 36750
rect 34642 36716 34698 36750
rect 34732 36716 34788 36750
rect 34822 36716 34878 36750
rect 34912 36716 34968 36750
rect 35002 36716 35061 36750
rect 34367 36692 35061 36716
rect 34367 36660 34440 36692
rect 34474 36660 34540 36692
rect 34574 36660 34640 36692
rect 34674 36660 34740 36692
rect 34367 36626 34428 36660
rect 34474 36658 34518 36660
rect 34574 36658 34608 36660
rect 34674 36658 34698 36660
rect 34462 36626 34518 36658
rect 34552 36626 34608 36658
rect 34642 36626 34698 36658
rect 34732 36658 34740 36660
rect 34774 36660 34840 36692
rect 34774 36658 34788 36660
rect 34732 36626 34788 36658
rect 34822 36658 34840 36660
rect 34874 36660 34940 36692
rect 34974 36660 35061 36692
rect 34874 36658 34878 36660
rect 34822 36626 34878 36658
rect 34912 36658 34940 36660
rect 34912 36626 34968 36658
rect 35002 36626 35061 36660
rect 34367 36592 35061 36626
rect 34367 36570 34440 36592
rect 34474 36570 34540 36592
rect 34574 36570 34640 36592
rect 34674 36570 34740 36592
rect 34367 36536 34428 36570
rect 34474 36558 34518 36570
rect 34574 36558 34608 36570
rect 34674 36558 34698 36570
rect 34462 36536 34518 36558
rect 34552 36536 34608 36558
rect 34642 36536 34698 36558
rect 34732 36558 34740 36570
rect 34774 36570 34840 36592
rect 34774 36558 34788 36570
rect 34732 36536 34788 36558
rect 34822 36558 34840 36570
rect 34874 36570 34940 36592
rect 34974 36570 35061 36592
rect 34874 36558 34878 36570
rect 34822 36536 34878 36558
rect 34912 36558 34940 36570
rect 34912 36536 34968 36558
rect 35002 36536 35061 36570
rect 34367 36492 35061 36536
rect 34367 36480 34440 36492
rect 34474 36480 34540 36492
rect 34574 36480 34640 36492
rect 34674 36480 34740 36492
rect 34367 36446 34428 36480
rect 34474 36458 34518 36480
rect 34574 36458 34608 36480
rect 34674 36458 34698 36480
rect 34462 36446 34518 36458
rect 34552 36446 34608 36458
rect 34642 36446 34698 36458
rect 34732 36458 34740 36480
rect 34774 36480 34840 36492
rect 34774 36458 34788 36480
rect 34732 36446 34788 36458
rect 34822 36458 34840 36480
rect 34874 36480 34940 36492
rect 34974 36480 35061 36492
rect 34874 36458 34878 36480
rect 34822 36446 34878 36458
rect 34912 36458 34940 36480
rect 34912 36446 34968 36458
rect 35002 36446 35061 36480
rect 34367 36385 35061 36446
rect 35123 37028 35195 37084
rect 35123 36994 35142 37028
rect 35176 36994 35195 37028
rect 35123 36938 35195 36994
rect 35123 36904 35142 36938
rect 35176 36904 35195 36938
rect 35123 36848 35195 36904
rect 35123 36814 35142 36848
rect 35176 36814 35195 36848
rect 35123 36758 35195 36814
rect 35123 36724 35142 36758
rect 35176 36724 35195 36758
rect 35123 36668 35195 36724
rect 35123 36634 35142 36668
rect 35176 36634 35195 36668
rect 35123 36578 35195 36634
rect 35123 36544 35142 36578
rect 35176 36544 35195 36578
rect 35123 36488 35195 36544
rect 35123 36454 35142 36488
rect 35176 36454 35195 36488
rect 35123 36398 35195 36454
rect 34233 36323 34305 36383
rect 35123 36364 35142 36398
rect 35176 36364 35195 36398
rect 35123 36323 35195 36364
rect 34233 36304 35195 36323
rect 34233 36270 34330 36304
rect 34364 36270 34420 36304
rect 34454 36270 34510 36304
rect 34544 36270 34600 36304
rect 34634 36270 34690 36304
rect 34724 36270 34780 36304
rect 34814 36270 34870 36304
rect 34904 36270 34960 36304
rect 34994 36270 35050 36304
rect 35084 36270 35195 36304
rect 34233 36251 35195 36270
rect 35259 37194 35291 37228
rect 35325 37194 35444 37228
rect 35478 37194 35509 37228
rect 36599 37228 36849 37277
rect 35259 37138 35509 37194
rect 35259 37104 35291 37138
rect 35325 37104 35444 37138
rect 35478 37104 35509 37138
rect 35259 37048 35509 37104
rect 35259 37014 35291 37048
rect 35325 37014 35444 37048
rect 35478 37014 35509 37048
rect 35259 36958 35509 37014
rect 35259 36924 35291 36958
rect 35325 36924 35444 36958
rect 35478 36924 35509 36958
rect 35259 36868 35509 36924
rect 35259 36834 35291 36868
rect 35325 36834 35444 36868
rect 35478 36834 35509 36868
rect 35259 36778 35509 36834
rect 35259 36744 35291 36778
rect 35325 36744 35444 36778
rect 35478 36744 35509 36778
rect 35259 36688 35509 36744
rect 35259 36654 35291 36688
rect 35325 36654 35444 36688
rect 35478 36654 35509 36688
rect 35259 36598 35509 36654
rect 35259 36564 35291 36598
rect 35325 36564 35444 36598
rect 35478 36564 35509 36598
rect 35259 36508 35509 36564
rect 35259 36474 35291 36508
rect 35325 36474 35444 36508
rect 35478 36474 35509 36508
rect 35259 36418 35509 36474
rect 35259 36384 35291 36418
rect 35325 36384 35444 36418
rect 35478 36384 35509 36418
rect 35259 36328 35509 36384
rect 35259 36294 35291 36328
rect 35325 36294 35444 36328
rect 35478 36294 35509 36328
rect 33919 36204 33951 36238
rect 33985 36204 34104 36238
rect 34138 36204 34169 36238
rect 33919 36187 34169 36204
rect 35259 36238 35509 36294
rect 35573 37196 36535 37213
rect 35573 37162 35594 37196
rect 35628 37162 35684 37196
rect 35718 37194 35774 37196
rect 35808 37194 35864 37196
rect 35898 37194 35954 37196
rect 35988 37194 36044 37196
rect 36078 37194 36134 37196
rect 36168 37194 36224 37196
rect 36258 37194 36314 37196
rect 36348 37194 36404 37196
rect 36438 37194 36494 37196
rect 35738 37162 35774 37194
rect 35828 37162 35864 37194
rect 35918 37162 35954 37194
rect 36008 37162 36044 37194
rect 36098 37162 36134 37194
rect 36188 37162 36224 37194
rect 36278 37162 36314 37194
rect 36368 37162 36404 37194
rect 36458 37162 36494 37194
rect 36528 37162 36535 37196
rect 35573 37160 35704 37162
rect 35738 37160 35794 37162
rect 35828 37160 35884 37162
rect 35918 37160 35974 37162
rect 36008 37160 36064 37162
rect 36098 37160 36154 37162
rect 36188 37160 36244 37162
rect 36278 37160 36334 37162
rect 36368 37160 36424 37162
rect 36458 37160 36535 37162
rect 35573 37141 36535 37160
rect 35573 37137 35645 37141
rect 35573 37103 35592 37137
rect 35626 37103 35645 37137
rect 35573 37047 35645 37103
rect 36463 37118 36535 37141
rect 36463 37084 36482 37118
rect 36516 37084 36535 37118
rect 35573 37013 35592 37047
rect 35626 37013 35645 37047
rect 35573 36957 35645 37013
rect 35573 36923 35592 36957
rect 35626 36923 35645 36957
rect 35573 36867 35645 36923
rect 35573 36833 35592 36867
rect 35626 36833 35645 36867
rect 35573 36777 35645 36833
rect 35573 36743 35592 36777
rect 35626 36743 35645 36777
rect 35573 36687 35645 36743
rect 35573 36653 35592 36687
rect 35626 36653 35645 36687
rect 35573 36597 35645 36653
rect 35573 36563 35592 36597
rect 35626 36563 35645 36597
rect 35573 36507 35645 36563
rect 35573 36473 35592 36507
rect 35626 36473 35645 36507
rect 35573 36417 35645 36473
rect 35573 36383 35592 36417
rect 35626 36383 35645 36417
rect 35707 37020 36401 37079
rect 35707 36986 35768 37020
rect 35802 36992 35858 37020
rect 35892 36992 35948 37020
rect 35982 36992 36038 37020
rect 35814 36986 35858 36992
rect 35914 36986 35948 36992
rect 36014 36986 36038 36992
rect 36072 36992 36128 37020
rect 36072 36986 36080 36992
rect 35707 36958 35780 36986
rect 35814 36958 35880 36986
rect 35914 36958 35980 36986
rect 36014 36958 36080 36986
rect 36114 36986 36128 36992
rect 36162 36992 36218 37020
rect 36162 36986 36180 36992
rect 36114 36958 36180 36986
rect 36214 36986 36218 36992
rect 36252 36992 36308 37020
rect 36252 36986 36280 36992
rect 36342 36986 36401 37020
rect 36214 36958 36280 36986
rect 36314 36958 36401 36986
rect 35707 36930 36401 36958
rect 35707 36896 35768 36930
rect 35802 36896 35858 36930
rect 35892 36896 35948 36930
rect 35982 36896 36038 36930
rect 36072 36896 36128 36930
rect 36162 36896 36218 36930
rect 36252 36896 36308 36930
rect 36342 36896 36401 36930
rect 35707 36892 36401 36896
rect 35707 36858 35780 36892
rect 35814 36858 35880 36892
rect 35914 36858 35980 36892
rect 36014 36858 36080 36892
rect 36114 36858 36180 36892
rect 36214 36858 36280 36892
rect 36314 36858 36401 36892
rect 35707 36840 36401 36858
rect 35707 36806 35768 36840
rect 35802 36806 35858 36840
rect 35892 36806 35948 36840
rect 35982 36806 36038 36840
rect 36072 36806 36128 36840
rect 36162 36806 36218 36840
rect 36252 36806 36308 36840
rect 36342 36806 36401 36840
rect 35707 36792 36401 36806
rect 35707 36758 35780 36792
rect 35814 36758 35880 36792
rect 35914 36758 35980 36792
rect 36014 36758 36080 36792
rect 36114 36758 36180 36792
rect 36214 36758 36280 36792
rect 36314 36758 36401 36792
rect 35707 36750 36401 36758
rect 35707 36716 35768 36750
rect 35802 36716 35858 36750
rect 35892 36716 35948 36750
rect 35982 36716 36038 36750
rect 36072 36716 36128 36750
rect 36162 36716 36218 36750
rect 36252 36716 36308 36750
rect 36342 36716 36401 36750
rect 35707 36692 36401 36716
rect 35707 36660 35780 36692
rect 35814 36660 35880 36692
rect 35914 36660 35980 36692
rect 36014 36660 36080 36692
rect 35707 36626 35768 36660
rect 35814 36658 35858 36660
rect 35914 36658 35948 36660
rect 36014 36658 36038 36660
rect 35802 36626 35858 36658
rect 35892 36626 35948 36658
rect 35982 36626 36038 36658
rect 36072 36658 36080 36660
rect 36114 36660 36180 36692
rect 36114 36658 36128 36660
rect 36072 36626 36128 36658
rect 36162 36658 36180 36660
rect 36214 36660 36280 36692
rect 36314 36660 36401 36692
rect 36214 36658 36218 36660
rect 36162 36626 36218 36658
rect 36252 36658 36280 36660
rect 36252 36626 36308 36658
rect 36342 36626 36401 36660
rect 35707 36592 36401 36626
rect 35707 36570 35780 36592
rect 35814 36570 35880 36592
rect 35914 36570 35980 36592
rect 36014 36570 36080 36592
rect 35707 36536 35768 36570
rect 35814 36558 35858 36570
rect 35914 36558 35948 36570
rect 36014 36558 36038 36570
rect 35802 36536 35858 36558
rect 35892 36536 35948 36558
rect 35982 36536 36038 36558
rect 36072 36558 36080 36570
rect 36114 36570 36180 36592
rect 36114 36558 36128 36570
rect 36072 36536 36128 36558
rect 36162 36558 36180 36570
rect 36214 36570 36280 36592
rect 36314 36570 36401 36592
rect 36214 36558 36218 36570
rect 36162 36536 36218 36558
rect 36252 36558 36280 36570
rect 36252 36536 36308 36558
rect 36342 36536 36401 36570
rect 35707 36492 36401 36536
rect 35707 36480 35780 36492
rect 35814 36480 35880 36492
rect 35914 36480 35980 36492
rect 36014 36480 36080 36492
rect 35707 36446 35768 36480
rect 35814 36458 35858 36480
rect 35914 36458 35948 36480
rect 36014 36458 36038 36480
rect 35802 36446 35858 36458
rect 35892 36446 35948 36458
rect 35982 36446 36038 36458
rect 36072 36458 36080 36480
rect 36114 36480 36180 36492
rect 36114 36458 36128 36480
rect 36072 36446 36128 36458
rect 36162 36458 36180 36480
rect 36214 36480 36280 36492
rect 36314 36480 36401 36492
rect 36214 36458 36218 36480
rect 36162 36446 36218 36458
rect 36252 36458 36280 36480
rect 36252 36446 36308 36458
rect 36342 36446 36401 36480
rect 35707 36385 36401 36446
rect 36463 37028 36535 37084
rect 36463 36994 36482 37028
rect 36516 36994 36535 37028
rect 36463 36938 36535 36994
rect 36463 36904 36482 36938
rect 36516 36904 36535 36938
rect 36463 36848 36535 36904
rect 36463 36814 36482 36848
rect 36516 36814 36535 36848
rect 36463 36758 36535 36814
rect 36463 36724 36482 36758
rect 36516 36724 36535 36758
rect 36463 36668 36535 36724
rect 36463 36634 36482 36668
rect 36516 36634 36535 36668
rect 36463 36578 36535 36634
rect 36463 36544 36482 36578
rect 36516 36544 36535 36578
rect 36463 36488 36535 36544
rect 36463 36454 36482 36488
rect 36516 36454 36535 36488
rect 36463 36398 36535 36454
rect 35573 36323 35645 36383
rect 36463 36364 36482 36398
rect 36516 36364 36535 36398
rect 36463 36323 36535 36364
rect 35573 36304 36535 36323
rect 35573 36270 35670 36304
rect 35704 36270 35760 36304
rect 35794 36270 35850 36304
rect 35884 36270 35940 36304
rect 35974 36270 36030 36304
rect 36064 36270 36120 36304
rect 36154 36270 36210 36304
rect 36244 36270 36300 36304
rect 36334 36270 36390 36304
rect 36424 36270 36535 36304
rect 35573 36251 36535 36270
rect 36599 37194 36631 37228
rect 36665 37194 36784 37228
rect 36818 37194 36849 37228
rect 37939 37228 38189 37277
rect 36599 37138 36849 37194
rect 36599 37104 36631 37138
rect 36665 37104 36784 37138
rect 36818 37104 36849 37138
rect 36599 37048 36849 37104
rect 36599 37014 36631 37048
rect 36665 37014 36784 37048
rect 36818 37014 36849 37048
rect 36599 36958 36849 37014
rect 36599 36924 36631 36958
rect 36665 36924 36784 36958
rect 36818 36924 36849 36958
rect 36599 36868 36849 36924
rect 36599 36834 36631 36868
rect 36665 36834 36784 36868
rect 36818 36834 36849 36868
rect 36599 36778 36849 36834
rect 36599 36744 36631 36778
rect 36665 36744 36784 36778
rect 36818 36744 36849 36778
rect 36599 36688 36849 36744
rect 36599 36654 36631 36688
rect 36665 36654 36784 36688
rect 36818 36654 36849 36688
rect 36599 36598 36849 36654
rect 36599 36564 36631 36598
rect 36665 36564 36784 36598
rect 36818 36564 36849 36598
rect 36599 36508 36849 36564
rect 36599 36474 36631 36508
rect 36665 36474 36784 36508
rect 36818 36474 36849 36508
rect 36599 36418 36849 36474
rect 36599 36384 36631 36418
rect 36665 36384 36784 36418
rect 36818 36384 36849 36418
rect 36599 36328 36849 36384
rect 36599 36294 36631 36328
rect 36665 36294 36784 36328
rect 36818 36294 36849 36328
rect 35259 36204 35291 36238
rect 35325 36204 35444 36238
rect 35478 36204 35509 36238
rect 35259 36187 35509 36204
rect 36599 36238 36849 36294
rect 36913 37196 37875 37213
rect 36913 37162 36934 37196
rect 36968 37162 37024 37196
rect 37058 37194 37114 37196
rect 37148 37194 37204 37196
rect 37238 37194 37294 37196
rect 37328 37194 37384 37196
rect 37418 37194 37474 37196
rect 37508 37194 37564 37196
rect 37598 37194 37654 37196
rect 37688 37194 37744 37196
rect 37778 37194 37834 37196
rect 37078 37162 37114 37194
rect 37168 37162 37204 37194
rect 37258 37162 37294 37194
rect 37348 37162 37384 37194
rect 37438 37162 37474 37194
rect 37528 37162 37564 37194
rect 37618 37162 37654 37194
rect 37708 37162 37744 37194
rect 37798 37162 37834 37194
rect 37868 37162 37875 37196
rect 36913 37160 37044 37162
rect 37078 37160 37134 37162
rect 37168 37160 37224 37162
rect 37258 37160 37314 37162
rect 37348 37160 37404 37162
rect 37438 37160 37494 37162
rect 37528 37160 37584 37162
rect 37618 37160 37674 37162
rect 37708 37160 37764 37162
rect 37798 37160 37875 37162
rect 36913 37141 37875 37160
rect 36913 37137 36985 37141
rect 36913 37103 36932 37137
rect 36966 37103 36985 37137
rect 36913 37047 36985 37103
rect 37803 37118 37875 37141
rect 37803 37084 37822 37118
rect 37856 37084 37875 37118
rect 36913 37013 36932 37047
rect 36966 37013 36985 37047
rect 36913 36957 36985 37013
rect 36913 36923 36932 36957
rect 36966 36923 36985 36957
rect 36913 36867 36985 36923
rect 36913 36833 36932 36867
rect 36966 36833 36985 36867
rect 36913 36777 36985 36833
rect 36913 36743 36932 36777
rect 36966 36743 36985 36777
rect 36913 36687 36985 36743
rect 36913 36653 36932 36687
rect 36966 36653 36985 36687
rect 36913 36597 36985 36653
rect 36913 36563 36932 36597
rect 36966 36563 36985 36597
rect 36913 36507 36985 36563
rect 36913 36473 36932 36507
rect 36966 36473 36985 36507
rect 36913 36417 36985 36473
rect 36913 36383 36932 36417
rect 36966 36383 36985 36417
rect 37047 37020 37741 37079
rect 37047 36986 37108 37020
rect 37142 36992 37198 37020
rect 37232 36992 37288 37020
rect 37322 36992 37378 37020
rect 37154 36986 37198 36992
rect 37254 36986 37288 36992
rect 37354 36986 37378 36992
rect 37412 36992 37468 37020
rect 37412 36986 37420 36992
rect 37047 36958 37120 36986
rect 37154 36958 37220 36986
rect 37254 36958 37320 36986
rect 37354 36958 37420 36986
rect 37454 36986 37468 36992
rect 37502 36992 37558 37020
rect 37502 36986 37520 36992
rect 37454 36958 37520 36986
rect 37554 36986 37558 36992
rect 37592 36992 37648 37020
rect 37592 36986 37620 36992
rect 37682 36986 37741 37020
rect 37554 36958 37620 36986
rect 37654 36958 37741 36986
rect 37047 36930 37741 36958
rect 37047 36896 37108 36930
rect 37142 36896 37198 36930
rect 37232 36896 37288 36930
rect 37322 36896 37378 36930
rect 37412 36896 37468 36930
rect 37502 36896 37558 36930
rect 37592 36896 37648 36930
rect 37682 36896 37741 36930
rect 37047 36892 37741 36896
rect 37047 36858 37120 36892
rect 37154 36858 37220 36892
rect 37254 36858 37320 36892
rect 37354 36858 37420 36892
rect 37454 36858 37520 36892
rect 37554 36858 37620 36892
rect 37654 36858 37741 36892
rect 37047 36840 37741 36858
rect 37047 36806 37108 36840
rect 37142 36806 37198 36840
rect 37232 36806 37288 36840
rect 37322 36806 37378 36840
rect 37412 36806 37468 36840
rect 37502 36806 37558 36840
rect 37592 36806 37648 36840
rect 37682 36806 37741 36840
rect 37047 36792 37741 36806
rect 37047 36758 37120 36792
rect 37154 36758 37220 36792
rect 37254 36758 37320 36792
rect 37354 36758 37420 36792
rect 37454 36758 37520 36792
rect 37554 36758 37620 36792
rect 37654 36758 37741 36792
rect 37047 36750 37741 36758
rect 37047 36716 37108 36750
rect 37142 36716 37198 36750
rect 37232 36716 37288 36750
rect 37322 36716 37378 36750
rect 37412 36716 37468 36750
rect 37502 36716 37558 36750
rect 37592 36716 37648 36750
rect 37682 36716 37741 36750
rect 37047 36692 37741 36716
rect 37047 36660 37120 36692
rect 37154 36660 37220 36692
rect 37254 36660 37320 36692
rect 37354 36660 37420 36692
rect 37047 36626 37108 36660
rect 37154 36658 37198 36660
rect 37254 36658 37288 36660
rect 37354 36658 37378 36660
rect 37142 36626 37198 36658
rect 37232 36626 37288 36658
rect 37322 36626 37378 36658
rect 37412 36658 37420 36660
rect 37454 36660 37520 36692
rect 37454 36658 37468 36660
rect 37412 36626 37468 36658
rect 37502 36658 37520 36660
rect 37554 36660 37620 36692
rect 37654 36660 37741 36692
rect 37554 36658 37558 36660
rect 37502 36626 37558 36658
rect 37592 36658 37620 36660
rect 37592 36626 37648 36658
rect 37682 36626 37741 36660
rect 37047 36592 37741 36626
rect 37047 36570 37120 36592
rect 37154 36570 37220 36592
rect 37254 36570 37320 36592
rect 37354 36570 37420 36592
rect 37047 36536 37108 36570
rect 37154 36558 37198 36570
rect 37254 36558 37288 36570
rect 37354 36558 37378 36570
rect 37142 36536 37198 36558
rect 37232 36536 37288 36558
rect 37322 36536 37378 36558
rect 37412 36558 37420 36570
rect 37454 36570 37520 36592
rect 37454 36558 37468 36570
rect 37412 36536 37468 36558
rect 37502 36558 37520 36570
rect 37554 36570 37620 36592
rect 37654 36570 37741 36592
rect 37554 36558 37558 36570
rect 37502 36536 37558 36558
rect 37592 36558 37620 36570
rect 37592 36536 37648 36558
rect 37682 36536 37741 36570
rect 37047 36492 37741 36536
rect 37047 36480 37120 36492
rect 37154 36480 37220 36492
rect 37254 36480 37320 36492
rect 37354 36480 37420 36492
rect 37047 36446 37108 36480
rect 37154 36458 37198 36480
rect 37254 36458 37288 36480
rect 37354 36458 37378 36480
rect 37142 36446 37198 36458
rect 37232 36446 37288 36458
rect 37322 36446 37378 36458
rect 37412 36458 37420 36480
rect 37454 36480 37520 36492
rect 37454 36458 37468 36480
rect 37412 36446 37468 36458
rect 37502 36458 37520 36480
rect 37554 36480 37620 36492
rect 37654 36480 37741 36492
rect 37554 36458 37558 36480
rect 37502 36446 37558 36458
rect 37592 36458 37620 36480
rect 37592 36446 37648 36458
rect 37682 36446 37741 36480
rect 37047 36385 37741 36446
rect 37803 37028 37875 37084
rect 37803 36994 37822 37028
rect 37856 36994 37875 37028
rect 37803 36938 37875 36994
rect 37803 36904 37822 36938
rect 37856 36904 37875 36938
rect 37803 36848 37875 36904
rect 37803 36814 37822 36848
rect 37856 36814 37875 36848
rect 37803 36758 37875 36814
rect 37803 36724 37822 36758
rect 37856 36724 37875 36758
rect 37803 36668 37875 36724
rect 37803 36634 37822 36668
rect 37856 36634 37875 36668
rect 37803 36578 37875 36634
rect 37803 36544 37822 36578
rect 37856 36544 37875 36578
rect 37803 36488 37875 36544
rect 37803 36454 37822 36488
rect 37856 36454 37875 36488
rect 37803 36398 37875 36454
rect 36913 36323 36985 36383
rect 37803 36364 37822 36398
rect 37856 36364 37875 36398
rect 37803 36323 37875 36364
rect 36913 36304 37875 36323
rect 36913 36270 37010 36304
rect 37044 36270 37100 36304
rect 37134 36270 37190 36304
rect 37224 36270 37280 36304
rect 37314 36270 37370 36304
rect 37404 36270 37460 36304
rect 37494 36270 37550 36304
rect 37584 36270 37640 36304
rect 37674 36270 37730 36304
rect 37764 36270 37875 36304
rect 36913 36251 37875 36270
rect 37939 37194 37971 37228
rect 38005 37194 38124 37228
rect 38158 37194 38189 37228
rect 39279 37228 39378 37277
rect 37939 37138 38189 37194
rect 37939 37104 37971 37138
rect 38005 37104 38124 37138
rect 38158 37104 38189 37138
rect 37939 37048 38189 37104
rect 37939 37014 37971 37048
rect 38005 37014 38124 37048
rect 38158 37014 38189 37048
rect 37939 36958 38189 37014
rect 37939 36924 37971 36958
rect 38005 36924 38124 36958
rect 38158 36924 38189 36958
rect 37939 36868 38189 36924
rect 37939 36834 37971 36868
rect 38005 36834 38124 36868
rect 38158 36834 38189 36868
rect 37939 36778 38189 36834
rect 37939 36744 37971 36778
rect 38005 36744 38124 36778
rect 38158 36744 38189 36778
rect 37939 36688 38189 36744
rect 37939 36654 37971 36688
rect 38005 36654 38124 36688
rect 38158 36654 38189 36688
rect 37939 36598 38189 36654
rect 37939 36564 37971 36598
rect 38005 36564 38124 36598
rect 38158 36564 38189 36598
rect 37939 36508 38189 36564
rect 37939 36474 37971 36508
rect 38005 36474 38124 36508
rect 38158 36474 38189 36508
rect 37939 36418 38189 36474
rect 37939 36384 37971 36418
rect 38005 36384 38124 36418
rect 38158 36384 38189 36418
rect 37939 36328 38189 36384
rect 37939 36294 37971 36328
rect 38005 36294 38124 36328
rect 38158 36294 38189 36328
rect 36599 36204 36631 36238
rect 36665 36204 36784 36238
rect 36818 36204 36849 36238
rect 36599 36187 36849 36204
rect 37939 36238 38189 36294
rect 38253 37196 39215 37213
rect 38253 37162 38274 37196
rect 38308 37162 38364 37196
rect 38398 37194 38454 37196
rect 38488 37194 38544 37196
rect 38578 37194 38634 37196
rect 38668 37194 38724 37196
rect 38758 37194 38814 37196
rect 38848 37194 38904 37196
rect 38938 37194 38994 37196
rect 39028 37194 39084 37196
rect 39118 37194 39174 37196
rect 38418 37162 38454 37194
rect 38508 37162 38544 37194
rect 38598 37162 38634 37194
rect 38688 37162 38724 37194
rect 38778 37162 38814 37194
rect 38868 37162 38904 37194
rect 38958 37162 38994 37194
rect 39048 37162 39084 37194
rect 39138 37162 39174 37194
rect 39208 37162 39215 37196
rect 38253 37160 38384 37162
rect 38418 37160 38474 37162
rect 38508 37160 38564 37162
rect 38598 37160 38654 37162
rect 38688 37160 38744 37162
rect 38778 37160 38834 37162
rect 38868 37160 38924 37162
rect 38958 37160 39014 37162
rect 39048 37160 39104 37162
rect 39138 37160 39215 37162
rect 38253 37141 39215 37160
rect 38253 37137 38325 37141
rect 38253 37103 38272 37137
rect 38306 37103 38325 37137
rect 38253 37047 38325 37103
rect 39143 37118 39215 37141
rect 39143 37084 39162 37118
rect 39196 37084 39215 37118
rect 38253 37013 38272 37047
rect 38306 37013 38325 37047
rect 38253 36957 38325 37013
rect 38253 36923 38272 36957
rect 38306 36923 38325 36957
rect 38253 36867 38325 36923
rect 38253 36833 38272 36867
rect 38306 36833 38325 36867
rect 38253 36777 38325 36833
rect 38253 36743 38272 36777
rect 38306 36743 38325 36777
rect 38253 36687 38325 36743
rect 38253 36653 38272 36687
rect 38306 36653 38325 36687
rect 38253 36597 38325 36653
rect 38253 36563 38272 36597
rect 38306 36563 38325 36597
rect 38253 36507 38325 36563
rect 38253 36473 38272 36507
rect 38306 36473 38325 36507
rect 38253 36417 38325 36473
rect 38253 36383 38272 36417
rect 38306 36383 38325 36417
rect 38387 37020 39081 37079
rect 38387 36986 38448 37020
rect 38482 36992 38538 37020
rect 38572 36992 38628 37020
rect 38662 36992 38718 37020
rect 38494 36986 38538 36992
rect 38594 36986 38628 36992
rect 38694 36986 38718 36992
rect 38752 36992 38808 37020
rect 38752 36986 38760 36992
rect 38387 36958 38460 36986
rect 38494 36958 38560 36986
rect 38594 36958 38660 36986
rect 38694 36958 38760 36986
rect 38794 36986 38808 36992
rect 38842 36992 38898 37020
rect 38842 36986 38860 36992
rect 38794 36958 38860 36986
rect 38894 36986 38898 36992
rect 38932 36992 38988 37020
rect 38932 36986 38960 36992
rect 39022 36986 39081 37020
rect 38894 36958 38960 36986
rect 38994 36958 39081 36986
rect 38387 36930 39081 36958
rect 38387 36896 38448 36930
rect 38482 36896 38538 36930
rect 38572 36896 38628 36930
rect 38662 36896 38718 36930
rect 38752 36896 38808 36930
rect 38842 36896 38898 36930
rect 38932 36896 38988 36930
rect 39022 36896 39081 36930
rect 38387 36892 39081 36896
rect 38387 36858 38460 36892
rect 38494 36858 38560 36892
rect 38594 36858 38660 36892
rect 38694 36858 38760 36892
rect 38794 36858 38860 36892
rect 38894 36858 38960 36892
rect 38994 36858 39081 36892
rect 38387 36840 39081 36858
rect 38387 36806 38448 36840
rect 38482 36806 38538 36840
rect 38572 36806 38628 36840
rect 38662 36806 38718 36840
rect 38752 36806 38808 36840
rect 38842 36806 38898 36840
rect 38932 36806 38988 36840
rect 39022 36806 39081 36840
rect 38387 36792 39081 36806
rect 38387 36758 38460 36792
rect 38494 36758 38560 36792
rect 38594 36758 38660 36792
rect 38694 36758 38760 36792
rect 38794 36758 38860 36792
rect 38894 36758 38960 36792
rect 38994 36758 39081 36792
rect 38387 36750 39081 36758
rect 38387 36716 38448 36750
rect 38482 36716 38538 36750
rect 38572 36716 38628 36750
rect 38662 36716 38718 36750
rect 38752 36716 38808 36750
rect 38842 36716 38898 36750
rect 38932 36716 38988 36750
rect 39022 36716 39081 36750
rect 38387 36692 39081 36716
rect 38387 36660 38460 36692
rect 38494 36660 38560 36692
rect 38594 36660 38660 36692
rect 38694 36660 38760 36692
rect 38387 36626 38448 36660
rect 38494 36658 38538 36660
rect 38594 36658 38628 36660
rect 38694 36658 38718 36660
rect 38482 36626 38538 36658
rect 38572 36626 38628 36658
rect 38662 36626 38718 36658
rect 38752 36658 38760 36660
rect 38794 36660 38860 36692
rect 38794 36658 38808 36660
rect 38752 36626 38808 36658
rect 38842 36658 38860 36660
rect 38894 36660 38960 36692
rect 38994 36660 39081 36692
rect 38894 36658 38898 36660
rect 38842 36626 38898 36658
rect 38932 36658 38960 36660
rect 38932 36626 38988 36658
rect 39022 36626 39081 36660
rect 38387 36592 39081 36626
rect 38387 36570 38460 36592
rect 38494 36570 38560 36592
rect 38594 36570 38660 36592
rect 38694 36570 38760 36592
rect 38387 36536 38448 36570
rect 38494 36558 38538 36570
rect 38594 36558 38628 36570
rect 38694 36558 38718 36570
rect 38482 36536 38538 36558
rect 38572 36536 38628 36558
rect 38662 36536 38718 36558
rect 38752 36558 38760 36570
rect 38794 36570 38860 36592
rect 38794 36558 38808 36570
rect 38752 36536 38808 36558
rect 38842 36558 38860 36570
rect 38894 36570 38960 36592
rect 38994 36570 39081 36592
rect 38894 36558 38898 36570
rect 38842 36536 38898 36558
rect 38932 36558 38960 36570
rect 38932 36536 38988 36558
rect 39022 36536 39081 36570
rect 38387 36492 39081 36536
rect 38387 36480 38460 36492
rect 38494 36480 38560 36492
rect 38594 36480 38660 36492
rect 38694 36480 38760 36492
rect 38387 36446 38448 36480
rect 38494 36458 38538 36480
rect 38594 36458 38628 36480
rect 38694 36458 38718 36480
rect 38482 36446 38538 36458
rect 38572 36446 38628 36458
rect 38662 36446 38718 36458
rect 38752 36458 38760 36480
rect 38794 36480 38860 36492
rect 38794 36458 38808 36480
rect 38752 36446 38808 36458
rect 38842 36458 38860 36480
rect 38894 36480 38960 36492
rect 38994 36480 39081 36492
rect 38894 36458 38898 36480
rect 38842 36446 38898 36458
rect 38932 36458 38960 36480
rect 38932 36446 38988 36458
rect 39022 36446 39081 36480
rect 38387 36385 39081 36446
rect 39143 37028 39215 37084
rect 39143 36994 39162 37028
rect 39196 36994 39215 37028
rect 39143 36938 39215 36994
rect 39143 36904 39162 36938
rect 39196 36904 39215 36938
rect 39143 36848 39215 36904
rect 39143 36814 39162 36848
rect 39196 36814 39215 36848
rect 39143 36758 39215 36814
rect 39143 36724 39162 36758
rect 39196 36724 39215 36758
rect 39143 36668 39215 36724
rect 39143 36634 39162 36668
rect 39196 36634 39215 36668
rect 39143 36578 39215 36634
rect 39143 36544 39162 36578
rect 39196 36544 39215 36578
rect 39143 36488 39215 36544
rect 39143 36454 39162 36488
rect 39196 36454 39215 36488
rect 39143 36398 39215 36454
rect 38253 36323 38325 36383
rect 39143 36364 39162 36398
rect 39196 36364 39215 36398
rect 39143 36323 39215 36364
rect 38253 36304 39215 36323
rect 38253 36270 38350 36304
rect 38384 36270 38440 36304
rect 38474 36270 38530 36304
rect 38564 36270 38620 36304
rect 38654 36270 38710 36304
rect 38744 36270 38800 36304
rect 38834 36270 38890 36304
rect 38924 36270 38980 36304
rect 39014 36270 39070 36304
rect 39104 36270 39215 36304
rect 38253 36251 39215 36270
rect 39279 37194 39311 37228
rect 39345 37194 39378 37228
rect 39279 37138 39378 37194
rect 39279 37104 39311 37138
rect 39345 37104 39378 37138
rect 39279 37048 39378 37104
rect 39279 37014 39311 37048
rect 39345 37014 39378 37048
rect 39279 36958 39378 37014
rect 39279 36924 39311 36958
rect 39345 36924 39378 36958
rect 39279 36868 39378 36924
rect 39279 36834 39311 36868
rect 39345 36834 39378 36868
rect 39279 36778 39378 36834
rect 39279 36744 39311 36778
rect 39345 36744 39378 36778
rect 39279 36688 39378 36744
rect 39279 36654 39311 36688
rect 39345 36654 39378 36688
rect 39279 36598 39378 36654
rect 39279 36564 39311 36598
rect 39345 36564 39378 36598
rect 39279 36508 39378 36564
rect 39279 36474 39311 36508
rect 39345 36474 39378 36508
rect 40658 36723 41274 36762
rect 40658 36621 40745 36723
rect 41187 36621 41274 36723
rect 39279 36418 39378 36474
rect 39279 36384 39311 36418
rect 39345 36384 39378 36418
rect 39279 36328 39378 36384
rect 39279 36294 39311 36328
rect 39345 36294 39378 36328
rect 37939 36204 37971 36238
rect 38005 36204 38124 36238
rect 38158 36204 38189 36238
rect 37939 36187 38189 36204
rect 39279 36238 39378 36294
rect 39279 36204 39311 36238
rect 39345 36204 39378 36238
rect 39279 36187 39378 36204
rect 30050 36154 39378 36187
rect 30050 36120 30180 36154
rect 30214 36120 30270 36154
rect 30304 36120 30360 36154
rect 30394 36120 30450 36154
rect 30484 36120 30540 36154
rect 30574 36120 30630 36154
rect 30664 36120 30720 36154
rect 30754 36120 30810 36154
rect 30844 36120 30900 36154
rect 30934 36120 30990 36154
rect 31024 36120 31080 36154
rect 31114 36120 31170 36154
rect 31204 36120 31520 36154
rect 31554 36120 31610 36154
rect 31644 36120 31700 36154
rect 31734 36120 31790 36154
rect 31824 36120 31880 36154
rect 31914 36120 31970 36154
rect 32004 36120 32060 36154
rect 32094 36120 32150 36154
rect 32184 36120 32240 36154
rect 32274 36120 32330 36154
rect 32364 36120 32420 36154
rect 32454 36120 32510 36154
rect 32544 36120 32860 36154
rect 32894 36120 32950 36154
rect 32984 36120 33040 36154
rect 33074 36120 33130 36154
rect 33164 36120 33220 36154
rect 33254 36120 33310 36154
rect 33344 36120 33400 36154
rect 33434 36120 33490 36154
rect 33524 36120 33580 36154
rect 33614 36120 33670 36154
rect 33704 36120 33760 36154
rect 33794 36120 33850 36154
rect 33884 36120 34200 36154
rect 34234 36120 34290 36154
rect 34324 36120 34380 36154
rect 34414 36120 34470 36154
rect 34504 36120 34560 36154
rect 34594 36120 34650 36154
rect 34684 36120 34740 36154
rect 34774 36120 34830 36154
rect 34864 36120 34920 36154
rect 34954 36120 35010 36154
rect 35044 36120 35100 36154
rect 35134 36120 35190 36154
rect 35224 36120 35540 36154
rect 35574 36120 35630 36154
rect 35664 36120 35720 36154
rect 35754 36120 35810 36154
rect 35844 36120 35900 36154
rect 35934 36120 35990 36154
rect 36024 36120 36080 36154
rect 36114 36120 36170 36154
rect 36204 36120 36260 36154
rect 36294 36120 36350 36154
rect 36384 36120 36440 36154
rect 36474 36120 36530 36154
rect 36564 36120 36880 36154
rect 36914 36120 36970 36154
rect 37004 36120 37060 36154
rect 37094 36120 37150 36154
rect 37184 36120 37240 36154
rect 37274 36120 37330 36154
rect 37364 36120 37420 36154
rect 37454 36120 37510 36154
rect 37544 36120 37600 36154
rect 37634 36120 37690 36154
rect 37724 36120 37780 36154
rect 37814 36120 37870 36154
rect 37904 36120 38220 36154
rect 38254 36120 38310 36154
rect 38344 36120 38400 36154
rect 38434 36120 38490 36154
rect 38524 36120 38580 36154
rect 38614 36120 38670 36154
rect 38704 36120 38760 36154
rect 38794 36120 38850 36154
rect 38884 36120 38940 36154
rect 38974 36120 39030 36154
rect 39064 36120 39120 36154
rect 39154 36120 39210 36154
rect 39244 36120 39378 36154
rect 30050 36088 39378 36120
rect 28258 35949 28318 36032
rect 28258 35915 28271 35949
rect 28305 35915 28318 35949
rect 28408 35983 28844 35996
rect 28408 35955 28511 35983
rect 28408 35936 28457 35955
rect 28491 35949 28511 35955
rect 28545 35949 28844 35983
rect 28491 35936 28844 35949
rect 28258 35822 28318 35915
rect 40658 35822 41274 36621
rect 41754 36477 42186 36867
rect 5918 35809 13086 35822
rect 5918 35775 6101 35809
rect 6135 35775 6501 35809
rect 6535 35775 6901 35809
rect 6935 35775 7301 35809
rect 7335 35775 7701 35809
rect 7735 35775 8101 35809
rect 8135 35775 8501 35809
rect 8535 35775 8901 35809
rect 8935 35775 9301 35809
rect 9335 35775 9701 35809
rect 9735 35775 10101 35809
rect 10135 35775 10501 35809
rect 10535 35775 10901 35809
rect 10935 35775 11301 35809
rect 11335 35775 11701 35809
rect 11735 35775 12101 35809
rect 12135 35775 12501 35809
rect 12535 35775 12901 35809
rect 12935 35775 13086 35809
rect 5918 35762 13086 35775
rect 13366 35809 20534 35822
rect 13366 35775 13549 35809
rect 13583 35775 13949 35809
rect 13983 35775 14349 35809
rect 14383 35775 14749 35809
rect 14783 35775 15149 35809
rect 15183 35775 15549 35809
rect 15583 35775 15949 35809
rect 15983 35775 16349 35809
rect 16383 35775 16749 35809
rect 16783 35775 17149 35809
rect 17183 35775 17549 35809
rect 17583 35775 17949 35809
rect 17983 35775 18349 35809
rect 18383 35775 18749 35809
rect 18783 35775 19149 35809
rect 19183 35775 19549 35809
rect 19583 35775 19949 35809
rect 19983 35775 20349 35809
rect 20383 35775 20534 35809
rect 13366 35762 20534 35775
rect 20814 35809 27982 35822
rect 20814 35775 20997 35809
rect 21031 35775 21397 35809
rect 21431 35775 21797 35809
rect 21831 35775 22197 35809
rect 22231 35775 22597 35809
rect 22631 35775 22997 35809
rect 23031 35775 23397 35809
rect 23431 35775 23797 35809
rect 23831 35775 24197 35809
rect 24231 35775 24597 35809
rect 24631 35775 24997 35809
rect 25031 35775 25397 35809
rect 25431 35775 25797 35809
rect 25831 35775 26197 35809
rect 26231 35775 26597 35809
rect 26631 35775 26997 35809
rect 27031 35775 27397 35809
rect 27431 35775 27797 35809
rect 27831 35775 27982 35809
rect 20814 35762 27982 35775
rect 28230 35809 28844 35822
rect 28230 35775 28511 35809
rect 28545 35775 28844 35809
rect 28230 35762 28844 35775
rect 30024 35809 39404 35822
rect 30024 35775 30207 35809
rect 30241 35775 30407 35809
rect 30441 35775 30607 35809
rect 30641 35775 30807 35809
rect 30841 35775 31007 35809
rect 31041 35775 31207 35809
rect 31241 35775 31407 35809
rect 31441 35775 31607 35809
rect 31641 35775 31807 35809
rect 31841 35775 32007 35809
rect 32041 35775 32207 35809
rect 32241 35775 32407 35809
rect 32441 35775 32607 35809
rect 32641 35775 32807 35809
rect 32841 35775 33007 35809
rect 33041 35775 33207 35809
rect 33241 35775 33407 35809
rect 33441 35775 33607 35809
rect 33641 35775 33807 35809
rect 33841 35775 34007 35809
rect 34041 35775 34207 35809
rect 34241 35775 34407 35809
rect 34441 35775 34607 35809
rect 34641 35775 34807 35809
rect 34841 35775 35007 35809
rect 35041 35775 35207 35809
rect 35241 35775 35407 35809
rect 35441 35775 35607 35809
rect 35641 35775 35807 35809
rect 35841 35775 36007 35809
rect 36041 35775 36207 35809
rect 36241 35775 36407 35809
rect 36441 35775 36607 35809
rect 36641 35775 36807 35809
rect 36841 35775 37007 35809
rect 37041 35775 37207 35809
rect 37241 35775 37407 35809
rect 37441 35775 37607 35809
rect 37641 35775 37807 35809
rect 37841 35775 38007 35809
rect 38041 35775 38207 35809
rect 38241 35775 38407 35809
rect 38441 35775 38607 35809
rect 38641 35775 38807 35809
rect 38841 35775 39007 35809
rect 39041 35775 39207 35809
rect 39241 35775 39404 35809
rect 30024 35762 39404 35775
rect 39746 35809 42186 35822
rect 39746 35775 39929 35809
rect 39963 35775 40129 35809
rect 40163 35775 40329 35809
rect 40363 35775 40529 35809
rect 40563 35775 40729 35809
rect 40763 35775 40929 35809
rect 40963 35775 41129 35809
rect 41163 35775 41329 35809
rect 41363 35775 41529 35809
rect 41563 35775 41729 35809
rect 41763 35775 41929 35809
rect 41963 35775 42186 35809
rect 39746 35762 42186 35775
rect 6604 33929 13772 33942
rect 6604 33895 6787 33929
rect 6821 33895 7187 33929
rect 7221 33895 7587 33929
rect 7621 33895 7987 33929
rect 8021 33895 8387 33929
rect 8421 33895 8787 33929
rect 8821 33895 9187 33929
rect 9221 33895 9587 33929
rect 9621 33895 9987 33929
rect 10021 33895 10387 33929
rect 10421 33895 10787 33929
rect 10821 33895 11187 33929
rect 11221 33895 11587 33929
rect 11621 33895 11987 33929
rect 12021 33895 12387 33929
rect 12421 33895 12787 33929
rect 12821 33895 13187 33929
rect 13221 33895 13587 33929
rect 13621 33895 13772 33929
rect 6604 33882 13772 33895
rect 14050 33929 41756 33942
rect 14050 33895 14331 33929
rect 14365 33895 14731 33929
rect 14765 33895 15131 33929
rect 15165 33895 15531 33929
rect 15565 33895 15931 33929
rect 15965 33895 16331 33929
rect 16365 33895 16731 33929
rect 16765 33895 17131 33929
rect 17165 33895 17531 33929
rect 17565 33895 17931 33929
rect 17965 33895 18331 33929
rect 18365 33895 18731 33929
rect 18765 33895 19131 33929
rect 19165 33895 19531 33929
rect 19565 33895 19931 33929
rect 19965 33895 20331 33929
rect 20365 33895 20731 33929
rect 20765 33895 21131 33929
rect 21165 33895 21531 33929
rect 21565 33895 21931 33929
rect 21965 33895 22331 33929
rect 22365 33895 22731 33929
rect 22765 33895 23131 33929
rect 23165 33895 23531 33929
rect 23565 33895 23931 33929
rect 23965 33895 24331 33929
rect 24365 33895 24731 33929
rect 24765 33895 25131 33929
rect 25165 33895 25531 33929
rect 25565 33895 25931 33929
rect 25965 33895 26331 33929
rect 26365 33895 26731 33929
rect 26765 33895 27131 33929
rect 27165 33895 27531 33929
rect 27565 33895 27931 33929
rect 27965 33895 28331 33929
rect 28365 33895 28731 33929
rect 28765 33895 29131 33929
rect 29165 33895 29531 33929
rect 29565 33895 29931 33929
rect 29965 33895 30331 33929
rect 30365 33895 30731 33929
rect 30765 33895 31131 33929
rect 31165 33895 31531 33929
rect 31565 33895 31931 33929
rect 31965 33895 32331 33929
rect 32365 33895 32731 33929
rect 32765 33895 33131 33929
rect 33165 33895 33531 33929
rect 33565 33895 33931 33929
rect 33965 33895 34331 33929
rect 34365 33895 34731 33929
rect 34765 33895 35131 33929
rect 35165 33895 35531 33929
rect 35565 33895 35931 33929
rect 35965 33895 36331 33929
rect 36365 33895 36731 33929
rect 36765 33895 37131 33929
rect 37165 33895 37531 33929
rect 37565 33895 37931 33929
rect 37965 33895 38331 33929
rect 38365 33895 38731 33929
rect 38765 33895 39131 33929
rect 39165 33895 39531 33929
rect 39565 33895 39931 33929
rect 39965 33895 40331 33929
rect 40365 33895 40731 33929
rect 40765 33895 41131 33929
rect 41165 33895 41531 33929
rect 41565 33895 41756 33929
rect 14050 33882 41756 33895
rect 14078 33789 14138 33882
rect 15126 33839 15286 33882
rect 15126 33805 15191 33839
rect 15225 33805 15286 33839
rect 15126 33802 15286 33805
rect 16426 33839 16586 33882
rect 16426 33805 16491 33839
rect 16525 33805 16586 33839
rect 16426 33802 16586 33805
rect 17726 33839 17886 33882
rect 17726 33805 17791 33839
rect 17825 33805 17886 33839
rect 17726 33802 17886 33805
rect 19026 33839 19186 33882
rect 19026 33805 19091 33839
rect 19125 33805 19186 33839
rect 19026 33802 19186 33805
rect 20326 33839 20486 33882
rect 20326 33805 20391 33839
rect 20425 33805 20486 33839
rect 20326 33802 20486 33805
rect 21626 33839 21786 33882
rect 21626 33805 21691 33839
rect 21725 33805 21786 33839
rect 21626 33802 21786 33805
rect 22926 33839 23086 33882
rect 22926 33805 22991 33839
rect 23025 33805 23086 33839
rect 22926 33802 23086 33805
rect 24226 33839 24386 33882
rect 24226 33805 24291 33839
rect 24325 33805 24386 33839
rect 24226 33802 24386 33805
rect 25526 33839 25686 33882
rect 25526 33805 25591 33839
rect 25625 33805 25686 33839
rect 25526 33802 25686 33805
rect 26826 33839 26986 33882
rect 26826 33805 26891 33839
rect 26925 33805 26986 33839
rect 26826 33802 26986 33805
rect 28126 33839 28286 33882
rect 28126 33805 28191 33839
rect 28225 33805 28286 33839
rect 28126 33802 28286 33805
rect 29426 33839 29586 33882
rect 29426 33805 29491 33839
rect 29525 33805 29586 33839
rect 29426 33802 29586 33805
rect 30726 33839 30886 33882
rect 30726 33805 30791 33839
rect 30825 33805 30886 33839
rect 30726 33802 30886 33805
rect 32026 33839 32186 33882
rect 32026 33805 32091 33839
rect 32125 33805 32186 33839
rect 32026 33802 32186 33805
rect 33326 33839 33486 33882
rect 33326 33805 33391 33839
rect 33425 33805 33486 33839
rect 33326 33802 33486 33805
rect 34626 33839 34786 33882
rect 34626 33805 34691 33839
rect 34725 33805 34786 33839
rect 34626 33802 34786 33805
rect 35926 33839 36086 33882
rect 35926 33805 35991 33839
rect 36025 33805 36086 33839
rect 35926 33802 36086 33805
rect 37226 33839 37386 33882
rect 37226 33805 37291 33839
rect 37325 33805 37386 33839
rect 37226 33802 37386 33805
rect 38526 33839 38686 33882
rect 38526 33805 38591 33839
rect 38625 33805 38686 33839
rect 38526 33802 38686 33805
rect 39826 33839 39986 33882
rect 39826 33805 39891 33839
rect 39925 33805 39986 33839
rect 39826 33802 39986 33805
rect 14078 33755 14091 33789
rect 14125 33755 14138 33789
rect 14078 33672 14138 33755
rect 14208 33722 41756 33762
rect 14195 33661 14229 33681
rect 14195 33593 14229 33627
rect 14195 33525 14229 33555
rect 14195 33457 14229 33483
rect 14195 33389 14229 33411
rect 14195 33321 14229 33339
rect 14195 33253 14229 33267
rect 14195 33185 14229 33195
rect 14195 33117 14229 33123
rect 14195 33049 14229 33051
rect 14195 33013 14229 33015
rect 14195 32941 14229 32947
rect 14195 32869 14229 32879
rect 14195 32797 14229 32811
rect 14195 32725 14229 32743
rect 14195 32653 14229 32675
rect 14195 32581 14229 32607
rect 14195 32509 14229 32539
rect 14195 32437 14229 32471
rect 14195 32302 14229 32403
rect 14653 33661 14687 33722
rect 14653 33593 14687 33627
rect 14653 33525 14687 33555
rect 14653 33457 14687 33483
rect 14653 33389 14687 33411
rect 14653 33321 14687 33339
rect 14653 33253 14687 33267
rect 14653 33185 14687 33195
rect 14653 33117 14687 33123
rect 14653 33049 14687 33051
rect 14653 33013 14687 33015
rect 14653 32941 14687 32947
rect 14653 32869 14687 32879
rect 14653 32797 14687 32811
rect 14653 32725 14687 32743
rect 14653 32653 14687 32675
rect 14653 32581 14687 32607
rect 14653 32509 14687 32539
rect 14653 32437 14687 32471
rect 14653 32383 14687 32403
rect 15111 33661 15145 33681
rect 15111 33593 15145 33627
rect 15111 33525 15145 33555
rect 15111 33457 15145 33483
rect 15111 33389 15145 33411
rect 15111 33321 15145 33339
rect 15111 33253 15145 33267
rect 15111 33185 15145 33195
rect 15111 33117 15145 33123
rect 15111 33049 15145 33051
rect 15111 33013 15145 33015
rect 15111 32941 15145 32947
rect 15111 32869 15145 32879
rect 15111 32797 15145 32811
rect 15111 32725 15145 32743
rect 15111 32653 15145 32675
rect 15111 32581 15145 32607
rect 15111 32509 15145 32539
rect 15111 32437 15145 32471
rect 15111 32302 15145 32403
rect 15569 33661 15603 33722
rect 15569 33593 15603 33627
rect 15569 33525 15603 33555
rect 15569 33457 15603 33483
rect 15569 33389 15603 33411
rect 15569 33321 15603 33339
rect 15569 33253 15603 33267
rect 15569 33185 15603 33195
rect 15569 33117 15603 33123
rect 15569 33049 15603 33051
rect 15569 33013 15603 33015
rect 15569 32941 15603 32947
rect 15569 32869 15603 32879
rect 15569 32797 15603 32811
rect 15569 32725 15603 32743
rect 15569 32653 15603 32675
rect 15569 32581 15603 32607
rect 15569 32509 15603 32539
rect 15569 32437 15603 32471
rect 15569 32383 15603 32403
rect 16027 33661 16061 33681
rect 16027 33593 16061 33627
rect 16027 33525 16061 33555
rect 16027 33457 16061 33483
rect 16027 33389 16061 33411
rect 16027 33321 16061 33339
rect 16027 33253 16061 33267
rect 16027 33185 16061 33195
rect 16027 33117 16061 33123
rect 16027 33049 16061 33051
rect 16027 33013 16061 33015
rect 16027 32941 16061 32947
rect 16027 32869 16061 32879
rect 16027 32797 16061 32811
rect 16027 32725 16061 32743
rect 16027 32653 16061 32675
rect 16027 32581 16061 32607
rect 16027 32509 16061 32539
rect 16027 32437 16061 32471
rect 16027 32302 16061 32403
rect 16485 33661 16519 33722
rect 16485 33593 16519 33627
rect 16485 33525 16519 33555
rect 16485 33457 16519 33483
rect 16485 33389 16519 33411
rect 16485 33321 16519 33339
rect 16485 33253 16519 33267
rect 16485 33185 16519 33195
rect 16485 33117 16519 33123
rect 16485 33049 16519 33051
rect 16485 33013 16519 33015
rect 16485 32941 16519 32947
rect 16485 32869 16519 32879
rect 16485 32797 16519 32811
rect 16485 32725 16519 32743
rect 16485 32653 16519 32675
rect 16485 32581 16519 32607
rect 16485 32509 16519 32539
rect 16485 32437 16519 32471
rect 16485 32383 16519 32403
rect 16943 33661 16977 33681
rect 16943 33593 16977 33627
rect 16943 33525 16977 33555
rect 16943 33457 16977 33483
rect 16943 33389 16977 33411
rect 16943 33321 16977 33339
rect 16943 33253 16977 33267
rect 16943 33185 16977 33195
rect 16943 33117 16977 33123
rect 16943 33049 16977 33051
rect 16943 33013 16977 33015
rect 16943 32941 16977 32947
rect 16943 32869 16977 32879
rect 16943 32797 16977 32811
rect 16943 32725 16977 32743
rect 16943 32653 16977 32675
rect 16943 32581 16977 32607
rect 16943 32509 16977 32539
rect 16943 32437 16977 32471
rect 16943 32302 16977 32403
rect 17401 33661 17435 33722
rect 17401 33593 17435 33627
rect 17401 33525 17435 33555
rect 17401 33457 17435 33483
rect 17401 33389 17435 33411
rect 17401 33321 17435 33339
rect 17401 33253 17435 33267
rect 17401 33185 17435 33195
rect 17401 33117 17435 33123
rect 17401 33049 17435 33051
rect 17401 33013 17435 33015
rect 17401 32941 17435 32947
rect 17401 32869 17435 32879
rect 17401 32797 17435 32811
rect 17401 32725 17435 32743
rect 17401 32653 17435 32675
rect 17401 32581 17435 32607
rect 17401 32509 17435 32539
rect 17401 32437 17435 32471
rect 17401 32383 17435 32403
rect 17859 33661 17893 33681
rect 17859 33593 17893 33627
rect 17859 33525 17893 33555
rect 17859 33457 17893 33483
rect 17859 33389 17893 33411
rect 17859 33321 17893 33339
rect 17859 33253 17893 33267
rect 17859 33185 17893 33195
rect 17859 33117 17893 33123
rect 17859 33049 17893 33051
rect 17859 33013 17893 33015
rect 17859 32941 17893 32947
rect 17859 32869 17893 32879
rect 17859 32797 17893 32811
rect 17859 32725 17893 32743
rect 17859 32653 17893 32675
rect 17859 32581 17893 32607
rect 17859 32509 17893 32539
rect 17859 32437 17893 32471
rect 17859 32302 17893 32403
rect 18317 33661 18351 33722
rect 18317 33593 18351 33627
rect 18317 33525 18351 33555
rect 18317 33457 18351 33483
rect 18317 33389 18351 33411
rect 18317 33321 18351 33339
rect 18317 33253 18351 33267
rect 18317 33185 18351 33195
rect 18317 33117 18351 33123
rect 18317 33049 18351 33051
rect 18317 33013 18351 33015
rect 18317 32941 18351 32947
rect 18317 32869 18351 32879
rect 18317 32797 18351 32811
rect 18317 32725 18351 32743
rect 18317 32653 18351 32675
rect 18317 32581 18351 32607
rect 18317 32509 18351 32539
rect 18317 32437 18351 32471
rect 18317 32383 18351 32403
rect 18775 33661 18809 33681
rect 18775 33593 18809 33627
rect 18775 33525 18809 33555
rect 18775 33457 18809 33483
rect 18775 33389 18809 33411
rect 18775 33321 18809 33339
rect 18775 33253 18809 33267
rect 18775 33185 18809 33195
rect 18775 33117 18809 33123
rect 18775 33049 18809 33051
rect 18775 33013 18809 33015
rect 18775 32941 18809 32947
rect 18775 32869 18809 32879
rect 18775 32797 18809 32811
rect 18775 32725 18809 32743
rect 18775 32653 18809 32675
rect 18775 32581 18809 32607
rect 18775 32509 18809 32539
rect 18775 32437 18809 32471
rect 18775 32302 18809 32403
rect 19233 33661 19267 33722
rect 19233 33593 19267 33627
rect 19233 33525 19267 33555
rect 19233 33457 19267 33483
rect 19233 33389 19267 33411
rect 19233 33321 19267 33339
rect 19233 33253 19267 33267
rect 19233 33185 19267 33195
rect 19233 33117 19267 33123
rect 19233 33049 19267 33051
rect 19233 33013 19267 33015
rect 19233 32941 19267 32947
rect 19233 32869 19267 32879
rect 19233 32797 19267 32811
rect 19233 32725 19267 32743
rect 19233 32653 19267 32675
rect 19233 32581 19267 32607
rect 19233 32509 19267 32539
rect 19233 32437 19267 32471
rect 19233 32383 19267 32403
rect 19691 33661 19725 33681
rect 19691 33593 19725 33627
rect 19691 33525 19725 33555
rect 19691 33457 19725 33483
rect 19691 33389 19725 33411
rect 19691 33321 19725 33339
rect 19691 33253 19725 33267
rect 19691 33185 19725 33195
rect 19691 33117 19725 33123
rect 19691 33049 19725 33051
rect 19691 33013 19725 33015
rect 19691 32941 19725 32947
rect 19691 32869 19725 32879
rect 19691 32797 19725 32811
rect 19691 32725 19725 32743
rect 19691 32653 19725 32675
rect 19691 32581 19725 32607
rect 19691 32509 19725 32539
rect 19691 32437 19725 32471
rect 19691 32302 19725 32403
rect 20149 33661 20183 33722
rect 20149 33593 20183 33627
rect 20149 33525 20183 33555
rect 20149 33457 20183 33483
rect 20149 33389 20183 33411
rect 20149 33321 20183 33339
rect 20149 33253 20183 33267
rect 20149 33185 20183 33195
rect 20149 33117 20183 33123
rect 20149 33049 20183 33051
rect 20149 33013 20183 33015
rect 20149 32941 20183 32947
rect 20149 32869 20183 32879
rect 20149 32797 20183 32811
rect 20149 32725 20183 32743
rect 20149 32653 20183 32675
rect 20149 32581 20183 32607
rect 20149 32509 20183 32539
rect 20149 32437 20183 32471
rect 20149 32383 20183 32403
rect 20607 33661 20641 33681
rect 20607 33593 20641 33627
rect 20607 33525 20641 33555
rect 20607 33457 20641 33483
rect 20607 33389 20641 33411
rect 20607 33321 20641 33339
rect 20607 33253 20641 33267
rect 20607 33185 20641 33195
rect 20607 33117 20641 33123
rect 20607 33049 20641 33051
rect 20607 33013 20641 33015
rect 20607 32941 20641 32947
rect 20607 32869 20641 32879
rect 20607 32797 20641 32811
rect 20607 32725 20641 32743
rect 20607 32653 20641 32675
rect 20607 32581 20641 32607
rect 20607 32509 20641 32539
rect 20607 32437 20641 32471
rect 20607 32302 20641 32403
rect 21065 33661 21099 33722
rect 21065 33593 21099 33627
rect 21065 33525 21099 33555
rect 21065 33457 21099 33483
rect 21065 33389 21099 33411
rect 21065 33321 21099 33339
rect 21065 33253 21099 33267
rect 21065 33185 21099 33195
rect 21065 33117 21099 33123
rect 21065 33049 21099 33051
rect 21065 33013 21099 33015
rect 21065 32941 21099 32947
rect 21065 32869 21099 32879
rect 21065 32797 21099 32811
rect 21065 32725 21099 32743
rect 21065 32653 21099 32675
rect 21065 32581 21099 32607
rect 21065 32509 21099 32539
rect 21065 32437 21099 32471
rect 21065 32383 21099 32403
rect 21523 33661 21557 33681
rect 21523 33593 21557 33627
rect 21523 33525 21557 33555
rect 21523 33457 21557 33483
rect 21523 33389 21557 33411
rect 21523 33321 21557 33339
rect 21523 33253 21557 33267
rect 21523 33185 21557 33195
rect 21523 33117 21557 33123
rect 21523 33049 21557 33051
rect 21523 33013 21557 33015
rect 21523 32941 21557 32947
rect 21523 32869 21557 32879
rect 21523 32797 21557 32811
rect 21523 32725 21557 32743
rect 21523 32653 21557 32675
rect 21523 32581 21557 32607
rect 21523 32509 21557 32539
rect 21523 32437 21557 32471
rect 21523 32302 21557 32403
rect 21981 33661 22015 33722
rect 21981 33593 22015 33627
rect 21981 33525 22015 33555
rect 21981 33457 22015 33483
rect 21981 33389 22015 33411
rect 21981 33321 22015 33339
rect 21981 33253 22015 33267
rect 21981 33185 22015 33195
rect 21981 33117 22015 33123
rect 21981 33049 22015 33051
rect 21981 33013 22015 33015
rect 21981 32941 22015 32947
rect 21981 32869 22015 32879
rect 21981 32797 22015 32811
rect 21981 32725 22015 32743
rect 21981 32653 22015 32675
rect 21981 32581 22015 32607
rect 21981 32509 22015 32539
rect 21981 32437 22015 32471
rect 21981 32383 22015 32403
rect 22439 33661 22473 33681
rect 22439 33593 22473 33627
rect 22439 33525 22473 33555
rect 22439 33457 22473 33483
rect 22439 33389 22473 33411
rect 22439 33321 22473 33339
rect 22439 33253 22473 33267
rect 22439 33185 22473 33195
rect 22439 33117 22473 33123
rect 22439 33049 22473 33051
rect 22439 33013 22473 33015
rect 22439 32941 22473 32947
rect 22439 32869 22473 32879
rect 22439 32797 22473 32811
rect 22439 32725 22473 32743
rect 22439 32653 22473 32675
rect 22439 32581 22473 32607
rect 22439 32509 22473 32539
rect 22439 32437 22473 32471
rect 22439 32302 22473 32403
rect 22897 33661 22931 33722
rect 22897 33593 22931 33627
rect 22897 33525 22931 33555
rect 22897 33457 22931 33483
rect 22897 33389 22931 33411
rect 22897 33321 22931 33339
rect 22897 33253 22931 33267
rect 22897 33185 22931 33195
rect 22897 33117 22931 33123
rect 22897 33049 22931 33051
rect 22897 33013 22931 33015
rect 22897 32941 22931 32947
rect 22897 32869 22931 32879
rect 22897 32797 22931 32811
rect 22897 32725 22931 32743
rect 22897 32653 22931 32675
rect 22897 32581 22931 32607
rect 22897 32509 22931 32539
rect 22897 32437 22931 32471
rect 22897 32383 22931 32403
rect 23355 33661 23389 33681
rect 23355 33593 23389 33627
rect 23355 33525 23389 33555
rect 23355 33457 23389 33483
rect 23355 33389 23389 33411
rect 23355 33321 23389 33339
rect 23355 33253 23389 33267
rect 23355 33185 23389 33195
rect 23355 33117 23389 33123
rect 23355 33049 23389 33051
rect 23355 33013 23389 33015
rect 23355 32941 23389 32947
rect 23355 32869 23389 32879
rect 23355 32797 23389 32811
rect 23355 32725 23389 32743
rect 23355 32653 23389 32675
rect 23355 32581 23389 32607
rect 23355 32509 23389 32539
rect 23355 32437 23389 32471
rect 23355 32302 23389 32403
rect 23813 33661 23847 33722
rect 23813 33593 23847 33627
rect 23813 33525 23847 33555
rect 23813 33457 23847 33483
rect 23813 33389 23847 33411
rect 23813 33321 23847 33339
rect 23813 33253 23847 33267
rect 23813 33185 23847 33195
rect 23813 33117 23847 33123
rect 23813 33049 23847 33051
rect 23813 33013 23847 33015
rect 23813 32941 23847 32947
rect 23813 32869 23847 32879
rect 23813 32797 23847 32811
rect 23813 32725 23847 32743
rect 23813 32653 23847 32675
rect 23813 32581 23847 32607
rect 23813 32509 23847 32539
rect 23813 32437 23847 32471
rect 23813 32383 23847 32403
rect 24271 33661 24305 33681
rect 24271 33593 24305 33627
rect 24271 33525 24305 33555
rect 24271 33457 24305 33483
rect 24271 33389 24305 33411
rect 24271 33321 24305 33339
rect 24271 33253 24305 33267
rect 24271 33185 24305 33195
rect 24271 33117 24305 33123
rect 24271 33049 24305 33051
rect 24271 33013 24305 33015
rect 24271 32941 24305 32947
rect 24271 32869 24305 32879
rect 24271 32797 24305 32811
rect 24271 32725 24305 32743
rect 24271 32653 24305 32675
rect 24271 32581 24305 32607
rect 24271 32509 24305 32539
rect 24271 32437 24305 32471
rect 24271 32302 24305 32403
rect 24729 33661 24763 33722
rect 24729 33593 24763 33627
rect 24729 33525 24763 33555
rect 24729 33457 24763 33483
rect 24729 33389 24763 33411
rect 24729 33321 24763 33339
rect 24729 33253 24763 33267
rect 24729 33185 24763 33195
rect 24729 33117 24763 33123
rect 24729 33049 24763 33051
rect 24729 33013 24763 33015
rect 24729 32941 24763 32947
rect 24729 32869 24763 32879
rect 24729 32797 24763 32811
rect 24729 32725 24763 32743
rect 24729 32653 24763 32675
rect 24729 32581 24763 32607
rect 24729 32509 24763 32539
rect 24729 32437 24763 32471
rect 24729 32383 24763 32403
rect 25187 33661 25221 33681
rect 25187 33593 25221 33627
rect 25187 33525 25221 33555
rect 25187 33457 25221 33483
rect 25187 33389 25221 33411
rect 25187 33321 25221 33339
rect 25187 33253 25221 33267
rect 25187 33185 25221 33195
rect 25187 33117 25221 33123
rect 25187 33049 25221 33051
rect 25187 33013 25221 33015
rect 25187 32941 25221 32947
rect 25187 32869 25221 32879
rect 25187 32797 25221 32811
rect 25187 32725 25221 32743
rect 25187 32653 25221 32675
rect 25187 32581 25221 32607
rect 25187 32509 25221 32539
rect 25187 32437 25221 32471
rect 25187 32302 25221 32403
rect 25645 33661 25679 33722
rect 25645 33593 25679 33627
rect 25645 33525 25679 33555
rect 25645 33457 25679 33483
rect 25645 33389 25679 33411
rect 25645 33321 25679 33339
rect 25645 33253 25679 33267
rect 25645 33185 25679 33195
rect 25645 33117 25679 33123
rect 25645 33049 25679 33051
rect 25645 33013 25679 33015
rect 25645 32941 25679 32947
rect 25645 32869 25679 32879
rect 25645 32797 25679 32811
rect 25645 32725 25679 32743
rect 25645 32653 25679 32675
rect 25645 32581 25679 32607
rect 25645 32509 25679 32539
rect 25645 32437 25679 32471
rect 25645 32383 25679 32403
rect 26103 33661 26137 33681
rect 26103 33593 26137 33627
rect 26103 33525 26137 33555
rect 26103 33457 26137 33483
rect 26103 33389 26137 33411
rect 26103 33321 26137 33339
rect 26103 33253 26137 33267
rect 26103 33185 26137 33195
rect 26103 33117 26137 33123
rect 26103 33049 26137 33051
rect 26103 33013 26137 33015
rect 26103 32941 26137 32947
rect 26103 32869 26137 32879
rect 26103 32797 26137 32811
rect 26103 32725 26137 32743
rect 26103 32653 26137 32675
rect 26103 32581 26137 32607
rect 26103 32509 26137 32539
rect 26103 32437 26137 32471
rect 26103 32302 26137 32403
rect 26561 33661 26595 33722
rect 26561 33593 26595 33627
rect 26561 33525 26595 33555
rect 26561 33457 26595 33483
rect 26561 33389 26595 33411
rect 26561 33321 26595 33339
rect 26561 33253 26595 33267
rect 26561 33185 26595 33195
rect 26561 33117 26595 33123
rect 26561 33049 26595 33051
rect 26561 33013 26595 33015
rect 26561 32941 26595 32947
rect 26561 32869 26595 32879
rect 26561 32797 26595 32811
rect 26561 32725 26595 32743
rect 26561 32653 26595 32675
rect 26561 32581 26595 32607
rect 26561 32509 26595 32539
rect 26561 32437 26595 32471
rect 26561 32383 26595 32403
rect 27019 33661 27053 33681
rect 27019 33593 27053 33627
rect 27019 33525 27053 33555
rect 27019 33457 27053 33483
rect 27019 33389 27053 33411
rect 27019 33321 27053 33339
rect 27019 33253 27053 33267
rect 27019 33185 27053 33195
rect 27019 33117 27053 33123
rect 27019 33049 27053 33051
rect 27019 33013 27053 33015
rect 27019 32941 27053 32947
rect 27019 32869 27053 32879
rect 27019 32797 27053 32811
rect 27019 32725 27053 32743
rect 27019 32653 27053 32675
rect 27019 32581 27053 32607
rect 27019 32509 27053 32539
rect 27019 32437 27053 32471
rect 27019 32302 27053 32403
rect 27477 33661 27511 33722
rect 27477 33593 27511 33627
rect 27477 33525 27511 33555
rect 27477 33457 27511 33483
rect 27477 33389 27511 33411
rect 27477 33321 27511 33339
rect 27477 33253 27511 33267
rect 27477 33185 27511 33195
rect 27477 33117 27511 33123
rect 27477 33049 27511 33051
rect 27477 33013 27511 33015
rect 27477 32941 27511 32947
rect 27477 32869 27511 32879
rect 27477 32797 27511 32811
rect 27477 32725 27511 32743
rect 27477 32653 27511 32675
rect 27477 32581 27511 32607
rect 27477 32509 27511 32539
rect 27477 32437 27511 32471
rect 27477 32383 27511 32403
rect 27935 33661 27969 33681
rect 27935 33593 27969 33627
rect 27935 33525 27969 33555
rect 27935 33457 27969 33483
rect 27935 33389 27969 33411
rect 27935 33321 27969 33339
rect 27935 33253 27969 33267
rect 27935 33185 27969 33195
rect 27935 33117 27969 33123
rect 27935 33049 27969 33051
rect 27935 33013 27969 33015
rect 27935 32941 27969 32947
rect 27935 32869 27969 32879
rect 27935 32797 27969 32811
rect 27935 32725 27969 32743
rect 27935 32653 27969 32675
rect 27935 32581 27969 32607
rect 27935 32509 27969 32539
rect 27935 32437 27969 32471
rect 27935 32302 27969 32403
rect 28393 33661 28427 33722
rect 28393 33593 28427 33627
rect 28393 33525 28427 33555
rect 28393 33457 28427 33483
rect 28393 33389 28427 33411
rect 28393 33321 28427 33339
rect 28393 33253 28427 33267
rect 28393 33185 28427 33195
rect 28393 33117 28427 33123
rect 28393 33049 28427 33051
rect 28393 33013 28427 33015
rect 28393 32941 28427 32947
rect 28393 32869 28427 32879
rect 28393 32797 28427 32811
rect 28393 32725 28427 32743
rect 28393 32653 28427 32675
rect 28393 32581 28427 32607
rect 28393 32509 28427 32539
rect 28393 32437 28427 32471
rect 28393 32383 28427 32403
rect 28851 33661 28885 33681
rect 28851 33593 28885 33627
rect 28851 33525 28885 33555
rect 28851 33457 28885 33483
rect 28851 33389 28885 33411
rect 28851 33321 28885 33339
rect 28851 33253 28885 33267
rect 28851 33185 28885 33195
rect 28851 33117 28885 33123
rect 28851 33049 28885 33051
rect 28851 33013 28885 33015
rect 28851 32941 28885 32947
rect 28851 32869 28885 32879
rect 28851 32797 28885 32811
rect 28851 32725 28885 32743
rect 28851 32653 28885 32675
rect 28851 32581 28885 32607
rect 28851 32509 28885 32539
rect 28851 32437 28885 32471
rect 28851 32302 28885 32403
rect 29309 33661 29343 33722
rect 29309 33593 29343 33627
rect 29309 33525 29343 33555
rect 29309 33457 29343 33483
rect 29309 33389 29343 33411
rect 29309 33321 29343 33339
rect 29309 33253 29343 33267
rect 29309 33185 29343 33195
rect 29309 33117 29343 33123
rect 29309 33049 29343 33051
rect 29309 33013 29343 33015
rect 29309 32941 29343 32947
rect 29309 32869 29343 32879
rect 29309 32797 29343 32811
rect 29309 32725 29343 32743
rect 29309 32653 29343 32675
rect 29309 32581 29343 32607
rect 29309 32509 29343 32539
rect 29309 32437 29343 32471
rect 29309 32383 29343 32403
rect 29767 33661 29801 33681
rect 29767 33593 29801 33627
rect 29767 33525 29801 33555
rect 29767 33457 29801 33483
rect 29767 33389 29801 33411
rect 29767 33321 29801 33339
rect 29767 33253 29801 33267
rect 29767 33185 29801 33195
rect 29767 33117 29801 33123
rect 29767 33049 29801 33051
rect 29767 33013 29801 33015
rect 29767 32941 29801 32947
rect 29767 32869 29801 32879
rect 29767 32797 29801 32811
rect 29767 32725 29801 32743
rect 29767 32653 29801 32675
rect 29767 32581 29801 32607
rect 29767 32509 29801 32539
rect 29767 32437 29801 32471
rect 29767 32302 29801 32403
rect 30225 33661 30259 33722
rect 30225 33593 30259 33627
rect 30225 33525 30259 33555
rect 30225 33457 30259 33483
rect 30225 33389 30259 33411
rect 30225 33321 30259 33339
rect 30225 33253 30259 33267
rect 30225 33185 30259 33195
rect 30225 33117 30259 33123
rect 30225 33049 30259 33051
rect 30225 33013 30259 33015
rect 30225 32941 30259 32947
rect 30225 32869 30259 32879
rect 30225 32797 30259 32811
rect 30225 32725 30259 32743
rect 30225 32653 30259 32675
rect 30225 32581 30259 32607
rect 30225 32509 30259 32539
rect 30225 32437 30259 32471
rect 30225 32383 30259 32403
rect 30683 33661 30717 33681
rect 30683 33593 30717 33627
rect 30683 33525 30717 33555
rect 30683 33457 30717 33483
rect 30683 33389 30717 33411
rect 30683 33321 30717 33339
rect 30683 33253 30717 33267
rect 30683 33185 30717 33195
rect 30683 33117 30717 33123
rect 30683 33049 30717 33051
rect 30683 33013 30717 33015
rect 30683 32941 30717 32947
rect 30683 32869 30717 32879
rect 30683 32797 30717 32811
rect 30683 32725 30717 32743
rect 30683 32653 30717 32675
rect 30683 32581 30717 32607
rect 30683 32509 30717 32539
rect 30683 32437 30717 32471
rect 30683 32302 30717 32403
rect 31141 33661 31175 33722
rect 31141 33593 31175 33627
rect 31141 33525 31175 33555
rect 31141 33457 31175 33483
rect 31141 33389 31175 33411
rect 31141 33321 31175 33339
rect 31141 33253 31175 33267
rect 31141 33185 31175 33195
rect 31141 33117 31175 33123
rect 31141 33049 31175 33051
rect 31141 33013 31175 33015
rect 31141 32941 31175 32947
rect 31141 32869 31175 32879
rect 31141 32797 31175 32811
rect 31141 32725 31175 32743
rect 31141 32653 31175 32675
rect 31141 32581 31175 32607
rect 31141 32509 31175 32539
rect 31141 32437 31175 32471
rect 31141 32383 31175 32403
rect 31599 33661 31633 33681
rect 31599 33593 31633 33627
rect 31599 33525 31633 33555
rect 31599 33457 31633 33483
rect 31599 33389 31633 33411
rect 31599 33321 31633 33339
rect 31599 33253 31633 33267
rect 31599 33185 31633 33195
rect 31599 33117 31633 33123
rect 31599 33049 31633 33051
rect 31599 33013 31633 33015
rect 31599 32941 31633 32947
rect 31599 32869 31633 32879
rect 31599 32797 31633 32811
rect 31599 32725 31633 32743
rect 31599 32653 31633 32675
rect 31599 32581 31633 32607
rect 31599 32509 31633 32539
rect 31599 32437 31633 32471
rect 31599 32302 31633 32403
rect 32057 33661 32091 33722
rect 32057 33593 32091 33627
rect 32057 33525 32091 33555
rect 32057 33457 32091 33483
rect 32057 33389 32091 33411
rect 32057 33321 32091 33339
rect 32057 33253 32091 33267
rect 32057 33185 32091 33195
rect 32057 33117 32091 33123
rect 32057 33049 32091 33051
rect 32057 33013 32091 33015
rect 32057 32941 32091 32947
rect 32057 32869 32091 32879
rect 32057 32797 32091 32811
rect 32057 32725 32091 32743
rect 32057 32653 32091 32675
rect 32057 32581 32091 32607
rect 32057 32509 32091 32539
rect 32057 32437 32091 32471
rect 32057 32383 32091 32403
rect 32515 33661 32549 33681
rect 32515 33593 32549 33627
rect 32515 33525 32549 33555
rect 32515 33457 32549 33483
rect 32515 33389 32549 33411
rect 32515 33321 32549 33339
rect 32515 33253 32549 33267
rect 32515 33185 32549 33195
rect 32515 33117 32549 33123
rect 32515 33049 32549 33051
rect 32515 33013 32549 33015
rect 32515 32941 32549 32947
rect 32515 32869 32549 32879
rect 32515 32797 32549 32811
rect 32515 32725 32549 32743
rect 32515 32653 32549 32675
rect 32515 32581 32549 32607
rect 32515 32509 32549 32539
rect 32515 32437 32549 32471
rect 32515 32302 32549 32403
rect 32973 33661 33007 33722
rect 32973 33593 33007 33627
rect 32973 33525 33007 33555
rect 32973 33457 33007 33483
rect 32973 33389 33007 33411
rect 32973 33321 33007 33339
rect 32973 33253 33007 33267
rect 32973 33185 33007 33195
rect 32973 33117 33007 33123
rect 32973 33049 33007 33051
rect 32973 33013 33007 33015
rect 32973 32941 33007 32947
rect 32973 32869 33007 32879
rect 32973 32797 33007 32811
rect 32973 32725 33007 32743
rect 32973 32653 33007 32675
rect 32973 32581 33007 32607
rect 32973 32509 33007 32539
rect 32973 32437 33007 32471
rect 32973 32383 33007 32403
rect 33431 33661 33465 33681
rect 33431 33593 33465 33627
rect 33431 33525 33465 33555
rect 33431 33457 33465 33483
rect 33431 33389 33465 33411
rect 33431 33321 33465 33339
rect 33431 33253 33465 33267
rect 33431 33185 33465 33195
rect 33431 33117 33465 33123
rect 33431 33049 33465 33051
rect 33431 33013 33465 33015
rect 33431 32941 33465 32947
rect 33431 32869 33465 32879
rect 33431 32797 33465 32811
rect 33431 32725 33465 32743
rect 33431 32653 33465 32675
rect 33431 32581 33465 32607
rect 33431 32509 33465 32539
rect 33431 32437 33465 32471
rect 33431 32302 33465 32403
rect 33889 33661 33923 33722
rect 33889 33593 33923 33627
rect 33889 33525 33923 33555
rect 33889 33457 33923 33483
rect 33889 33389 33923 33411
rect 33889 33321 33923 33339
rect 33889 33253 33923 33267
rect 33889 33185 33923 33195
rect 33889 33117 33923 33123
rect 33889 33049 33923 33051
rect 33889 33013 33923 33015
rect 33889 32941 33923 32947
rect 33889 32869 33923 32879
rect 33889 32797 33923 32811
rect 33889 32725 33923 32743
rect 33889 32653 33923 32675
rect 33889 32581 33923 32607
rect 33889 32509 33923 32539
rect 33889 32437 33923 32471
rect 33889 32383 33923 32403
rect 34347 33661 34381 33681
rect 34347 33593 34381 33627
rect 34347 33525 34381 33555
rect 34347 33457 34381 33483
rect 34347 33389 34381 33411
rect 34347 33321 34381 33339
rect 34347 33253 34381 33267
rect 34347 33185 34381 33195
rect 34347 33117 34381 33123
rect 34347 33049 34381 33051
rect 34347 33013 34381 33015
rect 34347 32941 34381 32947
rect 34347 32869 34381 32879
rect 34347 32797 34381 32811
rect 34347 32725 34381 32743
rect 34347 32653 34381 32675
rect 34347 32581 34381 32607
rect 34347 32509 34381 32539
rect 34347 32437 34381 32471
rect 34347 32302 34381 32403
rect 34805 33661 34839 33722
rect 34805 33593 34839 33627
rect 34805 33525 34839 33555
rect 34805 33457 34839 33483
rect 34805 33389 34839 33411
rect 34805 33321 34839 33339
rect 34805 33253 34839 33267
rect 34805 33185 34839 33195
rect 34805 33117 34839 33123
rect 34805 33049 34839 33051
rect 34805 33013 34839 33015
rect 34805 32941 34839 32947
rect 34805 32869 34839 32879
rect 34805 32797 34839 32811
rect 34805 32725 34839 32743
rect 34805 32653 34839 32675
rect 34805 32581 34839 32607
rect 34805 32509 34839 32539
rect 34805 32437 34839 32471
rect 34805 32383 34839 32403
rect 35263 33661 35297 33681
rect 35263 33593 35297 33627
rect 35263 33525 35297 33555
rect 35263 33457 35297 33483
rect 35263 33389 35297 33411
rect 35263 33321 35297 33339
rect 35263 33253 35297 33267
rect 35263 33185 35297 33195
rect 35263 33117 35297 33123
rect 35263 33049 35297 33051
rect 35263 33013 35297 33015
rect 35263 32941 35297 32947
rect 35263 32869 35297 32879
rect 35263 32797 35297 32811
rect 35263 32725 35297 32743
rect 35263 32653 35297 32675
rect 35263 32581 35297 32607
rect 35263 32509 35297 32539
rect 35263 32437 35297 32471
rect 35263 32302 35297 32403
rect 35721 33661 35755 33722
rect 35721 33593 35755 33627
rect 35721 33525 35755 33555
rect 35721 33457 35755 33483
rect 35721 33389 35755 33411
rect 35721 33321 35755 33339
rect 35721 33253 35755 33267
rect 35721 33185 35755 33195
rect 35721 33117 35755 33123
rect 35721 33049 35755 33051
rect 35721 33013 35755 33015
rect 35721 32941 35755 32947
rect 35721 32869 35755 32879
rect 35721 32797 35755 32811
rect 35721 32725 35755 32743
rect 35721 32653 35755 32675
rect 35721 32581 35755 32607
rect 35721 32509 35755 32539
rect 35721 32437 35755 32471
rect 35721 32383 35755 32403
rect 36179 33661 36213 33681
rect 36179 33593 36213 33627
rect 36179 33525 36213 33555
rect 36179 33457 36213 33483
rect 36179 33389 36213 33411
rect 36179 33321 36213 33339
rect 36179 33253 36213 33267
rect 36179 33185 36213 33195
rect 36179 33117 36213 33123
rect 36179 33049 36213 33051
rect 36179 33013 36213 33015
rect 36179 32941 36213 32947
rect 36179 32869 36213 32879
rect 36179 32797 36213 32811
rect 36179 32725 36213 32743
rect 36179 32653 36213 32675
rect 36179 32581 36213 32607
rect 36179 32509 36213 32539
rect 36179 32437 36213 32471
rect 36179 32302 36213 32403
rect 36637 33661 36671 33722
rect 36637 33593 36671 33627
rect 36637 33525 36671 33555
rect 36637 33457 36671 33483
rect 36637 33389 36671 33411
rect 36637 33321 36671 33339
rect 36637 33253 36671 33267
rect 36637 33185 36671 33195
rect 36637 33117 36671 33123
rect 36637 33049 36671 33051
rect 36637 33013 36671 33015
rect 36637 32941 36671 32947
rect 36637 32869 36671 32879
rect 36637 32797 36671 32811
rect 36637 32725 36671 32743
rect 36637 32653 36671 32675
rect 36637 32581 36671 32607
rect 36637 32509 36671 32539
rect 36637 32437 36671 32471
rect 36637 32383 36671 32403
rect 37095 33661 37129 33681
rect 37095 33593 37129 33627
rect 37095 33525 37129 33555
rect 37095 33457 37129 33483
rect 37095 33389 37129 33411
rect 37095 33321 37129 33339
rect 37095 33253 37129 33267
rect 37095 33185 37129 33195
rect 37095 33117 37129 33123
rect 37095 33049 37129 33051
rect 37095 33013 37129 33015
rect 37095 32941 37129 32947
rect 37095 32869 37129 32879
rect 37095 32797 37129 32811
rect 37095 32725 37129 32743
rect 37095 32653 37129 32675
rect 37095 32581 37129 32607
rect 37095 32509 37129 32539
rect 37095 32437 37129 32471
rect 37095 32302 37129 32403
rect 37553 33661 37587 33722
rect 37553 33593 37587 33627
rect 37553 33525 37587 33555
rect 37553 33457 37587 33483
rect 37553 33389 37587 33411
rect 37553 33321 37587 33339
rect 37553 33253 37587 33267
rect 37553 33185 37587 33195
rect 37553 33117 37587 33123
rect 37553 33049 37587 33051
rect 37553 33013 37587 33015
rect 37553 32941 37587 32947
rect 37553 32869 37587 32879
rect 37553 32797 37587 32811
rect 37553 32725 37587 32743
rect 37553 32653 37587 32675
rect 37553 32581 37587 32607
rect 37553 32509 37587 32539
rect 37553 32437 37587 32471
rect 37553 32383 37587 32403
rect 38011 33661 38045 33681
rect 38011 33593 38045 33627
rect 38011 33525 38045 33555
rect 38011 33457 38045 33483
rect 38011 33389 38045 33411
rect 38011 33321 38045 33339
rect 38011 33253 38045 33267
rect 38011 33185 38045 33195
rect 38011 33117 38045 33123
rect 38011 33049 38045 33051
rect 38011 33013 38045 33015
rect 38011 32941 38045 32947
rect 38011 32869 38045 32879
rect 38011 32797 38045 32811
rect 38011 32725 38045 32743
rect 38011 32653 38045 32675
rect 38011 32581 38045 32607
rect 38011 32509 38045 32539
rect 38011 32437 38045 32471
rect 38011 32302 38045 32403
rect 38469 33661 38503 33722
rect 38469 33593 38503 33627
rect 38469 33525 38503 33555
rect 38469 33457 38503 33483
rect 38469 33389 38503 33411
rect 38469 33321 38503 33339
rect 38469 33253 38503 33267
rect 38469 33185 38503 33195
rect 38469 33117 38503 33123
rect 38469 33049 38503 33051
rect 38469 33013 38503 33015
rect 38469 32941 38503 32947
rect 38469 32869 38503 32879
rect 38469 32797 38503 32811
rect 38469 32725 38503 32743
rect 38469 32653 38503 32675
rect 38469 32581 38503 32607
rect 38469 32509 38503 32539
rect 38469 32437 38503 32471
rect 38469 32383 38503 32403
rect 38927 33661 38961 33681
rect 38927 33593 38961 33627
rect 38927 33525 38961 33555
rect 38927 33457 38961 33483
rect 38927 33389 38961 33411
rect 38927 33321 38961 33339
rect 38927 33253 38961 33267
rect 38927 33185 38961 33195
rect 38927 33117 38961 33123
rect 38927 33049 38961 33051
rect 38927 33013 38961 33015
rect 38927 32941 38961 32947
rect 38927 32869 38961 32879
rect 38927 32797 38961 32811
rect 38927 32725 38961 32743
rect 38927 32653 38961 32675
rect 38927 32581 38961 32607
rect 38927 32509 38961 32539
rect 38927 32437 38961 32471
rect 38927 32302 38961 32403
rect 39385 33661 39419 33722
rect 39385 33593 39419 33627
rect 39385 33525 39419 33555
rect 39385 33457 39419 33483
rect 39385 33389 39419 33411
rect 39385 33321 39419 33339
rect 39385 33253 39419 33267
rect 39385 33185 39419 33195
rect 39385 33117 39419 33123
rect 39385 33049 39419 33051
rect 39385 33013 39419 33015
rect 39385 32941 39419 32947
rect 39385 32869 39419 32879
rect 39385 32797 39419 32811
rect 39385 32725 39419 32743
rect 39385 32653 39419 32675
rect 39385 32581 39419 32607
rect 39385 32509 39419 32539
rect 39385 32437 39419 32471
rect 39385 32383 39419 32403
rect 39843 33661 39877 33681
rect 39843 33593 39877 33627
rect 39843 33525 39877 33555
rect 39843 33457 39877 33483
rect 39843 33389 39877 33411
rect 39843 33321 39877 33339
rect 39843 33253 39877 33267
rect 39843 33185 39877 33195
rect 39843 33117 39877 33123
rect 39843 33049 39877 33051
rect 39843 33013 39877 33015
rect 39843 32941 39877 32947
rect 39843 32869 39877 32879
rect 39843 32797 39877 32811
rect 39843 32725 39877 32743
rect 39843 32653 39877 32675
rect 39843 32581 39877 32607
rect 39843 32509 39877 32539
rect 39843 32437 39877 32471
rect 39843 32302 39877 32403
rect 40301 33661 40335 33722
rect 40301 33593 40335 33627
rect 40301 33525 40335 33555
rect 40301 33457 40335 33483
rect 40301 33389 40335 33411
rect 40301 33321 40335 33339
rect 40301 33253 40335 33267
rect 40301 33185 40335 33195
rect 40301 33117 40335 33123
rect 40301 33049 40335 33051
rect 40301 33013 40335 33015
rect 40301 32941 40335 32947
rect 40301 32869 40335 32879
rect 40301 32797 40335 32811
rect 40301 32725 40335 32743
rect 40301 32653 40335 32675
rect 40301 32581 40335 32607
rect 40301 32509 40335 32539
rect 40301 32437 40335 32471
rect 40301 32383 40335 32403
rect 40759 33661 40793 33681
rect 40759 33593 40793 33627
rect 40759 33525 40793 33555
rect 40759 33457 40793 33483
rect 40759 33389 40793 33411
rect 40759 33321 40793 33339
rect 40759 33253 40793 33267
rect 40759 33185 40793 33195
rect 40759 33117 40793 33123
rect 40759 33049 40793 33051
rect 40759 33013 40793 33015
rect 40759 32941 40793 32947
rect 40759 32869 40793 32879
rect 40759 32797 40793 32811
rect 40759 32725 40793 32743
rect 40759 32653 40793 32675
rect 40759 32581 40793 32607
rect 40759 32509 40793 32539
rect 40759 32437 40793 32471
rect 40759 32302 40793 32403
rect 41217 33661 41251 33722
rect 41217 33593 41251 33627
rect 41217 33525 41251 33555
rect 41217 33457 41251 33483
rect 41217 33389 41251 33411
rect 41217 33321 41251 33339
rect 41217 33253 41251 33267
rect 41217 33185 41251 33195
rect 41217 33117 41251 33123
rect 41217 33049 41251 33051
rect 41217 33013 41251 33015
rect 41217 32941 41251 32947
rect 41217 32869 41251 32879
rect 41217 32797 41251 32811
rect 41217 32725 41251 32743
rect 41217 32653 41251 32675
rect 41217 32581 41251 32607
rect 41217 32509 41251 32539
rect 41217 32437 41251 32471
rect 41217 32383 41251 32403
rect 41675 33661 41709 33681
rect 41675 33593 41709 33627
rect 41675 33525 41709 33555
rect 41675 33457 41709 33483
rect 41675 33389 41709 33411
rect 41675 33321 41709 33339
rect 41675 33253 41709 33267
rect 41675 33185 41709 33195
rect 41675 33117 41709 33123
rect 41675 33049 41709 33051
rect 41675 33013 41709 33015
rect 41675 32941 41709 32947
rect 41675 32869 41709 32879
rect 41675 32797 41709 32811
rect 41675 32725 41709 32743
rect 41675 32653 41709 32675
rect 41675 32581 41709 32607
rect 41675 32509 41709 32539
rect 41675 32437 41709 32471
rect 41675 32302 41709 32403
rect 14148 32283 41756 32302
rect 14148 32249 26893 32283
rect 26927 32249 41756 32283
rect 14148 32242 41756 32249
rect 14148 32183 41756 32196
rect 14148 32181 14331 32183
rect 14148 32147 14197 32181
rect 14231 32149 14331 32181
rect 14365 32149 14731 32183
rect 14765 32149 15131 32183
rect 15165 32149 15531 32183
rect 15565 32149 15931 32183
rect 15965 32149 16331 32183
rect 16365 32149 16731 32183
rect 16765 32149 17131 32183
rect 17165 32149 17531 32183
rect 17565 32149 17931 32183
rect 17965 32149 18331 32183
rect 18365 32149 18731 32183
rect 18765 32149 19131 32183
rect 19165 32149 19531 32183
rect 19565 32149 19931 32183
rect 19965 32149 20331 32183
rect 20365 32149 20731 32183
rect 20765 32149 21131 32183
rect 21165 32149 21531 32183
rect 21565 32149 21931 32183
rect 21965 32149 22331 32183
rect 22365 32149 22731 32183
rect 22765 32149 23131 32183
rect 23165 32149 23531 32183
rect 23565 32149 23931 32183
rect 23965 32149 24331 32183
rect 24365 32149 24731 32183
rect 24765 32149 25131 32183
rect 25165 32149 25531 32183
rect 25565 32149 25931 32183
rect 25965 32149 26331 32183
rect 26365 32149 26731 32183
rect 26765 32149 27131 32183
rect 27165 32149 27531 32183
rect 27565 32149 27931 32183
rect 27965 32149 28331 32183
rect 28365 32149 28731 32183
rect 28765 32149 29131 32183
rect 29165 32149 29531 32183
rect 29565 32149 29931 32183
rect 29965 32149 30331 32183
rect 30365 32149 30731 32183
rect 30765 32149 31131 32183
rect 31165 32149 31531 32183
rect 31565 32149 31931 32183
rect 31965 32149 32331 32183
rect 32365 32149 32731 32183
rect 32765 32149 33131 32183
rect 33165 32149 33531 32183
rect 33565 32149 33931 32183
rect 33965 32149 34331 32183
rect 34365 32149 34731 32183
rect 34765 32149 35131 32183
rect 35165 32149 35531 32183
rect 35565 32149 35931 32183
rect 35965 32149 36331 32183
rect 36365 32149 36731 32183
rect 36765 32149 37131 32183
rect 37165 32149 37531 32183
rect 37565 32149 37931 32183
rect 37965 32149 38331 32183
rect 38365 32149 38731 32183
rect 38765 32149 39131 32183
rect 39165 32149 39531 32183
rect 39565 32149 39931 32183
rect 39965 32149 40331 32183
rect 40365 32149 40731 32183
rect 40765 32149 41131 32183
rect 41165 32149 41531 32183
rect 41565 32149 41756 32183
rect 14231 32147 41756 32149
rect 14148 32136 41756 32147
rect 6604 32049 13772 32062
rect 6604 32015 6787 32049
rect 6821 32015 7187 32049
rect 7221 32015 7587 32049
rect 7621 32015 7987 32049
rect 8021 32015 8387 32049
rect 8421 32015 8787 32049
rect 8821 32015 9187 32049
rect 9221 32015 9587 32049
rect 9621 32015 9987 32049
rect 10021 32015 10387 32049
rect 10421 32015 10787 32049
rect 10821 32015 11187 32049
rect 11221 32015 11587 32049
rect 11621 32015 11987 32049
rect 12021 32015 12387 32049
rect 12421 32015 12787 32049
rect 12821 32015 13187 32049
rect 13221 32015 13587 32049
rect 13621 32015 13772 32049
rect 6604 32002 13772 32015
rect 14050 32049 41756 32062
rect 14050 32015 14331 32049
rect 14365 32015 14731 32049
rect 14765 32015 15131 32049
rect 15165 32015 15531 32049
rect 15565 32015 15931 32049
rect 15965 32015 16331 32049
rect 16365 32015 16731 32049
rect 16765 32015 17131 32049
rect 17165 32015 17531 32049
rect 17565 32015 17931 32049
rect 17965 32015 18331 32049
rect 18365 32015 18731 32049
rect 18765 32015 19131 32049
rect 19165 32015 19531 32049
rect 19565 32015 19931 32049
rect 19965 32015 20331 32049
rect 20365 32015 20731 32049
rect 20765 32015 21131 32049
rect 21165 32015 21531 32049
rect 21565 32015 21931 32049
rect 21965 32015 22331 32049
rect 22365 32015 22731 32049
rect 22765 32015 23131 32049
rect 23165 32015 23531 32049
rect 23565 32015 23931 32049
rect 23965 32015 24331 32049
rect 24365 32015 24731 32049
rect 24765 32015 25131 32049
rect 25165 32015 25531 32049
rect 25565 32015 25931 32049
rect 25965 32015 26331 32049
rect 26365 32015 26731 32049
rect 26765 32015 27131 32049
rect 27165 32015 27531 32049
rect 27565 32015 27931 32049
rect 27965 32015 28331 32049
rect 28365 32015 28731 32049
rect 28765 32015 29131 32049
rect 29165 32015 29531 32049
rect 29565 32015 29931 32049
rect 29965 32015 30331 32049
rect 30365 32015 30731 32049
rect 30765 32015 31131 32049
rect 31165 32015 31531 32049
rect 31565 32015 31931 32049
rect 31965 32015 32331 32049
rect 32365 32015 32731 32049
rect 32765 32015 33131 32049
rect 33165 32015 33531 32049
rect 33565 32015 33931 32049
rect 33965 32015 34331 32049
rect 34365 32015 34731 32049
rect 34765 32015 35131 32049
rect 35165 32015 35531 32049
rect 35565 32015 35931 32049
rect 35965 32015 36331 32049
rect 36365 32015 36731 32049
rect 36765 32015 37131 32049
rect 37165 32015 37531 32049
rect 37565 32015 37931 32049
rect 37965 32015 38331 32049
rect 38365 32015 38731 32049
rect 38765 32015 39131 32049
rect 39165 32015 39531 32049
rect 39565 32015 39931 32049
rect 39965 32015 40331 32049
rect 40365 32015 40731 32049
rect 40765 32015 41131 32049
rect 41165 32015 41531 32049
rect 41565 32015 41756 32049
rect 14050 32002 41756 32015
rect 5916 30169 33622 30182
rect 5916 30135 6197 30169
rect 6231 30135 6597 30169
rect 6631 30135 6997 30169
rect 7031 30135 7397 30169
rect 7431 30135 7797 30169
rect 7831 30135 8197 30169
rect 8231 30135 8597 30169
rect 8631 30135 8997 30169
rect 9031 30135 9397 30169
rect 9431 30135 9797 30169
rect 9831 30135 10197 30169
rect 10231 30135 10597 30169
rect 10631 30135 10997 30169
rect 11031 30135 11397 30169
rect 11431 30135 11797 30169
rect 11831 30135 12197 30169
rect 12231 30135 12597 30169
rect 12631 30135 12997 30169
rect 13031 30135 13397 30169
rect 13431 30135 13797 30169
rect 13831 30135 14197 30169
rect 14231 30135 14597 30169
rect 14631 30135 14997 30169
rect 15031 30135 15397 30169
rect 15431 30135 15797 30169
rect 15831 30135 16197 30169
rect 16231 30135 16597 30169
rect 16631 30135 16997 30169
rect 17031 30135 17397 30169
rect 17431 30135 17797 30169
rect 17831 30135 18197 30169
rect 18231 30135 18597 30169
rect 18631 30135 18997 30169
rect 19031 30135 19397 30169
rect 19431 30135 19797 30169
rect 19831 30135 20197 30169
rect 20231 30135 20597 30169
rect 20631 30135 20997 30169
rect 21031 30135 21397 30169
rect 21431 30135 21797 30169
rect 21831 30135 22197 30169
rect 22231 30135 22597 30169
rect 22631 30135 22997 30169
rect 23031 30135 23397 30169
rect 23431 30135 23797 30169
rect 23831 30135 24197 30169
rect 24231 30135 24597 30169
rect 24631 30135 24997 30169
rect 25031 30135 25397 30169
rect 25431 30135 25797 30169
rect 25831 30135 26197 30169
rect 26231 30135 26597 30169
rect 26631 30135 26997 30169
rect 27031 30135 27397 30169
rect 27431 30135 27797 30169
rect 27831 30135 28197 30169
rect 28231 30135 28597 30169
rect 28631 30135 28997 30169
rect 29031 30135 29397 30169
rect 29431 30135 29797 30169
rect 29831 30135 30197 30169
rect 30231 30135 30597 30169
rect 30631 30135 30997 30169
rect 31031 30135 31397 30169
rect 31431 30135 31797 30169
rect 31831 30135 32197 30169
rect 32231 30135 32597 30169
rect 32631 30135 32997 30169
rect 33031 30135 33397 30169
rect 33431 30135 33622 30169
rect 5916 30122 33622 30135
rect 33944 30169 36918 30182
rect 33944 30135 34225 30169
rect 34259 30135 34625 30169
rect 34659 30135 35025 30169
rect 35059 30135 35425 30169
rect 35459 30135 35825 30169
rect 35859 30135 36225 30169
rect 36259 30135 36625 30169
rect 36659 30135 36918 30169
rect 33944 30122 36918 30135
rect 37394 30169 39834 30182
rect 37394 30135 37577 30169
rect 37611 30135 37777 30169
rect 37811 30135 37977 30169
rect 38011 30135 38177 30169
rect 38211 30135 38377 30169
rect 38411 30135 38577 30169
rect 38611 30135 38777 30169
rect 38811 30135 38977 30169
rect 39011 30135 39177 30169
rect 39211 30135 39377 30169
rect 39411 30135 39577 30169
rect 39611 30135 39834 30169
rect 37394 30122 39834 30135
rect 40138 30169 42578 30182
rect 40138 30135 40321 30169
rect 40355 30135 40521 30169
rect 40555 30135 40721 30169
rect 40755 30135 40921 30169
rect 40955 30135 41121 30169
rect 41155 30135 41321 30169
rect 41355 30135 41521 30169
rect 41555 30135 41721 30169
rect 41755 30135 41921 30169
rect 41955 30135 42121 30169
rect 42155 30135 42321 30169
rect 42355 30135 42578 30169
rect 40138 30122 42578 30135
rect 5944 30029 6004 30122
rect 6992 30079 7152 30122
rect 6992 30045 7057 30079
rect 7091 30045 7152 30079
rect 6992 30042 7152 30045
rect 8292 30079 8452 30122
rect 8292 30045 8357 30079
rect 8391 30045 8452 30079
rect 8292 30042 8452 30045
rect 9592 30079 9752 30122
rect 9592 30045 9657 30079
rect 9691 30045 9752 30079
rect 9592 30042 9752 30045
rect 10892 30079 11052 30122
rect 10892 30045 10957 30079
rect 10991 30045 11052 30079
rect 10892 30042 11052 30045
rect 12192 30079 12352 30122
rect 12192 30045 12257 30079
rect 12291 30045 12352 30079
rect 12192 30042 12352 30045
rect 13492 30079 13652 30122
rect 13492 30045 13557 30079
rect 13591 30045 13652 30079
rect 13492 30042 13652 30045
rect 14792 30079 14952 30122
rect 14792 30045 14857 30079
rect 14891 30045 14952 30079
rect 14792 30042 14952 30045
rect 16092 30079 16252 30122
rect 16092 30045 16157 30079
rect 16191 30045 16252 30079
rect 16092 30042 16252 30045
rect 17392 30079 17552 30122
rect 17392 30045 17457 30079
rect 17491 30045 17552 30079
rect 17392 30042 17552 30045
rect 18692 30079 18852 30122
rect 18692 30045 18757 30079
rect 18791 30045 18852 30079
rect 18692 30042 18852 30045
rect 19992 30079 20152 30122
rect 19992 30045 20057 30079
rect 20091 30045 20152 30079
rect 19992 30042 20152 30045
rect 21292 30079 21452 30122
rect 21292 30045 21357 30079
rect 21391 30045 21452 30079
rect 21292 30042 21452 30045
rect 22592 30079 22752 30122
rect 22592 30045 22657 30079
rect 22691 30045 22752 30079
rect 22592 30042 22752 30045
rect 23892 30079 24052 30122
rect 23892 30045 23957 30079
rect 23991 30045 24052 30079
rect 23892 30042 24052 30045
rect 25192 30079 25352 30122
rect 25192 30045 25257 30079
rect 25291 30045 25352 30079
rect 25192 30042 25352 30045
rect 26492 30079 26652 30122
rect 26492 30045 26557 30079
rect 26591 30045 26652 30079
rect 26492 30042 26652 30045
rect 27792 30079 27952 30122
rect 27792 30045 27857 30079
rect 27891 30045 27952 30079
rect 27792 30042 27952 30045
rect 29092 30079 29252 30122
rect 29092 30045 29157 30079
rect 29191 30045 29252 30079
rect 29092 30042 29252 30045
rect 30392 30079 30552 30122
rect 30392 30045 30457 30079
rect 30491 30045 30552 30079
rect 30392 30042 30552 30045
rect 31692 30079 31852 30122
rect 31692 30045 31757 30079
rect 31791 30045 31852 30079
rect 31692 30042 31852 30045
rect 5944 29995 5957 30029
rect 5991 29995 6004 30029
rect 33972 30029 34032 30122
rect 35020 30079 35180 30122
rect 35020 30045 35085 30079
rect 35119 30045 35180 30079
rect 35020 30042 35180 30045
rect 5944 29912 6004 29995
rect 6074 29962 33622 30002
rect 33972 29995 33985 30029
rect 34019 29995 34032 30029
rect 6061 29901 6095 29921
rect 6061 29833 6095 29867
rect 6061 29765 6095 29795
rect 6061 29697 6095 29723
rect 6061 29629 6095 29651
rect 6061 29561 6095 29579
rect 6061 29493 6095 29507
rect 6061 29425 6095 29435
rect 6061 29357 6095 29363
rect 6061 29289 6095 29291
rect 6061 29253 6095 29255
rect 6061 29181 6095 29187
rect 6061 29109 6095 29119
rect 6061 29037 6095 29051
rect 6061 28965 6095 28983
rect 6061 28893 6095 28915
rect 6061 28821 6095 28847
rect 6061 28749 6095 28779
rect 6061 28677 6095 28711
rect 6061 28542 6095 28643
rect 6519 29901 6553 29962
rect 6519 29833 6553 29867
rect 6519 29765 6553 29795
rect 6519 29697 6553 29723
rect 6519 29629 6553 29651
rect 6519 29561 6553 29579
rect 6519 29493 6553 29507
rect 6519 29425 6553 29435
rect 6519 29357 6553 29363
rect 6519 29289 6553 29291
rect 6519 29253 6553 29255
rect 6519 29181 6553 29187
rect 6519 29109 6553 29119
rect 6519 29037 6553 29051
rect 6519 28965 6553 28983
rect 6519 28893 6553 28915
rect 6519 28821 6553 28847
rect 6519 28749 6553 28779
rect 6519 28677 6553 28711
rect 6519 28623 6553 28643
rect 6977 29901 7011 29921
rect 6977 29833 7011 29867
rect 6977 29765 7011 29795
rect 6977 29697 7011 29723
rect 6977 29629 7011 29651
rect 6977 29561 7011 29579
rect 6977 29493 7011 29507
rect 6977 29425 7011 29435
rect 6977 29357 7011 29363
rect 6977 29289 7011 29291
rect 6977 29253 7011 29255
rect 6977 29181 7011 29187
rect 6977 29109 7011 29119
rect 6977 29037 7011 29051
rect 6977 28965 7011 28983
rect 6977 28893 7011 28915
rect 6977 28821 7011 28847
rect 6977 28749 7011 28779
rect 6977 28677 7011 28711
rect 6977 28542 7011 28643
rect 7435 29901 7469 29962
rect 7435 29833 7469 29867
rect 7435 29765 7469 29795
rect 7435 29697 7469 29723
rect 7435 29629 7469 29651
rect 7435 29561 7469 29579
rect 7435 29493 7469 29507
rect 7435 29425 7469 29435
rect 7435 29357 7469 29363
rect 7435 29289 7469 29291
rect 7435 29253 7469 29255
rect 7435 29181 7469 29187
rect 7435 29109 7469 29119
rect 7435 29037 7469 29051
rect 7435 28965 7469 28983
rect 7435 28893 7469 28915
rect 7435 28821 7469 28847
rect 7435 28749 7469 28779
rect 7435 28677 7469 28711
rect 7435 28623 7469 28643
rect 7893 29901 7927 29921
rect 7893 29833 7927 29867
rect 7893 29765 7927 29795
rect 7893 29697 7927 29723
rect 7893 29629 7927 29651
rect 7893 29561 7927 29579
rect 7893 29493 7927 29507
rect 7893 29425 7927 29435
rect 7893 29357 7927 29363
rect 7893 29289 7927 29291
rect 7893 29253 7927 29255
rect 7893 29181 7927 29187
rect 7893 29109 7927 29119
rect 7893 29037 7927 29051
rect 7893 28965 7927 28983
rect 7893 28893 7927 28915
rect 7893 28821 7927 28847
rect 7893 28749 7927 28779
rect 7893 28677 7927 28711
rect 7893 28542 7927 28643
rect 8351 29901 8385 29962
rect 8351 29833 8385 29867
rect 8351 29765 8385 29795
rect 8351 29697 8385 29723
rect 8351 29629 8385 29651
rect 8351 29561 8385 29579
rect 8351 29493 8385 29507
rect 8351 29425 8385 29435
rect 8351 29357 8385 29363
rect 8351 29289 8385 29291
rect 8351 29253 8385 29255
rect 8351 29181 8385 29187
rect 8351 29109 8385 29119
rect 8351 29037 8385 29051
rect 8351 28965 8385 28983
rect 8351 28893 8385 28915
rect 8351 28821 8385 28847
rect 8351 28749 8385 28779
rect 8351 28677 8385 28711
rect 8351 28623 8385 28643
rect 8809 29901 8843 29921
rect 8809 29833 8843 29867
rect 8809 29765 8843 29795
rect 8809 29697 8843 29723
rect 8809 29629 8843 29651
rect 8809 29561 8843 29579
rect 8809 29493 8843 29507
rect 8809 29425 8843 29435
rect 8809 29357 8843 29363
rect 8809 29289 8843 29291
rect 8809 29253 8843 29255
rect 8809 29181 8843 29187
rect 8809 29109 8843 29119
rect 8809 29037 8843 29051
rect 8809 28965 8843 28983
rect 8809 28893 8843 28915
rect 8809 28821 8843 28847
rect 8809 28749 8843 28779
rect 8809 28677 8843 28711
rect 8809 28542 8843 28643
rect 9267 29901 9301 29962
rect 9267 29833 9301 29867
rect 9267 29765 9301 29795
rect 9267 29697 9301 29723
rect 9267 29629 9301 29651
rect 9267 29561 9301 29579
rect 9267 29493 9301 29507
rect 9267 29425 9301 29435
rect 9267 29357 9301 29363
rect 9267 29289 9301 29291
rect 9267 29253 9301 29255
rect 9267 29181 9301 29187
rect 9267 29109 9301 29119
rect 9267 29037 9301 29051
rect 9267 28965 9301 28983
rect 9267 28893 9301 28915
rect 9267 28821 9301 28847
rect 9267 28749 9301 28779
rect 9267 28677 9301 28711
rect 9267 28623 9301 28643
rect 9725 29901 9759 29921
rect 9725 29833 9759 29867
rect 9725 29765 9759 29795
rect 9725 29697 9759 29723
rect 9725 29629 9759 29651
rect 9725 29561 9759 29579
rect 9725 29493 9759 29507
rect 9725 29425 9759 29435
rect 9725 29357 9759 29363
rect 9725 29289 9759 29291
rect 9725 29253 9759 29255
rect 9725 29181 9759 29187
rect 9725 29109 9759 29119
rect 9725 29037 9759 29051
rect 9725 28965 9759 28983
rect 9725 28893 9759 28915
rect 9725 28821 9759 28847
rect 9725 28749 9759 28779
rect 9725 28677 9759 28711
rect 9725 28542 9759 28643
rect 10183 29901 10217 29962
rect 10183 29833 10217 29867
rect 10183 29765 10217 29795
rect 10183 29697 10217 29723
rect 10183 29629 10217 29651
rect 10183 29561 10217 29579
rect 10183 29493 10217 29507
rect 10183 29425 10217 29435
rect 10183 29357 10217 29363
rect 10183 29289 10217 29291
rect 10183 29253 10217 29255
rect 10183 29181 10217 29187
rect 10183 29109 10217 29119
rect 10183 29037 10217 29051
rect 10183 28965 10217 28983
rect 10183 28893 10217 28915
rect 10183 28821 10217 28847
rect 10183 28749 10217 28779
rect 10183 28677 10217 28711
rect 10183 28623 10217 28643
rect 10641 29901 10675 29921
rect 10641 29833 10675 29867
rect 10641 29765 10675 29795
rect 10641 29697 10675 29723
rect 10641 29629 10675 29651
rect 10641 29561 10675 29579
rect 10641 29493 10675 29507
rect 10641 29425 10675 29435
rect 10641 29357 10675 29363
rect 10641 29289 10675 29291
rect 10641 29253 10675 29255
rect 10641 29181 10675 29187
rect 10641 29109 10675 29119
rect 10641 29037 10675 29051
rect 10641 28965 10675 28983
rect 10641 28893 10675 28915
rect 10641 28821 10675 28847
rect 10641 28749 10675 28779
rect 10641 28677 10675 28711
rect 10641 28542 10675 28643
rect 11099 29901 11133 29962
rect 11099 29833 11133 29867
rect 11099 29765 11133 29795
rect 11099 29697 11133 29723
rect 11099 29629 11133 29651
rect 11099 29561 11133 29579
rect 11099 29493 11133 29507
rect 11099 29425 11133 29435
rect 11099 29357 11133 29363
rect 11099 29289 11133 29291
rect 11099 29253 11133 29255
rect 11099 29181 11133 29187
rect 11099 29109 11133 29119
rect 11099 29037 11133 29051
rect 11099 28965 11133 28983
rect 11099 28893 11133 28915
rect 11099 28821 11133 28847
rect 11099 28749 11133 28779
rect 11099 28677 11133 28711
rect 11099 28623 11133 28643
rect 11557 29901 11591 29921
rect 11557 29833 11591 29867
rect 11557 29765 11591 29795
rect 11557 29697 11591 29723
rect 11557 29629 11591 29651
rect 11557 29561 11591 29579
rect 11557 29493 11591 29507
rect 11557 29425 11591 29435
rect 11557 29357 11591 29363
rect 11557 29289 11591 29291
rect 11557 29253 11591 29255
rect 11557 29181 11591 29187
rect 11557 29109 11591 29119
rect 11557 29037 11591 29051
rect 11557 28965 11591 28983
rect 11557 28893 11591 28915
rect 11557 28821 11591 28847
rect 11557 28749 11591 28779
rect 11557 28677 11591 28711
rect 11557 28542 11591 28643
rect 12015 29901 12049 29962
rect 12015 29833 12049 29867
rect 12015 29765 12049 29795
rect 12015 29697 12049 29723
rect 12015 29629 12049 29651
rect 12015 29561 12049 29579
rect 12015 29493 12049 29507
rect 12015 29425 12049 29435
rect 12015 29357 12049 29363
rect 12015 29289 12049 29291
rect 12015 29253 12049 29255
rect 12015 29181 12049 29187
rect 12015 29109 12049 29119
rect 12015 29037 12049 29051
rect 12015 28965 12049 28983
rect 12015 28893 12049 28915
rect 12015 28821 12049 28847
rect 12015 28749 12049 28779
rect 12015 28677 12049 28711
rect 12015 28623 12049 28643
rect 12473 29901 12507 29921
rect 12473 29833 12507 29867
rect 12473 29765 12507 29795
rect 12473 29697 12507 29723
rect 12473 29629 12507 29651
rect 12473 29561 12507 29579
rect 12473 29493 12507 29507
rect 12473 29425 12507 29435
rect 12473 29357 12507 29363
rect 12473 29289 12507 29291
rect 12473 29253 12507 29255
rect 12473 29181 12507 29187
rect 12473 29109 12507 29119
rect 12473 29037 12507 29051
rect 12473 28965 12507 28983
rect 12473 28893 12507 28915
rect 12473 28821 12507 28847
rect 12473 28749 12507 28779
rect 12473 28677 12507 28711
rect 12473 28542 12507 28643
rect 12931 29901 12965 29962
rect 12931 29833 12965 29867
rect 12931 29765 12965 29795
rect 12931 29697 12965 29723
rect 12931 29629 12965 29651
rect 12931 29561 12965 29579
rect 12931 29493 12965 29507
rect 12931 29425 12965 29435
rect 12931 29357 12965 29363
rect 12931 29289 12965 29291
rect 12931 29253 12965 29255
rect 12931 29181 12965 29187
rect 12931 29109 12965 29119
rect 12931 29037 12965 29051
rect 12931 28965 12965 28983
rect 12931 28893 12965 28915
rect 12931 28821 12965 28847
rect 12931 28749 12965 28779
rect 12931 28677 12965 28711
rect 12931 28623 12965 28643
rect 13389 29901 13423 29921
rect 13389 29833 13423 29867
rect 13389 29765 13423 29795
rect 13389 29697 13423 29723
rect 13389 29629 13423 29651
rect 13389 29561 13423 29579
rect 13389 29493 13423 29507
rect 13389 29425 13423 29435
rect 13389 29357 13423 29363
rect 13389 29289 13423 29291
rect 13389 29253 13423 29255
rect 13389 29181 13423 29187
rect 13389 29109 13423 29119
rect 13389 29037 13423 29051
rect 13389 28965 13423 28983
rect 13389 28893 13423 28915
rect 13389 28821 13423 28847
rect 13389 28749 13423 28779
rect 13389 28677 13423 28711
rect 13389 28542 13423 28643
rect 13847 29901 13881 29962
rect 13847 29833 13881 29867
rect 13847 29765 13881 29795
rect 13847 29697 13881 29723
rect 13847 29629 13881 29651
rect 13847 29561 13881 29579
rect 13847 29493 13881 29507
rect 13847 29425 13881 29435
rect 13847 29357 13881 29363
rect 13847 29289 13881 29291
rect 13847 29253 13881 29255
rect 13847 29181 13881 29187
rect 13847 29109 13881 29119
rect 13847 29037 13881 29051
rect 13847 28965 13881 28983
rect 13847 28893 13881 28915
rect 13847 28821 13881 28847
rect 13847 28749 13881 28779
rect 13847 28677 13881 28711
rect 13847 28623 13881 28643
rect 14305 29901 14339 29921
rect 14305 29833 14339 29867
rect 14305 29765 14339 29795
rect 14305 29697 14339 29723
rect 14305 29629 14339 29651
rect 14305 29561 14339 29579
rect 14305 29493 14339 29507
rect 14305 29425 14339 29435
rect 14305 29357 14339 29363
rect 14305 29289 14339 29291
rect 14305 29253 14339 29255
rect 14305 29181 14339 29187
rect 14305 29109 14339 29119
rect 14305 29037 14339 29051
rect 14305 28965 14339 28983
rect 14305 28893 14339 28915
rect 14305 28821 14339 28847
rect 14305 28749 14339 28779
rect 14305 28677 14339 28711
rect 14305 28542 14339 28643
rect 14763 29901 14797 29962
rect 14763 29833 14797 29867
rect 14763 29765 14797 29795
rect 14763 29697 14797 29723
rect 14763 29629 14797 29651
rect 14763 29561 14797 29579
rect 14763 29493 14797 29507
rect 14763 29425 14797 29435
rect 14763 29357 14797 29363
rect 14763 29289 14797 29291
rect 14763 29253 14797 29255
rect 14763 29181 14797 29187
rect 14763 29109 14797 29119
rect 14763 29037 14797 29051
rect 14763 28965 14797 28983
rect 14763 28893 14797 28915
rect 14763 28821 14797 28847
rect 14763 28749 14797 28779
rect 14763 28677 14797 28711
rect 14763 28623 14797 28643
rect 15221 29901 15255 29921
rect 15221 29833 15255 29867
rect 15221 29765 15255 29795
rect 15221 29697 15255 29723
rect 15221 29629 15255 29651
rect 15221 29561 15255 29579
rect 15221 29493 15255 29507
rect 15221 29425 15255 29435
rect 15221 29357 15255 29363
rect 15221 29289 15255 29291
rect 15221 29253 15255 29255
rect 15221 29181 15255 29187
rect 15221 29109 15255 29119
rect 15221 29037 15255 29051
rect 15221 28965 15255 28983
rect 15221 28893 15255 28915
rect 15221 28821 15255 28847
rect 15221 28749 15255 28779
rect 15221 28677 15255 28711
rect 15221 28542 15255 28643
rect 15679 29901 15713 29962
rect 15679 29833 15713 29867
rect 15679 29765 15713 29795
rect 15679 29697 15713 29723
rect 15679 29629 15713 29651
rect 15679 29561 15713 29579
rect 15679 29493 15713 29507
rect 15679 29425 15713 29435
rect 15679 29357 15713 29363
rect 15679 29289 15713 29291
rect 15679 29253 15713 29255
rect 15679 29181 15713 29187
rect 15679 29109 15713 29119
rect 15679 29037 15713 29051
rect 15679 28965 15713 28983
rect 15679 28893 15713 28915
rect 15679 28821 15713 28847
rect 15679 28749 15713 28779
rect 15679 28677 15713 28711
rect 15679 28623 15713 28643
rect 16137 29901 16171 29921
rect 16137 29833 16171 29867
rect 16137 29765 16171 29795
rect 16137 29697 16171 29723
rect 16137 29629 16171 29651
rect 16137 29561 16171 29579
rect 16137 29493 16171 29507
rect 16137 29425 16171 29435
rect 16137 29357 16171 29363
rect 16137 29289 16171 29291
rect 16137 29253 16171 29255
rect 16137 29181 16171 29187
rect 16137 29109 16171 29119
rect 16137 29037 16171 29051
rect 16137 28965 16171 28983
rect 16137 28893 16171 28915
rect 16137 28821 16171 28847
rect 16137 28749 16171 28779
rect 16137 28677 16171 28711
rect 16137 28542 16171 28643
rect 16595 29901 16629 29962
rect 16595 29833 16629 29867
rect 16595 29765 16629 29795
rect 16595 29697 16629 29723
rect 16595 29629 16629 29651
rect 16595 29561 16629 29579
rect 16595 29493 16629 29507
rect 16595 29425 16629 29435
rect 16595 29357 16629 29363
rect 16595 29289 16629 29291
rect 16595 29253 16629 29255
rect 16595 29181 16629 29187
rect 16595 29109 16629 29119
rect 16595 29037 16629 29051
rect 16595 28965 16629 28983
rect 16595 28893 16629 28915
rect 16595 28821 16629 28847
rect 16595 28749 16629 28779
rect 16595 28677 16629 28711
rect 16595 28623 16629 28643
rect 17053 29901 17087 29921
rect 17053 29833 17087 29867
rect 17053 29765 17087 29795
rect 17053 29697 17087 29723
rect 17053 29629 17087 29651
rect 17053 29561 17087 29579
rect 17053 29493 17087 29507
rect 17053 29425 17087 29435
rect 17053 29357 17087 29363
rect 17053 29289 17087 29291
rect 17053 29253 17087 29255
rect 17053 29181 17087 29187
rect 17053 29109 17087 29119
rect 17053 29037 17087 29051
rect 17053 28965 17087 28983
rect 17053 28893 17087 28915
rect 17053 28821 17087 28847
rect 17053 28749 17087 28779
rect 17053 28677 17087 28711
rect 17053 28542 17087 28643
rect 17511 29901 17545 29962
rect 17511 29833 17545 29867
rect 17511 29765 17545 29795
rect 17511 29697 17545 29723
rect 17511 29629 17545 29651
rect 17511 29561 17545 29579
rect 17511 29493 17545 29507
rect 17511 29425 17545 29435
rect 17511 29357 17545 29363
rect 17511 29289 17545 29291
rect 17511 29253 17545 29255
rect 17511 29181 17545 29187
rect 17511 29109 17545 29119
rect 17511 29037 17545 29051
rect 17511 28965 17545 28983
rect 17511 28893 17545 28915
rect 17511 28821 17545 28847
rect 17511 28749 17545 28779
rect 17511 28677 17545 28711
rect 17511 28623 17545 28643
rect 17969 29901 18003 29921
rect 17969 29833 18003 29867
rect 17969 29765 18003 29795
rect 17969 29697 18003 29723
rect 17969 29629 18003 29651
rect 17969 29561 18003 29579
rect 17969 29493 18003 29507
rect 17969 29425 18003 29435
rect 17969 29357 18003 29363
rect 17969 29289 18003 29291
rect 17969 29253 18003 29255
rect 17969 29181 18003 29187
rect 17969 29109 18003 29119
rect 17969 29037 18003 29051
rect 17969 28965 18003 28983
rect 17969 28893 18003 28915
rect 17969 28821 18003 28847
rect 17969 28749 18003 28779
rect 17969 28677 18003 28711
rect 17969 28542 18003 28643
rect 18427 29901 18461 29962
rect 18427 29833 18461 29867
rect 18427 29765 18461 29795
rect 18427 29697 18461 29723
rect 18427 29629 18461 29651
rect 18427 29561 18461 29579
rect 18427 29493 18461 29507
rect 18427 29425 18461 29435
rect 18427 29357 18461 29363
rect 18427 29289 18461 29291
rect 18427 29253 18461 29255
rect 18427 29181 18461 29187
rect 18427 29109 18461 29119
rect 18427 29037 18461 29051
rect 18427 28965 18461 28983
rect 18427 28893 18461 28915
rect 18427 28821 18461 28847
rect 18427 28749 18461 28779
rect 18427 28677 18461 28711
rect 18427 28623 18461 28643
rect 18885 29901 18919 29921
rect 18885 29833 18919 29867
rect 18885 29765 18919 29795
rect 18885 29697 18919 29723
rect 18885 29629 18919 29651
rect 18885 29561 18919 29579
rect 18885 29493 18919 29507
rect 18885 29425 18919 29435
rect 18885 29357 18919 29363
rect 18885 29289 18919 29291
rect 18885 29253 18919 29255
rect 18885 29181 18919 29187
rect 18885 29109 18919 29119
rect 18885 29037 18919 29051
rect 18885 28965 18919 28983
rect 18885 28893 18919 28915
rect 18885 28821 18919 28847
rect 18885 28749 18919 28779
rect 18885 28677 18919 28711
rect 18885 28542 18919 28643
rect 19343 29901 19377 29962
rect 19343 29833 19377 29867
rect 19343 29765 19377 29795
rect 19343 29697 19377 29723
rect 19343 29629 19377 29651
rect 19343 29561 19377 29579
rect 19343 29493 19377 29507
rect 19343 29425 19377 29435
rect 19343 29357 19377 29363
rect 19343 29289 19377 29291
rect 19343 29253 19377 29255
rect 19343 29181 19377 29187
rect 19343 29109 19377 29119
rect 19343 29037 19377 29051
rect 19343 28965 19377 28983
rect 19343 28893 19377 28915
rect 19343 28821 19377 28847
rect 19343 28749 19377 28779
rect 19343 28677 19377 28711
rect 19343 28623 19377 28643
rect 19801 29901 19835 29921
rect 19801 29833 19835 29867
rect 19801 29765 19835 29795
rect 19801 29697 19835 29723
rect 19801 29629 19835 29651
rect 19801 29561 19835 29579
rect 19801 29493 19835 29507
rect 19801 29425 19835 29435
rect 19801 29357 19835 29363
rect 19801 29289 19835 29291
rect 19801 29253 19835 29255
rect 19801 29181 19835 29187
rect 19801 29109 19835 29119
rect 19801 29037 19835 29051
rect 19801 28965 19835 28983
rect 19801 28893 19835 28915
rect 19801 28821 19835 28847
rect 19801 28749 19835 28779
rect 19801 28677 19835 28711
rect 19801 28542 19835 28643
rect 20259 29901 20293 29962
rect 20259 29833 20293 29867
rect 20259 29765 20293 29795
rect 20259 29697 20293 29723
rect 20259 29629 20293 29651
rect 20259 29561 20293 29579
rect 20259 29493 20293 29507
rect 20259 29425 20293 29435
rect 20259 29357 20293 29363
rect 20259 29289 20293 29291
rect 20259 29253 20293 29255
rect 20259 29181 20293 29187
rect 20259 29109 20293 29119
rect 20259 29037 20293 29051
rect 20259 28965 20293 28983
rect 20259 28893 20293 28915
rect 20259 28821 20293 28847
rect 20259 28749 20293 28779
rect 20259 28677 20293 28711
rect 20259 28623 20293 28643
rect 20717 29901 20751 29921
rect 20717 29833 20751 29867
rect 20717 29765 20751 29795
rect 20717 29697 20751 29723
rect 20717 29629 20751 29651
rect 20717 29561 20751 29579
rect 20717 29493 20751 29507
rect 20717 29425 20751 29435
rect 20717 29357 20751 29363
rect 20717 29289 20751 29291
rect 20717 29253 20751 29255
rect 20717 29181 20751 29187
rect 20717 29109 20751 29119
rect 20717 29037 20751 29051
rect 20717 28965 20751 28983
rect 20717 28893 20751 28915
rect 20717 28821 20751 28847
rect 20717 28749 20751 28779
rect 20717 28677 20751 28711
rect 20717 28542 20751 28643
rect 21175 29901 21209 29962
rect 21175 29833 21209 29867
rect 21175 29765 21209 29795
rect 21175 29697 21209 29723
rect 21175 29629 21209 29651
rect 21175 29561 21209 29579
rect 21175 29493 21209 29507
rect 21175 29425 21209 29435
rect 21175 29357 21209 29363
rect 21175 29289 21209 29291
rect 21175 29253 21209 29255
rect 21175 29181 21209 29187
rect 21175 29109 21209 29119
rect 21175 29037 21209 29051
rect 21175 28965 21209 28983
rect 21175 28893 21209 28915
rect 21175 28821 21209 28847
rect 21175 28749 21209 28779
rect 21175 28677 21209 28711
rect 21175 28623 21209 28643
rect 21633 29901 21667 29921
rect 21633 29833 21667 29867
rect 21633 29765 21667 29795
rect 21633 29697 21667 29723
rect 21633 29629 21667 29651
rect 21633 29561 21667 29579
rect 21633 29493 21667 29507
rect 21633 29425 21667 29435
rect 21633 29357 21667 29363
rect 21633 29289 21667 29291
rect 21633 29253 21667 29255
rect 21633 29181 21667 29187
rect 21633 29109 21667 29119
rect 21633 29037 21667 29051
rect 21633 28965 21667 28983
rect 21633 28893 21667 28915
rect 21633 28821 21667 28847
rect 21633 28749 21667 28779
rect 21633 28677 21667 28711
rect 21633 28542 21667 28643
rect 22091 29901 22125 29962
rect 22091 29833 22125 29867
rect 22091 29765 22125 29795
rect 22091 29697 22125 29723
rect 22091 29629 22125 29651
rect 22091 29561 22125 29579
rect 22091 29493 22125 29507
rect 22091 29425 22125 29435
rect 22091 29357 22125 29363
rect 22091 29289 22125 29291
rect 22091 29253 22125 29255
rect 22091 29181 22125 29187
rect 22091 29109 22125 29119
rect 22091 29037 22125 29051
rect 22091 28965 22125 28983
rect 22091 28893 22125 28915
rect 22091 28821 22125 28847
rect 22091 28749 22125 28779
rect 22091 28677 22125 28711
rect 22091 28623 22125 28643
rect 22549 29901 22583 29921
rect 22549 29833 22583 29867
rect 22549 29765 22583 29795
rect 22549 29697 22583 29723
rect 22549 29629 22583 29651
rect 22549 29561 22583 29579
rect 22549 29493 22583 29507
rect 22549 29425 22583 29435
rect 22549 29357 22583 29363
rect 22549 29289 22583 29291
rect 22549 29253 22583 29255
rect 22549 29181 22583 29187
rect 22549 29109 22583 29119
rect 22549 29037 22583 29051
rect 22549 28965 22583 28983
rect 22549 28893 22583 28915
rect 22549 28821 22583 28847
rect 22549 28749 22583 28779
rect 22549 28677 22583 28711
rect 22549 28542 22583 28643
rect 23007 29901 23041 29962
rect 23007 29833 23041 29867
rect 23007 29765 23041 29795
rect 23007 29697 23041 29723
rect 23007 29629 23041 29651
rect 23007 29561 23041 29579
rect 23007 29493 23041 29507
rect 23007 29425 23041 29435
rect 23007 29357 23041 29363
rect 23007 29289 23041 29291
rect 23007 29253 23041 29255
rect 23007 29181 23041 29187
rect 23007 29109 23041 29119
rect 23007 29037 23041 29051
rect 23007 28965 23041 28983
rect 23007 28893 23041 28915
rect 23007 28821 23041 28847
rect 23007 28749 23041 28779
rect 23007 28677 23041 28711
rect 23007 28623 23041 28643
rect 23465 29901 23499 29921
rect 23465 29833 23499 29867
rect 23465 29765 23499 29795
rect 23465 29697 23499 29723
rect 23465 29629 23499 29651
rect 23465 29561 23499 29579
rect 23465 29493 23499 29507
rect 23465 29425 23499 29435
rect 23465 29357 23499 29363
rect 23465 29289 23499 29291
rect 23465 29253 23499 29255
rect 23465 29181 23499 29187
rect 23465 29109 23499 29119
rect 23465 29037 23499 29051
rect 23465 28965 23499 28983
rect 23465 28893 23499 28915
rect 23465 28821 23499 28847
rect 23465 28749 23499 28779
rect 23465 28677 23499 28711
rect 23465 28542 23499 28643
rect 23923 29901 23957 29962
rect 23923 29833 23957 29867
rect 23923 29765 23957 29795
rect 23923 29697 23957 29723
rect 23923 29629 23957 29651
rect 23923 29561 23957 29579
rect 23923 29493 23957 29507
rect 23923 29425 23957 29435
rect 23923 29357 23957 29363
rect 23923 29289 23957 29291
rect 23923 29253 23957 29255
rect 23923 29181 23957 29187
rect 23923 29109 23957 29119
rect 23923 29037 23957 29051
rect 23923 28965 23957 28983
rect 23923 28893 23957 28915
rect 23923 28821 23957 28847
rect 23923 28749 23957 28779
rect 23923 28677 23957 28711
rect 23923 28623 23957 28643
rect 24381 29901 24415 29921
rect 24381 29833 24415 29867
rect 24381 29765 24415 29795
rect 24381 29697 24415 29723
rect 24381 29629 24415 29651
rect 24381 29561 24415 29579
rect 24381 29493 24415 29507
rect 24381 29425 24415 29435
rect 24381 29357 24415 29363
rect 24381 29289 24415 29291
rect 24381 29253 24415 29255
rect 24381 29181 24415 29187
rect 24381 29109 24415 29119
rect 24381 29037 24415 29051
rect 24381 28965 24415 28983
rect 24381 28893 24415 28915
rect 24381 28821 24415 28847
rect 24381 28749 24415 28779
rect 24381 28677 24415 28711
rect 24381 28542 24415 28643
rect 24839 29901 24873 29962
rect 24839 29833 24873 29867
rect 24839 29765 24873 29795
rect 24839 29697 24873 29723
rect 24839 29629 24873 29651
rect 24839 29561 24873 29579
rect 24839 29493 24873 29507
rect 24839 29425 24873 29435
rect 24839 29357 24873 29363
rect 24839 29289 24873 29291
rect 24839 29253 24873 29255
rect 24839 29181 24873 29187
rect 24839 29109 24873 29119
rect 24839 29037 24873 29051
rect 24839 28965 24873 28983
rect 24839 28893 24873 28915
rect 24839 28821 24873 28847
rect 24839 28749 24873 28779
rect 24839 28677 24873 28711
rect 24839 28623 24873 28643
rect 25297 29901 25331 29921
rect 25297 29833 25331 29867
rect 25297 29765 25331 29795
rect 25297 29697 25331 29723
rect 25297 29629 25331 29651
rect 25297 29561 25331 29579
rect 25297 29493 25331 29507
rect 25297 29425 25331 29435
rect 25297 29357 25331 29363
rect 25297 29289 25331 29291
rect 25297 29253 25331 29255
rect 25297 29181 25331 29187
rect 25297 29109 25331 29119
rect 25297 29037 25331 29051
rect 25297 28965 25331 28983
rect 25297 28893 25331 28915
rect 25297 28821 25331 28847
rect 25297 28749 25331 28779
rect 25297 28677 25331 28711
rect 25297 28542 25331 28643
rect 25755 29901 25789 29962
rect 25755 29833 25789 29867
rect 25755 29765 25789 29795
rect 25755 29697 25789 29723
rect 25755 29629 25789 29651
rect 25755 29561 25789 29579
rect 25755 29493 25789 29507
rect 25755 29425 25789 29435
rect 25755 29357 25789 29363
rect 25755 29289 25789 29291
rect 25755 29253 25789 29255
rect 25755 29181 25789 29187
rect 25755 29109 25789 29119
rect 25755 29037 25789 29051
rect 25755 28965 25789 28983
rect 25755 28893 25789 28915
rect 25755 28821 25789 28847
rect 25755 28749 25789 28779
rect 25755 28677 25789 28711
rect 25755 28623 25789 28643
rect 26213 29901 26247 29921
rect 26213 29833 26247 29867
rect 26213 29765 26247 29795
rect 26213 29697 26247 29723
rect 26213 29629 26247 29651
rect 26213 29561 26247 29579
rect 26213 29493 26247 29507
rect 26213 29425 26247 29435
rect 26213 29357 26247 29363
rect 26213 29289 26247 29291
rect 26213 29253 26247 29255
rect 26213 29181 26247 29187
rect 26213 29109 26247 29119
rect 26213 29037 26247 29051
rect 26213 28965 26247 28983
rect 26213 28893 26247 28915
rect 26213 28821 26247 28847
rect 26213 28749 26247 28779
rect 26213 28677 26247 28711
rect 26213 28542 26247 28643
rect 26671 29901 26705 29962
rect 26671 29833 26705 29867
rect 26671 29765 26705 29795
rect 26671 29697 26705 29723
rect 26671 29629 26705 29651
rect 26671 29561 26705 29579
rect 26671 29493 26705 29507
rect 26671 29425 26705 29435
rect 26671 29357 26705 29363
rect 26671 29289 26705 29291
rect 26671 29253 26705 29255
rect 26671 29181 26705 29187
rect 26671 29109 26705 29119
rect 26671 29037 26705 29051
rect 26671 28965 26705 28983
rect 26671 28893 26705 28915
rect 26671 28821 26705 28847
rect 26671 28749 26705 28779
rect 26671 28677 26705 28711
rect 26671 28623 26705 28643
rect 27129 29901 27163 29921
rect 27129 29833 27163 29867
rect 27129 29765 27163 29795
rect 27129 29697 27163 29723
rect 27129 29629 27163 29651
rect 27129 29561 27163 29579
rect 27129 29493 27163 29507
rect 27129 29425 27163 29435
rect 27129 29357 27163 29363
rect 27129 29289 27163 29291
rect 27129 29253 27163 29255
rect 27129 29181 27163 29187
rect 27129 29109 27163 29119
rect 27129 29037 27163 29051
rect 27129 28965 27163 28983
rect 27129 28893 27163 28915
rect 27129 28821 27163 28847
rect 27129 28749 27163 28779
rect 27129 28677 27163 28711
rect 27129 28542 27163 28643
rect 27587 29901 27621 29962
rect 27587 29833 27621 29867
rect 27587 29765 27621 29795
rect 27587 29697 27621 29723
rect 27587 29629 27621 29651
rect 27587 29561 27621 29579
rect 27587 29493 27621 29507
rect 27587 29425 27621 29435
rect 27587 29357 27621 29363
rect 27587 29289 27621 29291
rect 27587 29253 27621 29255
rect 27587 29181 27621 29187
rect 27587 29109 27621 29119
rect 27587 29037 27621 29051
rect 27587 28965 27621 28983
rect 27587 28893 27621 28915
rect 27587 28821 27621 28847
rect 27587 28749 27621 28779
rect 27587 28677 27621 28711
rect 27587 28623 27621 28643
rect 28045 29901 28079 29921
rect 28045 29833 28079 29867
rect 28045 29765 28079 29795
rect 28045 29697 28079 29723
rect 28045 29629 28079 29651
rect 28045 29561 28079 29579
rect 28045 29493 28079 29507
rect 28045 29425 28079 29435
rect 28045 29357 28079 29363
rect 28045 29289 28079 29291
rect 28045 29253 28079 29255
rect 28045 29181 28079 29187
rect 28045 29109 28079 29119
rect 28045 29037 28079 29051
rect 28045 28965 28079 28983
rect 28045 28893 28079 28915
rect 28045 28821 28079 28847
rect 28045 28749 28079 28779
rect 28045 28677 28079 28711
rect 28045 28542 28079 28643
rect 28503 29901 28537 29962
rect 28503 29833 28537 29867
rect 28503 29765 28537 29795
rect 28503 29697 28537 29723
rect 28503 29629 28537 29651
rect 28503 29561 28537 29579
rect 28503 29493 28537 29507
rect 28503 29425 28537 29435
rect 28503 29357 28537 29363
rect 28503 29289 28537 29291
rect 28503 29253 28537 29255
rect 28503 29181 28537 29187
rect 28503 29109 28537 29119
rect 28503 29037 28537 29051
rect 28503 28965 28537 28983
rect 28503 28893 28537 28915
rect 28503 28821 28537 28847
rect 28503 28749 28537 28779
rect 28503 28677 28537 28711
rect 28503 28623 28537 28643
rect 28961 29901 28995 29921
rect 28961 29833 28995 29867
rect 28961 29765 28995 29795
rect 28961 29697 28995 29723
rect 28961 29629 28995 29651
rect 28961 29561 28995 29579
rect 28961 29493 28995 29507
rect 28961 29425 28995 29435
rect 28961 29357 28995 29363
rect 28961 29289 28995 29291
rect 28961 29253 28995 29255
rect 28961 29181 28995 29187
rect 28961 29109 28995 29119
rect 28961 29037 28995 29051
rect 28961 28965 28995 28983
rect 28961 28893 28995 28915
rect 28961 28821 28995 28847
rect 28961 28749 28995 28779
rect 28961 28677 28995 28711
rect 28961 28542 28995 28643
rect 29419 29901 29453 29962
rect 29419 29833 29453 29867
rect 29419 29765 29453 29795
rect 29419 29697 29453 29723
rect 29419 29629 29453 29651
rect 29419 29561 29453 29579
rect 29419 29493 29453 29507
rect 29419 29425 29453 29435
rect 29419 29357 29453 29363
rect 29419 29289 29453 29291
rect 29419 29253 29453 29255
rect 29419 29181 29453 29187
rect 29419 29109 29453 29119
rect 29419 29037 29453 29051
rect 29419 28965 29453 28983
rect 29419 28893 29453 28915
rect 29419 28821 29453 28847
rect 29419 28749 29453 28779
rect 29419 28677 29453 28711
rect 29419 28623 29453 28643
rect 29877 29901 29911 29921
rect 29877 29833 29911 29867
rect 29877 29765 29911 29795
rect 29877 29697 29911 29723
rect 29877 29629 29911 29651
rect 29877 29561 29911 29579
rect 29877 29493 29911 29507
rect 29877 29425 29911 29435
rect 29877 29357 29911 29363
rect 29877 29289 29911 29291
rect 29877 29253 29911 29255
rect 29877 29181 29911 29187
rect 29877 29109 29911 29119
rect 29877 29037 29911 29051
rect 29877 28965 29911 28983
rect 29877 28893 29911 28915
rect 29877 28821 29911 28847
rect 29877 28749 29911 28779
rect 29877 28677 29911 28711
rect 29877 28542 29911 28643
rect 30335 29901 30369 29962
rect 30335 29833 30369 29867
rect 30335 29765 30369 29795
rect 30335 29697 30369 29723
rect 30335 29629 30369 29651
rect 30335 29561 30369 29579
rect 30335 29493 30369 29507
rect 30335 29425 30369 29435
rect 30335 29357 30369 29363
rect 30335 29289 30369 29291
rect 30335 29253 30369 29255
rect 30335 29181 30369 29187
rect 30335 29109 30369 29119
rect 30335 29037 30369 29051
rect 30335 28965 30369 28983
rect 30335 28893 30369 28915
rect 30335 28821 30369 28847
rect 30335 28749 30369 28779
rect 30335 28677 30369 28711
rect 30335 28623 30369 28643
rect 30793 29901 30827 29921
rect 30793 29833 30827 29867
rect 30793 29765 30827 29795
rect 30793 29697 30827 29723
rect 30793 29629 30827 29651
rect 30793 29561 30827 29579
rect 30793 29493 30827 29507
rect 30793 29425 30827 29435
rect 30793 29357 30827 29363
rect 30793 29289 30827 29291
rect 30793 29253 30827 29255
rect 30793 29181 30827 29187
rect 30793 29109 30827 29119
rect 30793 29037 30827 29051
rect 30793 28965 30827 28983
rect 30793 28893 30827 28915
rect 30793 28821 30827 28847
rect 30793 28749 30827 28779
rect 30793 28677 30827 28711
rect 30793 28542 30827 28643
rect 31251 29901 31285 29962
rect 31251 29833 31285 29867
rect 31251 29765 31285 29795
rect 31251 29697 31285 29723
rect 31251 29629 31285 29651
rect 31251 29561 31285 29579
rect 31251 29493 31285 29507
rect 31251 29425 31285 29435
rect 31251 29357 31285 29363
rect 31251 29289 31285 29291
rect 31251 29253 31285 29255
rect 31251 29181 31285 29187
rect 31251 29109 31285 29119
rect 31251 29037 31285 29051
rect 31251 28965 31285 28983
rect 31251 28893 31285 28915
rect 31251 28821 31285 28847
rect 31251 28749 31285 28779
rect 31251 28677 31285 28711
rect 31251 28623 31285 28643
rect 31709 29901 31743 29921
rect 31709 29833 31743 29867
rect 31709 29765 31743 29795
rect 31709 29697 31743 29723
rect 31709 29629 31743 29651
rect 31709 29561 31743 29579
rect 31709 29493 31743 29507
rect 31709 29425 31743 29435
rect 31709 29357 31743 29363
rect 31709 29289 31743 29291
rect 31709 29253 31743 29255
rect 31709 29181 31743 29187
rect 31709 29109 31743 29119
rect 31709 29037 31743 29051
rect 31709 28965 31743 28983
rect 31709 28893 31743 28915
rect 31709 28821 31743 28847
rect 31709 28749 31743 28779
rect 31709 28677 31743 28711
rect 31709 28542 31743 28643
rect 32167 29901 32201 29962
rect 32167 29833 32201 29867
rect 32167 29765 32201 29795
rect 32167 29697 32201 29723
rect 32167 29629 32201 29651
rect 32167 29561 32201 29579
rect 32167 29493 32201 29507
rect 32167 29425 32201 29435
rect 32167 29357 32201 29363
rect 32167 29289 32201 29291
rect 32167 29253 32201 29255
rect 32167 29181 32201 29187
rect 32167 29109 32201 29119
rect 32167 29037 32201 29051
rect 32167 28965 32201 28983
rect 32167 28893 32201 28915
rect 32167 28821 32201 28847
rect 32167 28749 32201 28779
rect 32167 28677 32201 28711
rect 32167 28623 32201 28643
rect 32625 29901 32659 29921
rect 32625 29833 32659 29867
rect 32625 29765 32659 29795
rect 32625 29697 32659 29723
rect 32625 29629 32659 29651
rect 32625 29561 32659 29579
rect 32625 29493 32659 29507
rect 32625 29425 32659 29435
rect 32625 29357 32659 29363
rect 32625 29289 32659 29291
rect 32625 29253 32659 29255
rect 32625 29181 32659 29187
rect 32625 29109 32659 29119
rect 32625 29037 32659 29051
rect 32625 28965 32659 28983
rect 32625 28893 32659 28915
rect 32625 28821 32659 28847
rect 32625 28749 32659 28779
rect 32625 28677 32659 28711
rect 32625 28542 32659 28643
rect 33083 29901 33117 29962
rect 33083 29833 33117 29867
rect 33083 29765 33117 29795
rect 33083 29697 33117 29723
rect 33083 29629 33117 29651
rect 33083 29561 33117 29579
rect 33083 29493 33117 29507
rect 33083 29425 33117 29435
rect 33083 29357 33117 29363
rect 33083 29289 33117 29291
rect 33083 29253 33117 29255
rect 33083 29181 33117 29187
rect 33083 29109 33117 29119
rect 33083 29037 33117 29051
rect 33083 28965 33117 28983
rect 33083 28893 33117 28915
rect 33083 28821 33117 28847
rect 33083 28749 33117 28779
rect 33083 28677 33117 28711
rect 33083 28623 33117 28643
rect 33541 29901 33575 29921
rect 33972 29912 34032 29995
rect 34102 29962 36918 30002
rect 33541 29833 33575 29867
rect 33541 29765 33575 29795
rect 33541 29697 33575 29723
rect 33541 29629 33575 29651
rect 33541 29561 33575 29579
rect 33541 29493 33575 29507
rect 33541 29425 33575 29435
rect 33541 29357 33575 29363
rect 33541 29289 33575 29291
rect 33541 29253 33575 29255
rect 33541 29181 33575 29187
rect 33541 29109 33575 29119
rect 33541 29037 33575 29051
rect 33541 28965 33575 28983
rect 33541 28893 33575 28915
rect 33541 28821 33575 28847
rect 33541 28749 33575 28779
rect 33541 28677 33575 28711
rect 33541 28542 33575 28643
rect 34089 29901 34123 29921
rect 34089 29833 34123 29867
rect 34089 29765 34123 29795
rect 34089 29697 34123 29723
rect 34089 29629 34123 29651
rect 34089 29561 34123 29579
rect 34089 29493 34123 29507
rect 34089 29425 34123 29435
rect 34089 29357 34123 29363
rect 34089 29289 34123 29291
rect 34089 29253 34123 29255
rect 34089 29181 34123 29187
rect 34089 29109 34123 29119
rect 34089 29037 34123 29051
rect 34089 28965 34123 28983
rect 34089 28893 34123 28915
rect 34089 28821 34123 28847
rect 34089 28749 34123 28779
rect 34089 28677 34123 28711
rect 34089 28542 34123 28643
rect 34547 29901 34581 29962
rect 34547 29833 34581 29867
rect 34547 29765 34581 29795
rect 34547 29697 34581 29723
rect 34547 29629 34581 29651
rect 34547 29561 34581 29579
rect 34547 29493 34581 29507
rect 34547 29425 34581 29435
rect 34547 29357 34581 29363
rect 34547 29289 34581 29291
rect 34547 29253 34581 29255
rect 34547 29181 34581 29187
rect 34547 29109 34581 29119
rect 34547 29037 34581 29051
rect 34547 28965 34581 28983
rect 34547 28893 34581 28915
rect 34547 28821 34581 28847
rect 34547 28749 34581 28779
rect 34547 28677 34581 28711
rect 34547 28623 34581 28643
rect 35005 29901 35039 29921
rect 35005 29833 35039 29867
rect 35005 29765 35039 29795
rect 35005 29697 35039 29723
rect 35005 29629 35039 29651
rect 35005 29561 35039 29579
rect 35005 29493 35039 29507
rect 35005 29425 35039 29435
rect 35005 29357 35039 29363
rect 35005 29289 35039 29291
rect 35005 29253 35039 29255
rect 35005 29181 35039 29187
rect 35005 29109 35039 29119
rect 35005 29037 35039 29051
rect 35005 28965 35039 28983
rect 35005 28893 35039 28915
rect 35005 28821 35039 28847
rect 35005 28749 35039 28779
rect 35005 28677 35039 28711
rect 35005 28542 35039 28643
rect 35463 29901 35497 29962
rect 35463 29833 35497 29867
rect 35463 29765 35497 29795
rect 35463 29697 35497 29723
rect 35463 29629 35497 29651
rect 35463 29561 35497 29579
rect 35463 29493 35497 29507
rect 35463 29425 35497 29435
rect 35463 29357 35497 29363
rect 35463 29289 35497 29291
rect 35463 29253 35497 29255
rect 35463 29181 35497 29187
rect 35463 29109 35497 29119
rect 35463 29037 35497 29051
rect 35463 28965 35497 28983
rect 35463 28893 35497 28915
rect 35463 28821 35497 28847
rect 35463 28749 35497 28779
rect 35463 28677 35497 28711
rect 35463 28623 35497 28643
rect 35921 29901 35955 29921
rect 35921 29833 35955 29867
rect 35921 29765 35955 29795
rect 35921 29697 35955 29723
rect 35921 29629 35955 29651
rect 35921 29561 35955 29579
rect 35921 29493 35955 29507
rect 35921 29425 35955 29435
rect 35921 29357 35955 29363
rect 35921 29289 35955 29291
rect 35921 29253 35955 29255
rect 35921 29181 35955 29187
rect 35921 29109 35955 29119
rect 35921 29037 35955 29051
rect 35921 28965 35955 28983
rect 35921 28893 35955 28915
rect 35921 28821 35955 28847
rect 35921 28749 35955 28779
rect 35921 28677 35955 28711
rect 35921 28542 35955 28643
rect 36379 29901 36413 29962
rect 36379 29833 36413 29867
rect 36379 29765 36413 29795
rect 36379 29697 36413 29723
rect 36379 29629 36413 29651
rect 36379 29561 36413 29579
rect 36379 29493 36413 29507
rect 36379 29425 36413 29435
rect 36379 29357 36413 29363
rect 36379 29289 36413 29291
rect 36379 29253 36413 29255
rect 36379 29181 36413 29187
rect 36379 29109 36413 29119
rect 36379 29037 36413 29051
rect 36379 28965 36413 28983
rect 36379 28893 36413 28915
rect 36379 28821 36413 28847
rect 36379 28749 36413 28779
rect 36379 28677 36413 28711
rect 36379 28623 36413 28643
rect 36837 29901 36871 29921
rect 36837 29833 36871 29867
rect 36837 29765 36871 29795
rect 36837 29697 36871 29723
rect 36837 29629 36871 29651
rect 36837 29561 36871 29579
rect 36837 29493 36871 29507
rect 36837 29425 36871 29435
rect 36837 29357 36871 29363
rect 36837 29289 36871 29291
rect 36837 29253 36871 29255
rect 36837 29181 36871 29187
rect 36837 29109 36871 29119
rect 36837 29037 36871 29051
rect 36837 28965 36871 28983
rect 38306 29203 38922 29242
rect 38306 29101 38393 29203
rect 38835 29101 38922 29203
rect 36837 28893 36871 28915
rect 36837 28821 36871 28847
rect 36837 28749 36871 28779
rect 36837 28677 36871 28711
rect 36837 28542 36871 28643
rect 6014 28482 33622 28542
rect 34042 28482 36918 28542
rect 6014 28423 33622 28436
rect 6014 28389 6197 28423
rect 6231 28389 6597 28423
rect 6631 28389 6997 28423
rect 7031 28389 7397 28423
rect 7431 28389 7797 28423
rect 7831 28389 8197 28423
rect 8231 28389 8597 28423
rect 8631 28389 8997 28423
rect 9031 28389 9397 28423
rect 9431 28389 9797 28423
rect 9831 28389 10197 28423
rect 10231 28389 10597 28423
rect 10631 28389 10997 28423
rect 11031 28389 11397 28423
rect 11431 28389 11797 28423
rect 11831 28389 12197 28423
rect 12231 28407 12597 28423
rect 12231 28389 12541 28407
rect 6014 28376 12541 28389
rect 12575 28389 12597 28407
rect 12631 28389 12997 28423
rect 13031 28389 13397 28423
rect 13431 28389 13797 28423
rect 13831 28389 14197 28423
rect 14231 28389 14597 28423
rect 14631 28389 14997 28423
rect 15031 28389 15397 28423
rect 15431 28389 15797 28423
rect 15831 28389 16197 28423
rect 16231 28389 16597 28423
rect 16631 28389 16997 28423
rect 17031 28389 17397 28423
rect 17431 28389 17797 28423
rect 17831 28389 18197 28423
rect 18231 28389 18597 28423
rect 18631 28389 18997 28423
rect 19031 28389 19397 28423
rect 19431 28389 19797 28423
rect 19831 28389 20197 28423
rect 20231 28389 20597 28423
rect 20631 28389 20997 28423
rect 21031 28389 21397 28423
rect 21431 28389 21797 28423
rect 21831 28389 22197 28423
rect 22231 28389 22597 28423
rect 22631 28389 22997 28423
rect 23031 28389 23397 28423
rect 23431 28389 23797 28423
rect 23831 28389 24197 28423
rect 24231 28389 24597 28423
rect 24631 28389 24997 28423
rect 25031 28389 25397 28423
rect 25431 28389 25797 28423
rect 25831 28389 26197 28423
rect 26231 28389 26597 28423
rect 26631 28389 26997 28423
rect 27031 28389 27397 28423
rect 27431 28389 27797 28423
rect 27831 28389 28197 28423
rect 28231 28389 28597 28423
rect 28631 28389 28997 28423
rect 29031 28389 29397 28423
rect 29431 28389 29797 28423
rect 29831 28389 30197 28423
rect 30231 28389 30597 28423
rect 30631 28389 30997 28423
rect 31031 28389 31397 28423
rect 31431 28389 31797 28423
rect 31831 28389 32197 28423
rect 32231 28389 32597 28423
rect 32631 28389 32997 28423
rect 33031 28389 33397 28423
rect 33431 28389 33622 28423
rect 12575 28376 14197 28389
rect 14231 28376 23397 28389
rect 23431 28376 33622 28389
rect 34042 28423 36918 28436
rect 34042 28407 34225 28423
rect 34042 28376 34069 28407
rect 34103 28389 34225 28407
rect 34259 28389 34625 28423
rect 34659 28389 35025 28423
rect 35059 28389 35425 28423
rect 35459 28389 35825 28423
rect 35859 28389 36225 28423
rect 36259 28389 36625 28423
rect 36659 28389 36918 28423
rect 34103 28376 36918 28389
rect 38306 28302 38922 29101
rect 39402 28957 39834 29347
rect 41050 29203 41666 29242
rect 41050 29101 41137 29203
rect 41579 29101 41666 29203
rect 41050 28302 41666 29101
rect 42146 28957 42578 29347
rect 5916 28289 33622 28302
rect 5916 28255 6197 28289
rect 6231 28255 6597 28289
rect 6631 28255 6997 28289
rect 7031 28255 7397 28289
rect 7431 28255 7797 28289
rect 7831 28255 8197 28289
rect 8231 28255 8597 28289
rect 8631 28255 8997 28289
rect 9031 28255 9397 28289
rect 9431 28255 9797 28289
rect 9831 28255 10197 28289
rect 10231 28255 10597 28289
rect 10631 28255 10997 28289
rect 11031 28255 11397 28289
rect 11431 28255 11797 28289
rect 11831 28255 12197 28289
rect 12231 28255 12597 28289
rect 12631 28255 12997 28289
rect 13031 28255 13397 28289
rect 13431 28255 13797 28289
rect 13831 28255 14197 28289
rect 14231 28255 14597 28289
rect 14631 28255 14997 28289
rect 15031 28255 15397 28289
rect 15431 28255 15797 28289
rect 15831 28255 16197 28289
rect 16231 28255 16597 28289
rect 16631 28255 16997 28289
rect 17031 28255 17397 28289
rect 17431 28255 17797 28289
rect 17831 28255 18197 28289
rect 18231 28255 18597 28289
rect 18631 28255 18997 28289
rect 19031 28255 19397 28289
rect 19431 28255 19797 28289
rect 19831 28255 20197 28289
rect 20231 28255 20597 28289
rect 20631 28255 20997 28289
rect 21031 28255 21397 28289
rect 21431 28255 21797 28289
rect 21831 28255 22197 28289
rect 22231 28255 22597 28289
rect 22631 28255 22997 28289
rect 23031 28255 23397 28289
rect 23431 28255 23797 28289
rect 23831 28255 24197 28289
rect 24231 28255 24597 28289
rect 24631 28255 24997 28289
rect 25031 28255 25397 28289
rect 25431 28255 25797 28289
rect 25831 28255 26197 28289
rect 26231 28255 26597 28289
rect 26631 28255 26997 28289
rect 27031 28255 27397 28289
rect 27431 28255 27797 28289
rect 27831 28255 28197 28289
rect 28231 28255 28597 28289
rect 28631 28255 28997 28289
rect 29031 28255 29397 28289
rect 29431 28255 29797 28289
rect 29831 28255 30197 28289
rect 30231 28255 30597 28289
rect 30631 28255 30997 28289
rect 31031 28255 31397 28289
rect 31431 28255 31797 28289
rect 31831 28255 32197 28289
rect 32231 28255 32597 28289
rect 32631 28255 32997 28289
rect 33031 28255 33397 28289
rect 33431 28255 33622 28289
rect 5916 28242 33622 28255
rect 33944 28289 36918 28302
rect 33944 28255 34225 28289
rect 34259 28255 34625 28289
rect 34659 28255 35025 28289
rect 35059 28255 35425 28289
rect 35459 28255 35825 28289
rect 35859 28255 36225 28289
rect 36259 28255 36625 28289
rect 36659 28255 36918 28289
rect 33944 28242 36918 28255
rect 37394 28289 39834 28302
rect 37394 28255 37577 28289
rect 37611 28255 37777 28289
rect 37811 28255 37977 28289
rect 38011 28255 38177 28289
rect 38211 28255 38377 28289
rect 38411 28255 38577 28289
rect 38611 28255 38777 28289
rect 38811 28255 38977 28289
rect 39011 28255 39177 28289
rect 39211 28255 39377 28289
rect 39411 28255 39577 28289
rect 39611 28255 39834 28289
rect 37394 28242 39834 28255
rect 40138 28289 42578 28302
rect 40138 28255 40321 28289
rect 40355 28255 40521 28289
rect 40555 28255 40721 28289
rect 40755 28255 40921 28289
rect 40955 28255 41121 28289
rect 41155 28255 41321 28289
rect 41355 28255 41521 28289
rect 41555 28255 41721 28289
rect 41755 28255 41921 28289
rect 41955 28255 42121 28289
rect 42155 28255 42321 28289
rect 42355 28255 42578 28289
rect 40138 28242 42578 28255
rect 6720 26409 9160 26422
rect 6720 26375 6903 26409
rect 6937 26375 7103 26409
rect 7137 26375 7303 26409
rect 7337 26375 7503 26409
rect 7537 26375 7703 26409
rect 7737 26375 7903 26409
rect 7937 26375 8103 26409
rect 8137 26375 8303 26409
rect 8337 26375 8503 26409
rect 8537 26375 8703 26409
rect 8737 26375 8903 26409
rect 8937 26375 9160 26409
rect 6720 26362 9160 26375
rect 9444 26409 15166 26422
rect 9444 26375 9725 26409
rect 9759 26375 10125 26409
rect 10159 26375 10525 26409
rect 10559 26375 10925 26409
rect 10959 26375 11325 26409
rect 11359 26375 11725 26409
rect 11759 26375 12125 26409
rect 12159 26375 12525 26409
rect 12559 26375 12925 26409
rect 12959 26375 13325 26409
rect 13359 26375 13725 26409
rect 13759 26375 14125 26409
rect 14159 26375 14525 26409
rect 14559 26375 14925 26409
rect 14959 26375 15166 26409
rect 9444 26362 15166 26375
rect 15424 26409 22592 26422
rect 15424 26375 15607 26409
rect 15641 26375 16007 26409
rect 16041 26375 16407 26409
rect 16441 26375 16807 26409
rect 16841 26375 17207 26409
rect 17241 26375 17607 26409
rect 17641 26375 18007 26409
rect 18041 26375 18407 26409
rect 18441 26375 18807 26409
rect 18841 26375 19207 26409
rect 19241 26375 19607 26409
rect 19641 26375 20007 26409
rect 20041 26375 20407 26409
rect 20441 26375 20807 26409
rect 20841 26375 21207 26409
rect 21241 26375 21607 26409
rect 21641 26375 22007 26409
rect 22041 26375 22407 26409
rect 22441 26375 22592 26409
rect 15424 26362 22592 26375
rect 22870 26409 27148 26422
rect 22870 26375 23151 26409
rect 23185 26375 23551 26409
rect 23585 26375 23951 26409
rect 23985 26375 24351 26409
rect 24385 26375 24751 26409
rect 24785 26375 25151 26409
rect 25185 26375 25551 26409
rect 25585 26375 25951 26409
rect 25985 26375 26351 26409
rect 26385 26375 26751 26409
rect 26785 26375 27148 26409
rect 22870 26362 27148 26375
rect 28260 26409 38980 26422
rect 28260 26375 28443 26409
rect 28477 26375 28643 26409
rect 28677 26375 28843 26409
rect 28877 26375 29043 26409
rect 29077 26375 29243 26409
rect 29277 26375 29443 26409
rect 29477 26375 29643 26409
rect 29677 26375 29843 26409
rect 29877 26375 30043 26409
rect 30077 26375 30243 26409
rect 30277 26375 30443 26409
rect 30477 26375 30643 26409
rect 30677 26375 30843 26409
rect 30877 26375 31043 26409
rect 31077 26375 31243 26409
rect 31277 26375 31443 26409
rect 31477 26375 31643 26409
rect 31677 26375 31843 26409
rect 31877 26375 32043 26409
rect 32077 26375 32243 26409
rect 32277 26375 32443 26409
rect 32477 26375 32643 26409
rect 32677 26375 32843 26409
rect 32877 26375 33043 26409
rect 33077 26375 33243 26409
rect 33277 26375 33443 26409
rect 33477 26375 33643 26409
rect 33677 26375 33843 26409
rect 33877 26375 34043 26409
rect 34077 26375 34243 26409
rect 34277 26375 34443 26409
rect 34477 26375 34643 26409
rect 34677 26375 34843 26409
rect 34877 26375 35043 26409
rect 35077 26375 35243 26409
rect 35277 26375 35443 26409
rect 35477 26375 35643 26409
rect 35677 26375 35843 26409
rect 35877 26375 36043 26409
rect 36077 26375 36243 26409
rect 36277 26375 36443 26409
rect 36477 26375 36643 26409
rect 36677 26375 36843 26409
rect 36877 26375 37043 26409
rect 37077 26375 37243 26409
rect 37277 26375 37443 26409
rect 37477 26375 37643 26409
rect 37677 26375 37843 26409
rect 37877 26375 38043 26409
rect 38077 26375 38243 26409
rect 38277 26375 38443 26409
rect 38477 26375 38643 26409
rect 38677 26375 38843 26409
rect 38877 26375 38980 26409
rect 28260 26362 38980 26375
rect 39746 26409 42186 26422
rect 39746 26375 39929 26409
rect 39963 26375 40129 26409
rect 40163 26375 40329 26409
rect 40363 26375 40529 26409
rect 40563 26375 40729 26409
rect 40763 26375 40929 26409
rect 40963 26375 41129 26409
rect 41163 26375 41329 26409
rect 41363 26375 41529 26409
rect 41563 26375 41729 26409
rect 41763 26375 41929 26409
rect 41963 26375 42186 26409
rect 39746 26362 42186 26375
rect 9472 26269 9532 26362
rect 10520 26319 10680 26362
rect 10520 26285 10585 26319
rect 10619 26285 10680 26319
rect 10520 26282 10680 26285
rect 11820 26319 11980 26362
rect 11820 26285 11885 26319
rect 11919 26285 11980 26319
rect 11820 26282 11980 26285
rect 13120 26319 13280 26362
rect 13120 26285 13185 26319
rect 13219 26285 13280 26319
rect 13120 26282 13280 26285
rect 9472 26235 9485 26269
rect 9519 26235 9532 26269
rect 9472 26152 9532 26235
rect 9602 26202 15166 26242
rect 22968 26231 27148 26262
rect 22968 26202 26157 26231
rect 7632 25443 8248 25482
rect 7632 25341 7719 25443
rect 8161 25341 8248 25443
rect 7632 24542 8248 25341
rect 8728 25197 9160 25587
rect 9589 26141 9623 26161
rect 9589 26073 9623 26107
rect 9589 26005 9623 26035
rect 9589 25937 9623 25963
rect 9589 25869 9623 25891
rect 9589 25801 9623 25819
rect 9589 25733 9623 25747
rect 9589 25665 9623 25675
rect 9589 25597 9623 25603
rect 9589 25529 9623 25531
rect 9589 25493 9623 25495
rect 9589 25421 9623 25427
rect 9589 25349 9623 25359
rect 9589 25277 9623 25291
rect 9589 25205 9623 25223
rect 9589 25133 9623 25155
rect 9589 25061 9623 25087
rect 9589 24989 9623 25019
rect 9589 24917 9623 24951
rect 9589 24782 9623 24883
rect 10047 26141 10081 26202
rect 10047 26073 10081 26107
rect 10047 26005 10081 26035
rect 10047 25937 10081 25963
rect 10047 25869 10081 25891
rect 10047 25801 10081 25819
rect 10047 25733 10081 25747
rect 10047 25665 10081 25675
rect 10047 25597 10081 25603
rect 10047 25529 10081 25531
rect 10047 25493 10081 25495
rect 10047 25421 10081 25427
rect 10047 25349 10081 25359
rect 10047 25277 10081 25291
rect 10047 25205 10081 25223
rect 10047 25133 10081 25155
rect 10047 25061 10081 25087
rect 10047 24989 10081 25019
rect 10047 24917 10081 24951
rect 10047 24863 10081 24883
rect 10505 26141 10539 26161
rect 10505 26073 10539 26107
rect 10505 26005 10539 26035
rect 10505 25937 10539 25963
rect 10505 25869 10539 25891
rect 10505 25801 10539 25819
rect 10505 25733 10539 25747
rect 10505 25665 10539 25675
rect 10505 25597 10539 25603
rect 10505 25529 10539 25531
rect 10505 25493 10539 25495
rect 10505 25421 10539 25427
rect 10505 25349 10539 25359
rect 10505 25277 10539 25291
rect 10505 25205 10539 25223
rect 10505 25133 10539 25155
rect 10505 25061 10539 25087
rect 10505 24989 10539 25019
rect 10505 24917 10539 24951
rect 10505 24782 10539 24883
rect 10963 26141 10997 26202
rect 10963 26073 10997 26107
rect 10963 26005 10997 26035
rect 10963 25937 10997 25963
rect 10963 25869 10997 25891
rect 10963 25801 10997 25819
rect 10963 25733 10997 25747
rect 10963 25665 10997 25675
rect 10963 25597 10997 25603
rect 10963 25529 10997 25531
rect 10963 25493 10997 25495
rect 10963 25421 10997 25427
rect 10963 25349 10997 25359
rect 10963 25277 10997 25291
rect 10963 25205 10997 25223
rect 10963 25133 10997 25155
rect 10963 25061 10997 25087
rect 10963 24989 10997 25019
rect 10963 24917 10997 24951
rect 10963 24863 10997 24883
rect 11421 26141 11455 26161
rect 11421 26073 11455 26107
rect 11421 26005 11455 26035
rect 11421 25937 11455 25963
rect 11421 25869 11455 25891
rect 11421 25801 11455 25819
rect 11421 25733 11455 25747
rect 11421 25665 11455 25675
rect 11421 25597 11455 25603
rect 11421 25529 11455 25531
rect 11421 25493 11455 25495
rect 11421 25421 11455 25427
rect 11421 25349 11455 25359
rect 11421 25277 11455 25291
rect 11421 25205 11455 25223
rect 11421 25133 11455 25155
rect 11421 25061 11455 25087
rect 11421 24989 11455 25019
rect 11421 24917 11455 24951
rect 11421 24782 11455 24883
rect 11879 26141 11913 26202
rect 11879 26073 11913 26107
rect 11879 26005 11913 26035
rect 11879 25937 11913 25963
rect 11879 25869 11913 25891
rect 11879 25801 11913 25819
rect 11879 25733 11913 25747
rect 11879 25665 11913 25675
rect 11879 25597 11913 25603
rect 11879 25529 11913 25531
rect 11879 25493 11913 25495
rect 11879 25421 11913 25427
rect 11879 25349 11913 25359
rect 11879 25277 11913 25291
rect 11879 25205 11913 25223
rect 11879 25133 11913 25155
rect 11879 25061 11913 25087
rect 11879 24989 11913 25019
rect 11879 24917 11913 24951
rect 11879 24863 11913 24883
rect 12337 26141 12371 26161
rect 12337 26073 12371 26107
rect 12337 26005 12371 26035
rect 12337 25937 12371 25963
rect 12337 25869 12371 25891
rect 12337 25801 12371 25819
rect 12337 25733 12371 25747
rect 12337 25665 12371 25675
rect 12337 25597 12371 25603
rect 12337 25529 12371 25531
rect 12337 25493 12371 25495
rect 12337 25421 12371 25427
rect 12337 25349 12371 25359
rect 12337 25277 12371 25291
rect 12337 25205 12371 25223
rect 12337 25133 12371 25155
rect 12337 25061 12371 25087
rect 12337 24989 12371 25019
rect 12337 24917 12371 24951
rect 12337 24782 12371 24883
rect 12795 26141 12829 26202
rect 12795 26073 12829 26107
rect 12795 26005 12829 26035
rect 12795 25937 12829 25963
rect 12795 25869 12829 25891
rect 12795 25801 12829 25819
rect 12795 25733 12829 25747
rect 12795 25665 12829 25675
rect 12795 25597 12829 25603
rect 12795 25529 12829 25531
rect 12795 25493 12829 25495
rect 12795 25421 12829 25427
rect 12795 25349 12829 25359
rect 12795 25277 12829 25291
rect 12795 25205 12829 25223
rect 12795 25133 12829 25155
rect 12795 25061 12829 25087
rect 12795 24989 12829 25019
rect 12795 24917 12829 24951
rect 12795 24863 12829 24883
rect 13253 26141 13287 26161
rect 13253 26073 13287 26107
rect 13253 26005 13287 26035
rect 13253 25937 13287 25963
rect 13253 25869 13287 25891
rect 13253 25801 13287 25819
rect 13253 25733 13287 25747
rect 13253 25665 13287 25675
rect 13253 25597 13287 25603
rect 13253 25529 13287 25531
rect 13253 25493 13287 25495
rect 13253 25421 13287 25427
rect 13253 25349 13287 25359
rect 13253 25277 13287 25291
rect 13253 25205 13287 25223
rect 13253 25133 13287 25155
rect 13253 25061 13287 25087
rect 13253 24989 13287 25019
rect 13253 24917 13287 24951
rect 13253 24782 13287 24883
rect 13711 26141 13745 26202
rect 13711 26073 13745 26107
rect 13711 26005 13745 26035
rect 13711 25937 13745 25963
rect 13711 25869 13745 25891
rect 13711 25801 13745 25819
rect 13711 25733 13745 25747
rect 13711 25665 13745 25675
rect 13711 25597 13745 25603
rect 13711 25529 13745 25531
rect 13711 25493 13745 25495
rect 13711 25421 13745 25427
rect 13711 25349 13745 25359
rect 13711 25277 13745 25291
rect 13711 25205 13745 25223
rect 13711 25133 13745 25155
rect 13711 25061 13745 25087
rect 13711 24989 13745 25019
rect 13711 24917 13745 24951
rect 13711 24863 13745 24883
rect 14169 26141 14203 26161
rect 14169 26073 14203 26107
rect 14169 26005 14203 26035
rect 14169 25937 14203 25963
rect 14169 25869 14203 25891
rect 14169 25801 14203 25819
rect 14169 25733 14203 25747
rect 14169 25665 14203 25675
rect 14169 25597 14203 25603
rect 14169 25529 14203 25531
rect 14169 25493 14203 25495
rect 14169 25421 14203 25427
rect 14169 25349 14203 25359
rect 14169 25277 14203 25291
rect 14169 25205 14203 25223
rect 14169 25133 14203 25155
rect 14169 25061 14203 25087
rect 14169 24989 14203 25019
rect 14169 24917 14203 24951
rect 14169 24782 14203 24883
rect 14627 26141 14661 26202
rect 14627 26073 14661 26107
rect 14627 26005 14661 26035
rect 14627 25937 14661 25963
rect 14627 25869 14661 25891
rect 14627 25801 14661 25819
rect 14627 25733 14661 25747
rect 14627 25665 14661 25675
rect 14627 25597 14661 25603
rect 14627 25529 14661 25531
rect 14627 25493 14661 25495
rect 14627 25421 14661 25427
rect 14627 25349 14661 25359
rect 14627 25277 14661 25291
rect 14627 25205 14661 25223
rect 14627 25133 14661 25155
rect 14627 25061 14661 25087
rect 14627 24989 14661 25019
rect 14627 24917 14661 24951
rect 14627 24863 14661 24883
rect 15085 26141 15119 26161
rect 15085 26073 15119 26107
rect 15085 26005 15119 26035
rect 15085 25937 15119 25963
rect 23437 25916 23471 26202
rect 24353 25916 24387 26202
rect 25269 25916 25303 26202
rect 26191 26202 27148 26231
rect 26191 26197 26219 26202
rect 26185 25916 26219 26197
rect 27101 25916 27135 26202
rect 28286 26076 38954 26096
rect 28286 26042 28306 26076
rect 28340 26042 28396 26076
rect 28430 26061 28486 26076
rect 28520 26061 28576 26076
rect 28610 26061 28666 26076
rect 28700 26061 28756 26076
rect 28790 26061 28846 26076
rect 28880 26061 28936 26076
rect 28970 26061 29026 26076
rect 29060 26061 29116 26076
rect 29150 26061 29206 26076
rect 29240 26061 29296 26076
rect 29330 26061 29386 26076
rect 29420 26061 29476 26076
rect 28450 26042 28486 26061
rect 28540 26042 28576 26061
rect 28630 26042 28666 26061
rect 28720 26042 28756 26061
rect 28810 26042 28846 26061
rect 28900 26042 28936 26061
rect 28990 26042 29026 26061
rect 29080 26042 29116 26061
rect 29170 26042 29206 26061
rect 29260 26042 29296 26061
rect 29350 26042 29386 26061
rect 29440 26042 29476 26061
rect 29510 26042 29646 26076
rect 29680 26042 29736 26076
rect 29770 26061 29826 26076
rect 29860 26061 29916 26076
rect 29950 26061 30006 26076
rect 30040 26061 30096 26076
rect 30130 26061 30186 26076
rect 30220 26061 30276 26076
rect 30310 26061 30366 26076
rect 30400 26061 30456 26076
rect 30490 26061 30546 26076
rect 30580 26061 30636 26076
rect 30670 26061 30726 26076
rect 30760 26061 30816 26076
rect 29790 26042 29826 26061
rect 29880 26042 29916 26061
rect 29970 26042 30006 26061
rect 30060 26042 30096 26061
rect 30150 26042 30186 26061
rect 30240 26042 30276 26061
rect 30330 26042 30366 26061
rect 30420 26042 30456 26061
rect 30510 26042 30546 26061
rect 30600 26042 30636 26061
rect 30690 26042 30726 26061
rect 30780 26042 30816 26061
rect 30850 26042 30986 26076
rect 31020 26042 31076 26076
rect 31110 26061 31166 26076
rect 31200 26061 31256 26076
rect 31290 26061 31346 26076
rect 31380 26061 31436 26076
rect 31470 26061 31526 26076
rect 31560 26061 31616 26076
rect 31650 26061 31706 26076
rect 31740 26061 31796 26076
rect 31830 26061 31886 26076
rect 31920 26061 31976 26076
rect 32010 26061 32066 26076
rect 32100 26061 32156 26076
rect 31130 26042 31166 26061
rect 31220 26042 31256 26061
rect 31310 26042 31346 26061
rect 31400 26042 31436 26061
rect 31490 26042 31526 26061
rect 31580 26042 31616 26061
rect 31670 26042 31706 26061
rect 31760 26042 31796 26061
rect 31850 26042 31886 26061
rect 31940 26042 31976 26061
rect 32030 26042 32066 26061
rect 32120 26042 32156 26061
rect 32190 26042 32326 26076
rect 32360 26042 32416 26076
rect 32450 26061 32506 26076
rect 32540 26061 32596 26076
rect 32630 26061 32686 26076
rect 32720 26061 32776 26076
rect 32810 26061 32866 26076
rect 32900 26061 32956 26076
rect 32990 26061 33046 26076
rect 33080 26061 33136 26076
rect 33170 26061 33226 26076
rect 33260 26061 33316 26076
rect 33350 26061 33406 26076
rect 33440 26061 33496 26076
rect 32470 26042 32506 26061
rect 32560 26042 32596 26061
rect 32650 26042 32686 26061
rect 32740 26042 32776 26061
rect 32830 26042 32866 26061
rect 32920 26042 32956 26061
rect 33010 26042 33046 26061
rect 33100 26042 33136 26061
rect 33190 26042 33226 26061
rect 33280 26042 33316 26061
rect 33370 26042 33406 26061
rect 33460 26042 33496 26061
rect 33530 26042 33666 26076
rect 33700 26042 33756 26076
rect 33790 26061 33846 26076
rect 33880 26061 33936 26076
rect 33970 26061 34026 26076
rect 34060 26061 34116 26076
rect 34150 26061 34206 26076
rect 34240 26061 34296 26076
rect 34330 26061 34386 26076
rect 34420 26061 34476 26076
rect 34510 26061 34566 26076
rect 34600 26061 34656 26076
rect 34690 26061 34746 26076
rect 34780 26061 34836 26076
rect 33810 26042 33846 26061
rect 33900 26042 33936 26061
rect 33990 26042 34026 26061
rect 34080 26042 34116 26061
rect 34170 26042 34206 26061
rect 34260 26042 34296 26061
rect 34350 26042 34386 26061
rect 34440 26042 34476 26061
rect 34530 26042 34566 26061
rect 34620 26042 34656 26061
rect 34710 26042 34746 26061
rect 34800 26042 34836 26061
rect 34870 26042 35006 26076
rect 35040 26042 35096 26076
rect 35130 26061 35186 26076
rect 35220 26061 35276 26076
rect 35310 26061 35366 26076
rect 35400 26061 35456 26076
rect 35490 26061 35546 26076
rect 35580 26061 35636 26076
rect 35670 26061 35726 26076
rect 35760 26061 35816 26076
rect 35850 26061 35906 26076
rect 35940 26061 35996 26076
rect 36030 26061 36086 26076
rect 36120 26061 36176 26076
rect 35150 26042 35186 26061
rect 35240 26042 35276 26061
rect 35330 26042 35366 26061
rect 35420 26042 35456 26061
rect 35510 26042 35546 26061
rect 35600 26042 35636 26061
rect 35690 26042 35726 26061
rect 35780 26042 35816 26061
rect 35870 26042 35906 26061
rect 35960 26042 35996 26061
rect 36050 26042 36086 26061
rect 36140 26042 36176 26061
rect 36210 26042 36346 26076
rect 36380 26042 36436 26076
rect 36470 26061 36526 26076
rect 36560 26061 36616 26076
rect 36650 26061 36706 26076
rect 36740 26061 36796 26076
rect 36830 26061 36886 26076
rect 36920 26061 36976 26076
rect 37010 26061 37066 26076
rect 37100 26061 37156 26076
rect 37190 26061 37246 26076
rect 37280 26061 37336 26076
rect 37370 26061 37426 26076
rect 37460 26061 37516 26076
rect 36490 26042 36526 26061
rect 36580 26042 36616 26061
rect 36670 26042 36706 26061
rect 36760 26042 36796 26061
rect 36850 26042 36886 26061
rect 36940 26042 36976 26061
rect 37030 26042 37066 26061
rect 37120 26042 37156 26061
rect 37210 26042 37246 26061
rect 37300 26042 37336 26061
rect 37390 26042 37426 26061
rect 37480 26042 37516 26061
rect 37550 26042 37686 26076
rect 37720 26042 37776 26076
rect 37810 26061 37866 26076
rect 37900 26061 37956 26076
rect 37990 26061 38046 26076
rect 38080 26061 38136 26076
rect 38170 26061 38226 26076
rect 38260 26061 38316 26076
rect 38350 26061 38406 26076
rect 38440 26061 38496 26076
rect 38530 26061 38586 26076
rect 38620 26061 38676 26076
rect 38710 26061 38766 26076
rect 38800 26061 38856 26076
rect 37830 26042 37866 26061
rect 37920 26042 37956 26061
rect 38010 26042 38046 26061
rect 38100 26042 38136 26061
rect 38190 26042 38226 26061
rect 38280 26042 38316 26061
rect 38370 26042 38406 26061
rect 38460 26042 38496 26061
rect 38550 26042 38586 26061
rect 38640 26042 38676 26061
rect 38730 26042 38766 26061
rect 38820 26042 38856 26061
rect 38890 26042 38954 26076
rect 28286 26038 28416 26042
rect 28286 26004 28320 26038
rect 28354 26027 28416 26038
rect 28450 26027 28506 26042
rect 28540 26027 28596 26042
rect 28630 26027 28686 26042
rect 28720 26027 28776 26042
rect 28810 26027 28866 26042
rect 28900 26027 28956 26042
rect 28990 26027 29046 26042
rect 29080 26027 29136 26042
rect 29170 26027 29226 26042
rect 29260 26027 29316 26042
rect 29350 26027 29406 26042
rect 29440 26038 29756 26042
rect 29440 26027 29507 26038
rect 28354 26004 29507 26027
rect 29541 26004 29660 26038
rect 29694 26027 29756 26038
rect 29790 26027 29846 26042
rect 29880 26027 29936 26042
rect 29970 26027 30026 26042
rect 30060 26027 30116 26042
rect 30150 26027 30206 26042
rect 30240 26027 30296 26042
rect 30330 26027 30386 26042
rect 30420 26027 30476 26042
rect 30510 26027 30566 26042
rect 30600 26027 30656 26042
rect 30690 26027 30746 26042
rect 30780 26038 31096 26042
rect 30780 26027 30847 26038
rect 29694 26004 30847 26027
rect 30881 26004 31000 26038
rect 31034 26027 31096 26038
rect 31130 26027 31186 26042
rect 31220 26027 31276 26042
rect 31310 26027 31366 26042
rect 31400 26027 31456 26042
rect 31490 26027 31546 26042
rect 31580 26027 31636 26042
rect 31670 26027 31726 26042
rect 31760 26027 31816 26042
rect 31850 26027 31906 26042
rect 31940 26027 31996 26042
rect 32030 26027 32086 26042
rect 32120 26038 32436 26042
rect 32120 26027 32187 26038
rect 31034 26004 32187 26027
rect 32221 26004 32340 26038
rect 32374 26027 32436 26038
rect 32470 26027 32526 26042
rect 32560 26027 32616 26042
rect 32650 26027 32706 26042
rect 32740 26027 32796 26042
rect 32830 26027 32886 26042
rect 32920 26027 32976 26042
rect 33010 26027 33066 26042
rect 33100 26027 33156 26042
rect 33190 26027 33246 26042
rect 33280 26027 33336 26042
rect 33370 26027 33426 26042
rect 33460 26038 33776 26042
rect 33460 26027 33527 26038
rect 32374 26004 33527 26027
rect 33561 26004 33680 26038
rect 33714 26027 33776 26038
rect 33810 26027 33866 26042
rect 33900 26027 33956 26042
rect 33990 26027 34046 26042
rect 34080 26027 34136 26042
rect 34170 26027 34226 26042
rect 34260 26027 34316 26042
rect 34350 26027 34406 26042
rect 34440 26027 34496 26042
rect 34530 26027 34586 26042
rect 34620 26027 34676 26042
rect 34710 26027 34766 26042
rect 34800 26038 35116 26042
rect 34800 26027 34867 26038
rect 33714 26004 34867 26027
rect 34901 26004 35020 26038
rect 35054 26027 35116 26038
rect 35150 26027 35206 26042
rect 35240 26027 35296 26042
rect 35330 26027 35386 26042
rect 35420 26027 35476 26042
rect 35510 26027 35566 26042
rect 35600 26027 35656 26042
rect 35690 26027 35746 26042
rect 35780 26027 35836 26042
rect 35870 26027 35926 26042
rect 35960 26027 36016 26042
rect 36050 26027 36106 26042
rect 36140 26038 36456 26042
rect 36140 26027 36207 26038
rect 35054 26004 36207 26027
rect 36241 26004 36360 26038
rect 36394 26027 36456 26038
rect 36490 26027 36546 26042
rect 36580 26027 36636 26042
rect 36670 26027 36726 26042
rect 36760 26027 36816 26042
rect 36850 26027 36906 26042
rect 36940 26027 36996 26042
rect 37030 26027 37086 26042
rect 37120 26027 37176 26042
rect 37210 26027 37266 26042
rect 37300 26027 37356 26042
rect 37390 26027 37446 26042
rect 37480 26038 37796 26042
rect 37480 26027 37547 26038
rect 36394 26004 37547 26027
rect 37581 26004 37700 26038
rect 37734 26027 37796 26038
rect 37830 26027 37886 26042
rect 37920 26027 37976 26042
rect 38010 26027 38066 26042
rect 38100 26027 38156 26042
rect 38190 26027 38246 26042
rect 38280 26027 38336 26042
rect 38370 26027 38426 26042
rect 38460 26027 38516 26042
rect 38550 26027 38606 26042
rect 38640 26027 38696 26042
rect 38730 26027 38786 26042
rect 38820 26038 38954 26042
rect 38820 26027 38887 26038
rect 37734 26004 38887 26027
rect 38921 26004 38954 26038
rect 28286 25997 38954 26004
rect 28286 25948 28385 25997
rect 15085 25869 15119 25891
rect 15085 25801 15119 25819
rect 15085 25733 15119 25747
rect 15085 25665 15119 25675
rect 15085 25597 15119 25603
rect 15085 25529 15119 25531
rect 15085 25493 15119 25495
rect 15085 25421 15119 25427
rect 15085 25349 15119 25359
rect 15085 25277 15119 25291
rect 15085 25205 15119 25223
rect 22980 25889 23014 25916
rect 23437 25898 23472 25916
rect 22980 25817 23014 25835
rect 22980 25745 23014 25767
rect 22980 25673 23014 25699
rect 22980 25601 23014 25631
rect 22980 25529 23014 25563
rect 22980 25461 23014 25495
rect 22980 25393 23014 25423
rect 22980 25325 23014 25351
rect 22980 25257 23014 25279
rect 22980 25189 23014 25207
rect 15085 25133 15119 25155
rect 15085 25061 15119 25087
rect 22979 25135 22980 25166
rect 22979 25108 23014 25135
rect 23438 25889 23472 25898
rect 23438 25817 23472 25835
rect 23438 25745 23472 25767
rect 23438 25673 23472 25699
rect 23438 25601 23472 25631
rect 23438 25529 23472 25563
rect 23438 25461 23472 25495
rect 23438 25393 23472 25423
rect 23438 25325 23472 25351
rect 23438 25257 23472 25279
rect 23438 25189 23472 25207
rect 23896 25889 23930 25916
rect 24353 25898 24388 25916
rect 23896 25817 23930 25835
rect 23896 25745 23930 25767
rect 23896 25673 23930 25699
rect 23896 25601 23930 25631
rect 23896 25529 23930 25563
rect 23896 25461 23930 25495
rect 23896 25393 23930 25423
rect 23896 25325 23930 25351
rect 23896 25257 23930 25279
rect 23896 25189 23930 25207
rect 23438 25108 23472 25135
rect 23895 25135 23896 25166
rect 23895 25108 23930 25135
rect 24354 25889 24388 25898
rect 24354 25817 24388 25835
rect 24354 25745 24388 25767
rect 24354 25673 24388 25699
rect 24354 25601 24388 25631
rect 24354 25529 24388 25563
rect 24354 25461 24388 25495
rect 24354 25393 24388 25423
rect 24354 25325 24388 25351
rect 24354 25257 24388 25279
rect 24354 25189 24388 25207
rect 24812 25889 24846 25916
rect 25269 25898 25304 25916
rect 24812 25817 24846 25835
rect 24812 25745 24846 25767
rect 24812 25673 24846 25699
rect 24812 25601 24846 25631
rect 24812 25529 24846 25563
rect 24812 25461 24846 25495
rect 24812 25393 24846 25423
rect 24812 25325 24846 25351
rect 24812 25257 24846 25279
rect 24812 25189 24846 25207
rect 24354 25108 24388 25135
rect 24811 25135 24812 25166
rect 24811 25108 24846 25135
rect 25270 25889 25304 25898
rect 25270 25817 25304 25835
rect 25270 25745 25304 25767
rect 25270 25673 25304 25699
rect 25270 25601 25304 25631
rect 25270 25529 25304 25563
rect 25270 25461 25304 25495
rect 25270 25393 25304 25423
rect 25270 25325 25304 25351
rect 25270 25257 25304 25279
rect 25270 25189 25304 25207
rect 25728 25889 25762 25916
rect 26185 25898 26220 25916
rect 25728 25817 25762 25835
rect 25728 25745 25762 25767
rect 25728 25673 25762 25699
rect 25728 25601 25762 25631
rect 25728 25529 25762 25563
rect 25728 25461 25762 25495
rect 25728 25393 25762 25423
rect 25728 25325 25762 25351
rect 25728 25257 25762 25279
rect 25728 25189 25762 25207
rect 25270 25108 25304 25135
rect 25727 25135 25728 25166
rect 25727 25108 25762 25135
rect 26186 25889 26220 25898
rect 26186 25817 26220 25835
rect 26186 25745 26220 25767
rect 26186 25673 26220 25699
rect 26186 25601 26220 25631
rect 26186 25529 26220 25563
rect 26186 25461 26220 25495
rect 26186 25393 26220 25423
rect 26186 25325 26220 25351
rect 26186 25257 26220 25279
rect 26186 25189 26220 25207
rect 26644 25889 26678 25916
rect 27101 25898 27136 25916
rect 26644 25817 26678 25835
rect 26644 25745 26678 25767
rect 26644 25673 26678 25699
rect 26644 25601 26678 25631
rect 26644 25529 26678 25563
rect 26644 25461 26678 25495
rect 26644 25393 26678 25423
rect 26644 25325 26678 25351
rect 26644 25257 26678 25279
rect 26644 25189 26678 25207
rect 26186 25108 26220 25135
rect 26643 25135 26644 25166
rect 26643 25108 26678 25135
rect 27102 25889 27136 25898
rect 27102 25817 27136 25835
rect 27102 25745 27136 25767
rect 27102 25673 27136 25699
rect 27102 25601 27136 25631
rect 27102 25529 27136 25563
rect 27102 25461 27136 25495
rect 27102 25393 27136 25423
rect 27102 25325 27136 25351
rect 27102 25257 27136 25279
rect 27102 25189 27136 25207
rect 27102 25108 27136 25135
rect 28286 25914 28320 25948
rect 28354 25914 28385 25948
rect 29475 25948 29725 25997
rect 28286 25858 28385 25914
rect 28286 25824 28320 25858
rect 28354 25824 28385 25858
rect 28286 25768 28385 25824
rect 28286 25734 28320 25768
rect 28354 25734 28385 25768
rect 28286 25678 28385 25734
rect 28286 25644 28320 25678
rect 28354 25644 28385 25678
rect 28286 25588 28385 25644
rect 28286 25554 28320 25588
rect 28354 25554 28385 25588
rect 28286 25498 28385 25554
rect 28286 25464 28320 25498
rect 28354 25464 28385 25498
rect 28286 25408 28385 25464
rect 28286 25374 28320 25408
rect 28354 25374 28385 25408
rect 28286 25318 28385 25374
rect 28286 25284 28320 25318
rect 28354 25284 28385 25318
rect 28286 25228 28385 25284
rect 28286 25194 28320 25228
rect 28354 25194 28385 25228
rect 28286 25138 28385 25194
rect 22979 25042 23013 25108
rect 23895 25042 23929 25108
rect 24811 25042 24845 25108
rect 25727 25042 25761 25108
rect 26643 25042 26677 25108
rect 28286 25104 28320 25138
rect 28354 25104 28385 25138
rect 28286 25048 28385 25104
rect 15085 24989 15119 25019
rect 22968 25007 27148 25042
rect 22968 24982 23397 25007
rect 23431 24982 27148 25007
rect 28286 25014 28320 25048
rect 28354 25014 28385 25048
rect 15085 24917 15119 24951
rect 15085 24782 15119 24883
rect 28286 24958 28385 25014
rect 28449 25916 29411 25933
rect 28449 25882 28470 25916
rect 28504 25882 28560 25916
rect 28594 25914 28650 25916
rect 28684 25914 28740 25916
rect 28774 25914 28830 25916
rect 28864 25914 28920 25916
rect 28954 25914 29010 25916
rect 29044 25914 29100 25916
rect 29134 25914 29190 25916
rect 29224 25914 29280 25916
rect 29314 25914 29370 25916
rect 28614 25882 28650 25914
rect 28704 25882 28740 25914
rect 28794 25882 28830 25914
rect 28884 25882 28920 25914
rect 28974 25882 29010 25914
rect 29064 25882 29100 25914
rect 29154 25882 29190 25914
rect 29244 25882 29280 25914
rect 29334 25882 29370 25914
rect 29404 25882 29411 25916
rect 28449 25880 28580 25882
rect 28614 25880 28670 25882
rect 28704 25880 28760 25882
rect 28794 25880 28850 25882
rect 28884 25880 28940 25882
rect 28974 25880 29030 25882
rect 29064 25880 29120 25882
rect 29154 25880 29210 25882
rect 29244 25880 29300 25882
rect 29334 25880 29411 25882
rect 28449 25861 29411 25880
rect 28449 25857 28521 25861
rect 28449 25823 28468 25857
rect 28502 25823 28521 25857
rect 28449 25767 28521 25823
rect 29339 25838 29411 25861
rect 29339 25804 29358 25838
rect 29392 25804 29411 25838
rect 28449 25733 28468 25767
rect 28502 25733 28521 25767
rect 28449 25677 28521 25733
rect 28449 25643 28468 25677
rect 28502 25643 28521 25677
rect 28449 25587 28521 25643
rect 28449 25553 28468 25587
rect 28502 25553 28521 25587
rect 28449 25497 28521 25553
rect 28449 25463 28468 25497
rect 28502 25463 28521 25497
rect 28449 25407 28521 25463
rect 28449 25373 28468 25407
rect 28502 25373 28521 25407
rect 28449 25317 28521 25373
rect 28449 25283 28468 25317
rect 28502 25283 28521 25317
rect 28449 25227 28521 25283
rect 28449 25193 28468 25227
rect 28502 25193 28521 25227
rect 28449 25137 28521 25193
rect 28449 25103 28468 25137
rect 28502 25103 28521 25137
rect 28583 25740 29277 25799
rect 28583 25706 28644 25740
rect 28678 25712 28734 25740
rect 28768 25712 28824 25740
rect 28858 25712 28914 25740
rect 28690 25706 28734 25712
rect 28790 25706 28824 25712
rect 28890 25706 28914 25712
rect 28948 25712 29004 25740
rect 28948 25706 28956 25712
rect 28583 25678 28656 25706
rect 28690 25678 28756 25706
rect 28790 25678 28856 25706
rect 28890 25678 28956 25706
rect 28990 25706 29004 25712
rect 29038 25712 29094 25740
rect 29038 25706 29056 25712
rect 28990 25678 29056 25706
rect 29090 25706 29094 25712
rect 29128 25712 29184 25740
rect 29128 25706 29156 25712
rect 29218 25706 29277 25740
rect 29090 25678 29156 25706
rect 29190 25678 29277 25706
rect 28583 25650 29277 25678
rect 28583 25616 28644 25650
rect 28678 25616 28734 25650
rect 28768 25616 28824 25650
rect 28858 25616 28914 25650
rect 28948 25616 29004 25650
rect 29038 25616 29094 25650
rect 29128 25616 29184 25650
rect 29218 25616 29277 25650
rect 28583 25612 29277 25616
rect 28583 25578 28656 25612
rect 28690 25578 28756 25612
rect 28790 25578 28856 25612
rect 28890 25578 28956 25612
rect 28990 25578 29056 25612
rect 29090 25578 29156 25612
rect 29190 25578 29277 25612
rect 28583 25560 29277 25578
rect 28583 25526 28644 25560
rect 28678 25526 28734 25560
rect 28768 25526 28824 25560
rect 28858 25526 28914 25560
rect 28948 25526 29004 25560
rect 29038 25526 29094 25560
rect 29128 25526 29184 25560
rect 29218 25526 29277 25560
rect 28583 25512 29277 25526
rect 28583 25478 28656 25512
rect 28690 25478 28756 25512
rect 28790 25478 28856 25512
rect 28890 25478 28956 25512
rect 28990 25478 29056 25512
rect 29090 25478 29156 25512
rect 29190 25478 29277 25512
rect 28583 25470 29277 25478
rect 28583 25436 28644 25470
rect 28678 25436 28734 25470
rect 28768 25436 28824 25470
rect 28858 25436 28914 25470
rect 28948 25436 29004 25470
rect 29038 25436 29094 25470
rect 29128 25436 29184 25470
rect 29218 25436 29277 25470
rect 28583 25412 29277 25436
rect 28583 25380 28656 25412
rect 28690 25380 28756 25412
rect 28790 25380 28856 25412
rect 28890 25380 28956 25412
rect 28583 25346 28644 25380
rect 28690 25378 28734 25380
rect 28790 25378 28824 25380
rect 28890 25378 28914 25380
rect 28678 25346 28734 25378
rect 28768 25346 28824 25378
rect 28858 25346 28914 25378
rect 28948 25378 28956 25380
rect 28990 25380 29056 25412
rect 28990 25378 29004 25380
rect 28948 25346 29004 25378
rect 29038 25378 29056 25380
rect 29090 25380 29156 25412
rect 29190 25380 29277 25412
rect 29090 25378 29094 25380
rect 29038 25346 29094 25378
rect 29128 25378 29156 25380
rect 29128 25346 29184 25378
rect 29218 25346 29277 25380
rect 28583 25312 29277 25346
rect 28583 25290 28656 25312
rect 28690 25290 28756 25312
rect 28790 25290 28856 25312
rect 28890 25290 28956 25312
rect 28583 25256 28644 25290
rect 28690 25278 28734 25290
rect 28790 25278 28824 25290
rect 28890 25278 28914 25290
rect 28678 25256 28734 25278
rect 28768 25256 28824 25278
rect 28858 25256 28914 25278
rect 28948 25278 28956 25290
rect 28990 25290 29056 25312
rect 28990 25278 29004 25290
rect 28948 25256 29004 25278
rect 29038 25278 29056 25290
rect 29090 25290 29156 25312
rect 29190 25290 29277 25312
rect 29090 25278 29094 25290
rect 29038 25256 29094 25278
rect 29128 25278 29156 25290
rect 29128 25256 29184 25278
rect 29218 25256 29277 25290
rect 28583 25212 29277 25256
rect 28583 25200 28656 25212
rect 28690 25200 28756 25212
rect 28790 25200 28856 25212
rect 28890 25200 28956 25212
rect 28583 25166 28644 25200
rect 28690 25178 28734 25200
rect 28790 25178 28824 25200
rect 28890 25178 28914 25200
rect 28678 25166 28734 25178
rect 28768 25166 28824 25178
rect 28858 25166 28914 25178
rect 28948 25178 28956 25200
rect 28990 25200 29056 25212
rect 28990 25178 29004 25200
rect 28948 25166 29004 25178
rect 29038 25178 29056 25200
rect 29090 25200 29156 25212
rect 29190 25200 29277 25212
rect 29090 25178 29094 25200
rect 29038 25166 29094 25178
rect 29128 25178 29156 25200
rect 29128 25166 29184 25178
rect 29218 25166 29277 25200
rect 28583 25105 29277 25166
rect 29339 25748 29411 25804
rect 29339 25714 29358 25748
rect 29392 25714 29411 25748
rect 29339 25658 29411 25714
rect 29339 25624 29358 25658
rect 29392 25624 29411 25658
rect 29339 25568 29411 25624
rect 29339 25534 29358 25568
rect 29392 25534 29411 25568
rect 29339 25478 29411 25534
rect 29339 25444 29358 25478
rect 29392 25444 29411 25478
rect 29339 25388 29411 25444
rect 29339 25354 29358 25388
rect 29392 25354 29411 25388
rect 29339 25298 29411 25354
rect 29339 25264 29358 25298
rect 29392 25264 29411 25298
rect 29339 25208 29411 25264
rect 29339 25174 29358 25208
rect 29392 25174 29411 25208
rect 29339 25118 29411 25174
rect 28449 25043 28521 25103
rect 29339 25084 29358 25118
rect 29392 25084 29411 25118
rect 29339 25043 29411 25084
rect 28449 25024 29411 25043
rect 28449 24990 28546 25024
rect 28580 24990 28636 25024
rect 28670 24990 28726 25024
rect 28760 24990 28816 25024
rect 28850 24990 28906 25024
rect 28940 24990 28996 25024
rect 29030 24990 29086 25024
rect 29120 24990 29176 25024
rect 29210 24990 29266 25024
rect 29300 24990 29411 25024
rect 28449 24971 29411 24990
rect 29475 25914 29507 25948
rect 29541 25914 29660 25948
rect 29694 25914 29725 25948
rect 30815 25948 31065 25997
rect 29475 25858 29725 25914
rect 29475 25824 29507 25858
rect 29541 25824 29660 25858
rect 29694 25824 29725 25858
rect 29475 25768 29725 25824
rect 29475 25734 29507 25768
rect 29541 25734 29660 25768
rect 29694 25734 29725 25768
rect 29475 25678 29725 25734
rect 29475 25644 29507 25678
rect 29541 25644 29660 25678
rect 29694 25644 29725 25678
rect 29475 25588 29725 25644
rect 29475 25554 29507 25588
rect 29541 25554 29660 25588
rect 29694 25554 29725 25588
rect 29475 25498 29725 25554
rect 29475 25464 29507 25498
rect 29541 25464 29660 25498
rect 29694 25464 29725 25498
rect 29475 25408 29725 25464
rect 29475 25374 29507 25408
rect 29541 25374 29660 25408
rect 29694 25374 29725 25408
rect 29475 25318 29725 25374
rect 29475 25284 29507 25318
rect 29541 25284 29660 25318
rect 29694 25284 29725 25318
rect 29475 25228 29725 25284
rect 29475 25194 29507 25228
rect 29541 25194 29660 25228
rect 29694 25194 29725 25228
rect 29475 25138 29725 25194
rect 29475 25104 29507 25138
rect 29541 25104 29660 25138
rect 29694 25104 29725 25138
rect 29475 25048 29725 25104
rect 29475 25014 29507 25048
rect 29541 25014 29660 25048
rect 29694 25014 29725 25048
rect 28286 24924 28320 24958
rect 28354 24924 28385 24958
rect 28286 24907 28385 24924
rect 29475 24958 29725 25014
rect 29789 25916 30751 25933
rect 29789 25882 29810 25916
rect 29844 25882 29900 25916
rect 29934 25914 29990 25916
rect 30024 25914 30080 25916
rect 30114 25914 30170 25916
rect 30204 25914 30260 25916
rect 30294 25914 30350 25916
rect 30384 25914 30440 25916
rect 30474 25914 30530 25916
rect 30564 25914 30620 25916
rect 30654 25914 30710 25916
rect 29954 25882 29990 25914
rect 30044 25882 30080 25914
rect 30134 25882 30170 25914
rect 30224 25882 30260 25914
rect 30314 25882 30350 25914
rect 30404 25882 30440 25914
rect 30494 25882 30530 25914
rect 30584 25882 30620 25914
rect 30674 25882 30710 25914
rect 30744 25882 30751 25916
rect 29789 25880 29920 25882
rect 29954 25880 30010 25882
rect 30044 25880 30100 25882
rect 30134 25880 30190 25882
rect 30224 25880 30280 25882
rect 30314 25880 30370 25882
rect 30404 25880 30460 25882
rect 30494 25880 30550 25882
rect 30584 25880 30640 25882
rect 30674 25880 30751 25882
rect 29789 25861 30751 25880
rect 29789 25857 29861 25861
rect 29789 25823 29808 25857
rect 29842 25823 29861 25857
rect 29789 25767 29861 25823
rect 30679 25838 30751 25861
rect 30679 25804 30698 25838
rect 30732 25804 30751 25838
rect 29789 25733 29808 25767
rect 29842 25733 29861 25767
rect 29789 25677 29861 25733
rect 29789 25643 29808 25677
rect 29842 25643 29861 25677
rect 29789 25587 29861 25643
rect 29789 25553 29808 25587
rect 29842 25553 29861 25587
rect 29789 25497 29861 25553
rect 29789 25463 29808 25497
rect 29842 25463 29861 25497
rect 29789 25407 29861 25463
rect 29789 25373 29808 25407
rect 29842 25373 29861 25407
rect 29789 25317 29861 25373
rect 29789 25283 29808 25317
rect 29842 25283 29861 25317
rect 29789 25227 29861 25283
rect 29789 25193 29808 25227
rect 29842 25193 29861 25227
rect 29789 25137 29861 25193
rect 29789 25103 29808 25137
rect 29842 25103 29861 25137
rect 29923 25740 30617 25799
rect 29923 25706 29984 25740
rect 30018 25712 30074 25740
rect 30108 25712 30164 25740
rect 30198 25712 30254 25740
rect 30030 25706 30074 25712
rect 30130 25706 30164 25712
rect 30230 25706 30254 25712
rect 30288 25712 30344 25740
rect 30288 25706 30296 25712
rect 29923 25678 29996 25706
rect 30030 25678 30096 25706
rect 30130 25678 30196 25706
rect 30230 25678 30296 25706
rect 30330 25706 30344 25712
rect 30378 25712 30434 25740
rect 30378 25706 30396 25712
rect 30330 25678 30396 25706
rect 30430 25706 30434 25712
rect 30468 25712 30524 25740
rect 30468 25706 30496 25712
rect 30558 25706 30617 25740
rect 30430 25678 30496 25706
rect 30530 25678 30617 25706
rect 29923 25650 30617 25678
rect 29923 25616 29984 25650
rect 30018 25616 30074 25650
rect 30108 25616 30164 25650
rect 30198 25616 30254 25650
rect 30288 25616 30344 25650
rect 30378 25616 30434 25650
rect 30468 25616 30524 25650
rect 30558 25616 30617 25650
rect 29923 25612 30617 25616
rect 29923 25578 29996 25612
rect 30030 25578 30096 25612
rect 30130 25578 30196 25612
rect 30230 25578 30296 25612
rect 30330 25578 30396 25612
rect 30430 25578 30496 25612
rect 30530 25578 30617 25612
rect 29923 25560 30617 25578
rect 29923 25526 29984 25560
rect 30018 25526 30074 25560
rect 30108 25526 30164 25560
rect 30198 25526 30254 25560
rect 30288 25526 30344 25560
rect 30378 25526 30434 25560
rect 30468 25526 30524 25560
rect 30558 25526 30617 25560
rect 29923 25512 30617 25526
rect 29923 25478 29996 25512
rect 30030 25478 30096 25512
rect 30130 25478 30196 25512
rect 30230 25478 30296 25512
rect 30330 25478 30396 25512
rect 30430 25478 30496 25512
rect 30530 25478 30617 25512
rect 29923 25470 30617 25478
rect 29923 25436 29984 25470
rect 30018 25436 30074 25470
rect 30108 25436 30164 25470
rect 30198 25436 30254 25470
rect 30288 25436 30344 25470
rect 30378 25436 30434 25470
rect 30468 25436 30524 25470
rect 30558 25436 30617 25470
rect 29923 25412 30617 25436
rect 29923 25380 29996 25412
rect 30030 25380 30096 25412
rect 30130 25380 30196 25412
rect 30230 25380 30296 25412
rect 29923 25346 29984 25380
rect 30030 25378 30074 25380
rect 30130 25378 30164 25380
rect 30230 25378 30254 25380
rect 30018 25346 30074 25378
rect 30108 25346 30164 25378
rect 30198 25346 30254 25378
rect 30288 25378 30296 25380
rect 30330 25380 30396 25412
rect 30330 25378 30344 25380
rect 30288 25346 30344 25378
rect 30378 25378 30396 25380
rect 30430 25380 30496 25412
rect 30530 25380 30617 25412
rect 30430 25378 30434 25380
rect 30378 25346 30434 25378
rect 30468 25378 30496 25380
rect 30468 25346 30524 25378
rect 30558 25346 30617 25380
rect 29923 25312 30617 25346
rect 29923 25290 29996 25312
rect 30030 25290 30096 25312
rect 30130 25290 30196 25312
rect 30230 25290 30296 25312
rect 29923 25256 29984 25290
rect 30030 25278 30074 25290
rect 30130 25278 30164 25290
rect 30230 25278 30254 25290
rect 30018 25256 30074 25278
rect 30108 25256 30164 25278
rect 30198 25256 30254 25278
rect 30288 25278 30296 25290
rect 30330 25290 30396 25312
rect 30330 25278 30344 25290
rect 30288 25256 30344 25278
rect 30378 25278 30396 25290
rect 30430 25290 30496 25312
rect 30530 25290 30617 25312
rect 30430 25278 30434 25290
rect 30378 25256 30434 25278
rect 30468 25278 30496 25290
rect 30468 25256 30524 25278
rect 30558 25256 30617 25290
rect 29923 25212 30617 25256
rect 29923 25200 29996 25212
rect 30030 25200 30096 25212
rect 30130 25200 30196 25212
rect 30230 25200 30296 25212
rect 29923 25166 29984 25200
rect 30030 25178 30074 25200
rect 30130 25178 30164 25200
rect 30230 25178 30254 25200
rect 30018 25166 30074 25178
rect 30108 25166 30164 25178
rect 30198 25166 30254 25178
rect 30288 25178 30296 25200
rect 30330 25200 30396 25212
rect 30330 25178 30344 25200
rect 30288 25166 30344 25178
rect 30378 25178 30396 25200
rect 30430 25200 30496 25212
rect 30530 25200 30617 25212
rect 30430 25178 30434 25200
rect 30378 25166 30434 25178
rect 30468 25178 30496 25200
rect 30468 25166 30524 25178
rect 30558 25166 30617 25200
rect 29923 25105 30617 25166
rect 30679 25748 30751 25804
rect 30679 25714 30698 25748
rect 30732 25714 30751 25748
rect 30679 25658 30751 25714
rect 30679 25624 30698 25658
rect 30732 25624 30751 25658
rect 30679 25568 30751 25624
rect 30679 25534 30698 25568
rect 30732 25534 30751 25568
rect 30679 25478 30751 25534
rect 30679 25444 30698 25478
rect 30732 25444 30751 25478
rect 30679 25388 30751 25444
rect 30679 25354 30698 25388
rect 30732 25354 30751 25388
rect 30679 25298 30751 25354
rect 30679 25264 30698 25298
rect 30732 25264 30751 25298
rect 30679 25208 30751 25264
rect 30679 25174 30698 25208
rect 30732 25174 30751 25208
rect 30679 25118 30751 25174
rect 29789 25043 29861 25103
rect 30679 25084 30698 25118
rect 30732 25084 30751 25118
rect 30679 25043 30751 25084
rect 29789 25024 30751 25043
rect 29789 24990 29886 25024
rect 29920 24990 29976 25024
rect 30010 24990 30066 25024
rect 30100 24990 30156 25024
rect 30190 24990 30246 25024
rect 30280 24990 30336 25024
rect 30370 24990 30426 25024
rect 30460 24990 30516 25024
rect 30550 24990 30606 25024
rect 30640 24990 30751 25024
rect 29789 24971 30751 24990
rect 30815 25914 30847 25948
rect 30881 25914 31000 25948
rect 31034 25914 31065 25948
rect 32155 25948 32405 25997
rect 30815 25858 31065 25914
rect 30815 25824 30847 25858
rect 30881 25824 31000 25858
rect 31034 25824 31065 25858
rect 30815 25768 31065 25824
rect 30815 25734 30847 25768
rect 30881 25734 31000 25768
rect 31034 25734 31065 25768
rect 30815 25678 31065 25734
rect 30815 25644 30847 25678
rect 30881 25644 31000 25678
rect 31034 25644 31065 25678
rect 30815 25588 31065 25644
rect 30815 25554 30847 25588
rect 30881 25554 31000 25588
rect 31034 25554 31065 25588
rect 30815 25498 31065 25554
rect 30815 25464 30847 25498
rect 30881 25464 31000 25498
rect 31034 25464 31065 25498
rect 30815 25408 31065 25464
rect 30815 25374 30847 25408
rect 30881 25374 31000 25408
rect 31034 25374 31065 25408
rect 30815 25318 31065 25374
rect 30815 25284 30847 25318
rect 30881 25284 31000 25318
rect 31034 25284 31065 25318
rect 30815 25228 31065 25284
rect 30815 25194 30847 25228
rect 30881 25194 31000 25228
rect 31034 25194 31065 25228
rect 30815 25138 31065 25194
rect 30815 25104 30847 25138
rect 30881 25104 31000 25138
rect 31034 25104 31065 25138
rect 30815 25048 31065 25104
rect 30815 25014 30847 25048
rect 30881 25014 31000 25048
rect 31034 25014 31065 25048
rect 29475 24924 29507 24958
rect 29541 24924 29660 24958
rect 29694 24924 29725 24958
rect 29475 24907 29725 24924
rect 30815 24958 31065 25014
rect 31129 25916 32091 25933
rect 31129 25882 31150 25916
rect 31184 25882 31240 25916
rect 31274 25914 31330 25916
rect 31364 25914 31420 25916
rect 31454 25914 31510 25916
rect 31544 25914 31600 25916
rect 31634 25914 31690 25916
rect 31724 25914 31780 25916
rect 31814 25914 31870 25916
rect 31904 25914 31960 25916
rect 31994 25914 32050 25916
rect 31294 25882 31330 25914
rect 31384 25882 31420 25914
rect 31474 25882 31510 25914
rect 31564 25882 31600 25914
rect 31654 25882 31690 25914
rect 31744 25882 31780 25914
rect 31834 25882 31870 25914
rect 31924 25882 31960 25914
rect 32014 25882 32050 25914
rect 32084 25882 32091 25916
rect 31129 25880 31260 25882
rect 31294 25880 31350 25882
rect 31384 25880 31440 25882
rect 31474 25880 31530 25882
rect 31564 25880 31620 25882
rect 31654 25880 31710 25882
rect 31744 25880 31800 25882
rect 31834 25880 31890 25882
rect 31924 25880 31980 25882
rect 32014 25880 32091 25882
rect 31129 25861 32091 25880
rect 31129 25857 31201 25861
rect 31129 25823 31148 25857
rect 31182 25823 31201 25857
rect 31129 25767 31201 25823
rect 32019 25838 32091 25861
rect 32019 25804 32038 25838
rect 32072 25804 32091 25838
rect 31129 25733 31148 25767
rect 31182 25733 31201 25767
rect 31129 25677 31201 25733
rect 31129 25643 31148 25677
rect 31182 25643 31201 25677
rect 31129 25587 31201 25643
rect 31129 25553 31148 25587
rect 31182 25553 31201 25587
rect 31129 25497 31201 25553
rect 31129 25463 31148 25497
rect 31182 25463 31201 25497
rect 31129 25407 31201 25463
rect 31129 25373 31148 25407
rect 31182 25373 31201 25407
rect 31129 25317 31201 25373
rect 31129 25283 31148 25317
rect 31182 25283 31201 25317
rect 31129 25227 31201 25283
rect 31129 25193 31148 25227
rect 31182 25193 31201 25227
rect 31129 25137 31201 25193
rect 31129 25103 31148 25137
rect 31182 25103 31201 25137
rect 31263 25740 31957 25799
rect 31263 25706 31324 25740
rect 31358 25712 31414 25740
rect 31448 25712 31504 25740
rect 31538 25712 31594 25740
rect 31370 25706 31414 25712
rect 31470 25706 31504 25712
rect 31570 25706 31594 25712
rect 31628 25712 31684 25740
rect 31628 25706 31636 25712
rect 31263 25678 31336 25706
rect 31370 25678 31436 25706
rect 31470 25678 31536 25706
rect 31570 25678 31636 25706
rect 31670 25706 31684 25712
rect 31718 25712 31774 25740
rect 31718 25706 31736 25712
rect 31670 25678 31736 25706
rect 31770 25706 31774 25712
rect 31808 25712 31864 25740
rect 31808 25706 31836 25712
rect 31898 25706 31957 25740
rect 31770 25678 31836 25706
rect 31870 25678 31957 25706
rect 31263 25650 31957 25678
rect 31263 25616 31324 25650
rect 31358 25616 31414 25650
rect 31448 25616 31504 25650
rect 31538 25616 31594 25650
rect 31628 25616 31684 25650
rect 31718 25616 31774 25650
rect 31808 25616 31864 25650
rect 31898 25616 31957 25650
rect 31263 25612 31957 25616
rect 31263 25578 31336 25612
rect 31370 25578 31436 25612
rect 31470 25578 31536 25612
rect 31570 25578 31636 25612
rect 31670 25578 31736 25612
rect 31770 25578 31836 25612
rect 31870 25578 31957 25612
rect 31263 25560 31957 25578
rect 31263 25526 31324 25560
rect 31358 25526 31414 25560
rect 31448 25526 31504 25560
rect 31538 25526 31594 25560
rect 31628 25526 31684 25560
rect 31718 25526 31774 25560
rect 31808 25526 31864 25560
rect 31898 25526 31957 25560
rect 31263 25512 31957 25526
rect 31263 25478 31336 25512
rect 31370 25478 31436 25512
rect 31470 25478 31536 25512
rect 31570 25478 31636 25512
rect 31670 25478 31736 25512
rect 31770 25478 31836 25512
rect 31870 25478 31957 25512
rect 31263 25470 31957 25478
rect 31263 25436 31324 25470
rect 31358 25436 31414 25470
rect 31448 25436 31504 25470
rect 31538 25436 31594 25470
rect 31628 25436 31684 25470
rect 31718 25436 31774 25470
rect 31808 25436 31864 25470
rect 31898 25436 31957 25470
rect 31263 25412 31957 25436
rect 31263 25380 31336 25412
rect 31370 25380 31436 25412
rect 31470 25380 31536 25412
rect 31570 25380 31636 25412
rect 31263 25346 31324 25380
rect 31370 25378 31414 25380
rect 31470 25378 31504 25380
rect 31570 25378 31594 25380
rect 31358 25346 31414 25378
rect 31448 25346 31504 25378
rect 31538 25346 31594 25378
rect 31628 25378 31636 25380
rect 31670 25380 31736 25412
rect 31670 25378 31684 25380
rect 31628 25346 31684 25378
rect 31718 25378 31736 25380
rect 31770 25380 31836 25412
rect 31870 25380 31957 25412
rect 31770 25378 31774 25380
rect 31718 25346 31774 25378
rect 31808 25378 31836 25380
rect 31808 25346 31864 25378
rect 31898 25346 31957 25380
rect 31263 25312 31957 25346
rect 31263 25290 31336 25312
rect 31370 25290 31436 25312
rect 31470 25290 31536 25312
rect 31570 25290 31636 25312
rect 31263 25256 31324 25290
rect 31370 25278 31414 25290
rect 31470 25278 31504 25290
rect 31570 25278 31594 25290
rect 31358 25256 31414 25278
rect 31448 25256 31504 25278
rect 31538 25256 31594 25278
rect 31628 25278 31636 25290
rect 31670 25290 31736 25312
rect 31670 25278 31684 25290
rect 31628 25256 31684 25278
rect 31718 25278 31736 25290
rect 31770 25290 31836 25312
rect 31870 25290 31957 25312
rect 31770 25278 31774 25290
rect 31718 25256 31774 25278
rect 31808 25278 31836 25290
rect 31808 25256 31864 25278
rect 31898 25256 31957 25290
rect 31263 25212 31957 25256
rect 31263 25200 31336 25212
rect 31370 25200 31436 25212
rect 31470 25200 31536 25212
rect 31570 25200 31636 25212
rect 31263 25166 31324 25200
rect 31370 25178 31414 25200
rect 31470 25178 31504 25200
rect 31570 25178 31594 25200
rect 31358 25166 31414 25178
rect 31448 25166 31504 25178
rect 31538 25166 31594 25178
rect 31628 25178 31636 25200
rect 31670 25200 31736 25212
rect 31670 25178 31684 25200
rect 31628 25166 31684 25178
rect 31718 25178 31736 25200
rect 31770 25200 31836 25212
rect 31870 25200 31957 25212
rect 31770 25178 31774 25200
rect 31718 25166 31774 25178
rect 31808 25178 31836 25200
rect 31808 25166 31864 25178
rect 31898 25166 31957 25200
rect 31263 25105 31957 25166
rect 32019 25748 32091 25804
rect 32019 25714 32038 25748
rect 32072 25714 32091 25748
rect 32019 25658 32091 25714
rect 32019 25624 32038 25658
rect 32072 25624 32091 25658
rect 32019 25568 32091 25624
rect 32019 25534 32038 25568
rect 32072 25534 32091 25568
rect 32019 25478 32091 25534
rect 32019 25444 32038 25478
rect 32072 25444 32091 25478
rect 32019 25388 32091 25444
rect 32019 25354 32038 25388
rect 32072 25354 32091 25388
rect 32019 25298 32091 25354
rect 32019 25264 32038 25298
rect 32072 25264 32091 25298
rect 32019 25208 32091 25264
rect 32019 25174 32038 25208
rect 32072 25174 32091 25208
rect 32019 25118 32091 25174
rect 31129 25043 31201 25103
rect 32019 25084 32038 25118
rect 32072 25084 32091 25118
rect 32019 25043 32091 25084
rect 31129 25024 32091 25043
rect 31129 24990 31226 25024
rect 31260 24990 31316 25024
rect 31350 24990 31406 25024
rect 31440 24990 31496 25024
rect 31530 24990 31586 25024
rect 31620 24990 31676 25024
rect 31710 24990 31766 25024
rect 31800 24990 31856 25024
rect 31890 24990 31946 25024
rect 31980 24990 32091 25024
rect 31129 24971 32091 24990
rect 32155 25914 32187 25948
rect 32221 25914 32340 25948
rect 32374 25914 32405 25948
rect 33495 25948 33745 25997
rect 32155 25858 32405 25914
rect 32155 25824 32187 25858
rect 32221 25824 32340 25858
rect 32374 25824 32405 25858
rect 32155 25768 32405 25824
rect 32155 25734 32187 25768
rect 32221 25734 32340 25768
rect 32374 25734 32405 25768
rect 32155 25678 32405 25734
rect 32155 25644 32187 25678
rect 32221 25644 32340 25678
rect 32374 25644 32405 25678
rect 32155 25588 32405 25644
rect 32155 25554 32187 25588
rect 32221 25554 32340 25588
rect 32374 25554 32405 25588
rect 32155 25498 32405 25554
rect 32155 25464 32187 25498
rect 32221 25464 32340 25498
rect 32374 25464 32405 25498
rect 32155 25408 32405 25464
rect 32155 25374 32187 25408
rect 32221 25374 32340 25408
rect 32374 25374 32405 25408
rect 32155 25318 32405 25374
rect 32155 25284 32187 25318
rect 32221 25284 32340 25318
rect 32374 25284 32405 25318
rect 32155 25228 32405 25284
rect 32155 25194 32187 25228
rect 32221 25194 32340 25228
rect 32374 25194 32405 25228
rect 32155 25138 32405 25194
rect 32155 25104 32187 25138
rect 32221 25104 32340 25138
rect 32374 25104 32405 25138
rect 32155 25048 32405 25104
rect 32155 25014 32187 25048
rect 32221 25014 32340 25048
rect 32374 25014 32405 25048
rect 30815 24924 30847 24958
rect 30881 24924 31000 24958
rect 31034 24924 31065 24958
rect 30815 24907 31065 24924
rect 32155 24958 32405 25014
rect 32469 25916 33431 25933
rect 32469 25882 32490 25916
rect 32524 25882 32580 25916
rect 32614 25914 32670 25916
rect 32704 25914 32760 25916
rect 32794 25914 32850 25916
rect 32884 25914 32940 25916
rect 32974 25914 33030 25916
rect 33064 25914 33120 25916
rect 33154 25914 33210 25916
rect 33244 25914 33300 25916
rect 33334 25914 33390 25916
rect 32634 25882 32670 25914
rect 32724 25882 32760 25914
rect 32814 25882 32850 25914
rect 32904 25882 32940 25914
rect 32994 25882 33030 25914
rect 33084 25882 33120 25914
rect 33174 25882 33210 25914
rect 33264 25882 33300 25914
rect 33354 25882 33390 25914
rect 33424 25882 33431 25916
rect 32469 25880 32600 25882
rect 32634 25880 32690 25882
rect 32724 25880 32780 25882
rect 32814 25880 32870 25882
rect 32904 25880 32960 25882
rect 32994 25880 33050 25882
rect 33084 25880 33140 25882
rect 33174 25880 33230 25882
rect 33264 25880 33320 25882
rect 33354 25880 33431 25882
rect 32469 25861 33431 25880
rect 32469 25857 32541 25861
rect 32469 25823 32488 25857
rect 32522 25823 32541 25857
rect 32469 25767 32541 25823
rect 33359 25838 33431 25861
rect 33359 25804 33378 25838
rect 33412 25804 33431 25838
rect 32469 25733 32488 25767
rect 32522 25733 32541 25767
rect 32469 25677 32541 25733
rect 32469 25643 32488 25677
rect 32522 25643 32541 25677
rect 32469 25587 32541 25643
rect 32469 25553 32488 25587
rect 32522 25553 32541 25587
rect 32469 25497 32541 25553
rect 32469 25463 32488 25497
rect 32522 25463 32541 25497
rect 32469 25407 32541 25463
rect 32469 25373 32488 25407
rect 32522 25373 32541 25407
rect 32469 25317 32541 25373
rect 32469 25283 32488 25317
rect 32522 25283 32541 25317
rect 32469 25227 32541 25283
rect 32469 25193 32488 25227
rect 32522 25193 32541 25227
rect 32469 25137 32541 25193
rect 32469 25103 32488 25137
rect 32522 25103 32541 25137
rect 32603 25740 33297 25799
rect 32603 25706 32664 25740
rect 32698 25712 32754 25740
rect 32788 25712 32844 25740
rect 32878 25712 32934 25740
rect 32710 25706 32754 25712
rect 32810 25706 32844 25712
rect 32910 25706 32934 25712
rect 32968 25712 33024 25740
rect 32968 25706 32976 25712
rect 32603 25678 32676 25706
rect 32710 25678 32776 25706
rect 32810 25678 32876 25706
rect 32910 25678 32976 25706
rect 33010 25706 33024 25712
rect 33058 25712 33114 25740
rect 33058 25706 33076 25712
rect 33010 25678 33076 25706
rect 33110 25706 33114 25712
rect 33148 25712 33204 25740
rect 33148 25706 33176 25712
rect 33238 25706 33297 25740
rect 33110 25678 33176 25706
rect 33210 25678 33297 25706
rect 32603 25650 33297 25678
rect 32603 25616 32664 25650
rect 32698 25616 32754 25650
rect 32788 25616 32844 25650
rect 32878 25616 32934 25650
rect 32968 25616 33024 25650
rect 33058 25616 33114 25650
rect 33148 25616 33204 25650
rect 33238 25616 33297 25650
rect 32603 25612 33297 25616
rect 32603 25578 32676 25612
rect 32710 25578 32776 25612
rect 32810 25578 32876 25612
rect 32910 25578 32976 25612
rect 33010 25578 33076 25612
rect 33110 25578 33176 25612
rect 33210 25578 33297 25612
rect 32603 25560 33297 25578
rect 32603 25526 32664 25560
rect 32698 25526 32754 25560
rect 32788 25526 32844 25560
rect 32878 25526 32934 25560
rect 32968 25526 33024 25560
rect 33058 25526 33114 25560
rect 33148 25526 33204 25560
rect 33238 25526 33297 25560
rect 32603 25512 33297 25526
rect 32603 25478 32676 25512
rect 32710 25478 32776 25512
rect 32810 25478 32876 25512
rect 32910 25478 32976 25512
rect 33010 25478 33076 25512
rect 33110 25478 33176 25512
rect 33210 25478 33297 25512
rect 32603 25470 33297 25478
rect 32603 25436 32664 25470
rect 32698 25436 32754 25470
rect 32788 25436 32844 25470
rect 32878 25436 32934 25470
rect 32968 25436 33024 25470
rect 33058 25436 33114 25470
rect 33148 25436 33204 25470
rect 33238 25436 33297 25470
rect 32603 25412 33297 25436
rect 32603 25380 32676 25412
rect 32710 25380 32776 25412
rect 32810 25380 32876 25412
rect 32910 25380 32976 25412
rect 32603 25346 32664 25380
rect 32710 25378 32754 25380
rect 32810 25378 32844 25380
rect 32910 25378 32934 25380
rect 32698 25346 32754 25378
rect 32788 25346 32844 25378
rect 32878 25346 32934 25378
rect 32968 25378 32976 25380
rect 33010 25380 33076 25412
rect 33010 25378 33024 25380
rect 32968 25346 33024 25378
rect 33058 25378 33076 25380
rect 33110 25380 33176 25412
rect 33210 25380 33297 25412
rect 33110 25378 33114 25380
rect 33058 25346 33114 25378
rect 33148 25378 33176 25380
rect 33148 25346 33204 25378
rect 33238 25346 33297 25380
rect 32603 25312 33297 25346
rect 32603 25290 32676 25312
rect 32710 25290 32776 25312
rect 32810 25290 32876 25312
rect 32910 25290 32976 25312
rect 32603 25256 32664 25290
rect 32710 25278 32754 25290
rect 32810 25278 32844 25290
rect 32910 25278 32934 25290
rect 32698 25256 32754 25278
rect 32788 25256 32844 25278
rect 32878 25256 32934 25278
rect 32968 25278 32976 25290
rect 33010 25290 33076 25312
rect 33010 25278 33024 25290
rect 32968 25256 33024 25278
rect 33058 25278 33076 25290
rect 33110 25290 33176 25312
rect 33210 25290 33297 25312
rect 33110 25278 33114 25290
rect 33058 25256 33114 25278
rect 33148 25278 33176 25290
rect 33148 25256 33204 25278
rect 33238 25256 33297 25290
rect 32603 25212 33297 25256
rect 32603 25200 32676 25212
rect 32710 25200 32776 25212
rect 32810 25200 32876 25212
rect 32910 25200 32976 25212
rect 32603 25166 32664 25200
rect 32710 25178 32754 25200
rect 32810 25178 32844 25200
rect 32910 25178 32934 25200
rect 32698 25166 32754 25178
rect 32788 25166 32844 25178
rect 32878 25166 32934 25178
rect 32968 25178 32976 25200
rect 33010 25200 33076 25212
rect 33010 25178 33024 25200
rect 32968 25166 33024 25178
rect 33058 25178 33076 25200
rect 33110 25200 33176 25212
rect 33210 25200 33297 25212
rect 33110 25178 33114 25200
rect 33058 25166 33114 25178
rect 33148 25178 33176 25200
rect 33148 25166 33204 25178
rect 33238 25166 33297 25200
rect 32603 25105 33297 25166
rect 33359 25748 33431 25804
rect 33359 25714 33378 25748
rect 33412 25714 33431 25748
rect 33359 25658 33431 25714
rect 33359 25624 33378 25658
rect 33412 25624 33431 25658
rect 33359 25568 33431 25624
rect 33359 25534 33378 25568
rect 33412 25534 33431 25568
rect 33359 25478 33431 25534
rect 33359 25444 33378 25478
rect 33412 25444 33431 25478
rect 33359 25388 33431 25444
rect 33359 25354 33378 25388
rect 33412 25354 33431 25388
rect 33359 25298 33431 25354
rect 33359 25264 33378 25298
rect 33412 25264 33431 25298
rect 33359 25208 33431 25264
rect 33359 25174 33378 25208
rect 33412 25174 33431 25208
rect 33359 25118 33431 25174
rect 32469 25043 32541 25103
rect 33359 25084 33378 25118
rect 33412 25084 33431 25118
rect 33359 25043 33431 25084
rect 32469 25024 33431 25043
rect 32469 24990 32566 25024
rect 32600 24990 32656 25024
rect 32690 24990 32746 25024
rect 32780 24990 32836 25024
rect 32870 24990 32926 25024
rect 32960 24990 33016 25024
rect 33050 24990 33106 25024
rect 33140 24990 33196 25024
rect 33230 24990 33286 25024
rect 33320 24990 33431 25024
rect 32469 24971 33431 24990
rect 33495 25914 33527 25948
rect 33561 25914 33680 25948
rect 33714 25914 33745 25948
rect 34835 25948 35085 25997
rect 33495 25858 33745 25914
rect 33495 25824 33527 25858
rect 33561 25824 33680 25858
rect 33714 25824 33745 25858
rect 33495 25768 33745 25824
rect 33495 25734 33527 25768
rect 33561 25734 33680 25768
rect 33714 25734 33745 25768
rect 33495 25678 33745 25734
rect 33495 25644 33527 25678
rect 33561 25644 33680 25678
rect 33714 25644 33745 25678
rect 33495 25588 33745 25644
rect 33495 25554 33527 25588
rect 33561 25554 33680 25588
rect 33714 25554 33745 25588
rect 33495 25498 33745 25554
rect 33495 25464 33527 25498
rect 33561 25464 33680 25498
rect 33714 25464 33745 25498
rect 33495 25408 33745 25464
rect 33495 25374 33527 25408
rect 33561 25374 33680 25408
rect 33714 25374 33745 25408
rect 33495 25318 33745 25374
rect 33495 25284 33527 25318
rect 33561 25284 33680 25318
rect 33714 25284 33745 25318
rect 33495 25228 33745 25284
rect 33495 25194 33527 25228
rect 33561 25194 33680 25228
rect 33714 25194 33745 25228
rect 33495 25138 33745 25194
rect 33495 25104 33527 25138
rect 33561 25104 33680 25138
rect 33714 25104 33745 25138
rect 33495 25048 33745 25104
rect 33495 25014 33527 25048
rect 33561 25014 33680 25048
rect 33714 25014 33745 25048
rect 32155 24924 32187 24958
rect 32221 24924 32340 24958
rect 32374 24924 32405 24958
rect 32155 24907 32405 24924
rect 33495 24958 33745 25014
rect 33809 25916 34771 25933
rect 33809 25882 33830 25916
rect 33864 25882 33920 25916
rect 33954 25914 34010 25916
rect 34044 25914 34100 25916
rect 34134 25914 34190 25916
rect 34224 25914 34280 25916
rect 34314 25914 34370 25916
rect 34404 25914 34460 25916
rect 34494 25914 34550 25916
rect 34584 25914 34640 25916
rect 34674 25914 34730 25916
rect 33974 25882 34010 25914
rect 34064 25882 34100 25914
rect 34154 25882 34190 25914
rect 34244 25882 34280 25914
rect 34334 25882 34370 25914
rect 34424 25882 34460 25914
rect 34514 25882 34550 25914
rect 34604 25882 34640 25914
rect 34694 25882 34730 25914
rect 34764 25882 34771 25916
rect 33809 25880 33940 25882
rect 33974 25880 34030 25882
rect 34064 25880 34120 25882
rect 34154 25880 34210 25882
rect 34244 25880 34300 25882
rect 34334 25880 34390 25882
rect 34424 25880 34480 25882
rect 34514 25880 34570 25882
rect 34604 25880 34660 25882
rect 34694 25880 34771 25882
rect 33809 25861 34771 25880
rect 33809 25857 33881 25861
rect 33809 25823 33828 25857
rect 33862 25823 33881 25857
rect 33809 25767 33881 25823
rect 34699 25838 34771 25861
rect 34699 25804 34718 25838
rect 34752 25804 34771 25838
rect 33809 25733 33828 25767
rect 33862 25733 33881 25767
rect 33809 25677 33881 25733
rect 33809 25643 33828 25677
rect 33862 25643 33881 25677
rect 33809 25587 33881 25643
rect 33809 25553 33828 25587
rect 33862 25553 33881 25587
rect 33809 25497 33881 25553
rect 33809 25463 33828 25497
rect 33862 25463 33881 25497
rect 33809 25407 33881 25463
rect 33809 25373 33828 25407
rect 33862 25373 33881 25407
rect 33809 25317 33881 25373
rect 33809 25283 33828 25317
rect 33862 25283 33881 25317
rect 33809 25227 33881 25283
rect 33809 25193 33828 25227
rect 33862 25193 33881 25227
rect 33809 25137 33881 25193
rect 33809 25103 33828 25137
rect 33862 25103 33881 25137
rect 33943 25740 34637 25799
rect 33943 25706 34004 25740
rect 34038 25712 34094 25740
rect 34128 25712 34184 25740
rect 34218 25712 34274 25740
rect 34050 25706 34094 25712
rect 34150 25706 34184 25712
rect 34250 25706 34274 25712
rect 34308 25712 34364 25740
rect 34308 25706 34316 25712
rect 33943 25678 34016 25706
rect 34050 25678 34116 25706
rect 34150 25678 34216 25706
rect 34250 25678 34316 25706
rect 34350 25706 34364 25712
rect 34398 25712 34454 25740
rect 34398 25706 34416 25712
rect 34350 25678 34416 25706
rect 34450 25706 34454 25712
rect 34488 25712 34544 25740
rect 34488 25706 34516 25712
rect 34578 25706 34637 25740
rect 34450 25678 34516 25706
rect 34550 25678 34637 25706
rect 33943 25650 34637 25678
rect 33943 25616 34004 25650
rect 34038 25616 34094 25650
rect 34128 25616 34184 25650
rect 34218 25616 34274 25650
rect 34308 25616 34364 25650
rect 34398 25616 34454 25650
rect 34488 25616 34544 25650
rect 34578 25616 34637 25650
rect 33943 25612 34637 25616
rect 33943 25578 34016 25612
rect 34050 25578 34116 25612
rect 34150 25578 34216 25612
rect 34250 25578 34316 25612
rect 34350 25578 34416 25612
rect 34450 25578 34516 25612
rect 34550 25578 34637 25612
rect 33943 25560 34637 25578
rect 33943 25526 34004 25560
rect 34038 25526 34094 25560
rect 34128 25526 34184 25560
rect 34218 25526 34274 25560
rect 34308 25526 34364 25560
rect 34398 25526 34454 25560
rect 34488 25526 34544 25560
rect 34578 25526 34637 25560
rect 33943 25512 34637 25526
rect 33943 25478 34016 25512
rect 34050 25478 34116 25512
rect 34150 25478 34216 25512
rect 34250 25478 34316 25512
rect 34350 25478 34416 25512
rect 34450 25478 34516 25512
rect 34550 25478 34637 25512
rect 33943 25470 34637 25478
rect 33943 25436 34004 25470
rect 34038 25436 34094 25470
rect 34128 25436 34184 25470
rect 34218 25436 34274 25470
rect 34308 25436 34364 25470
rect 34398 25436 34454 25470
rect 34488 25436 34544 25470
rect 34578 25436 34637 25470
rect 33943 25412 34637 25436
rect 33943 25380 34016 25412
rect 34050 25380 34116 25412
rect 34150 25380 34216 25412
rect 34250 25380 34316 25412
rect 33943 25346 34004 25380
rect 34050 25378 34094 25380
rect 34150 25378 34184 25380
rect 34250 25378 34274 25380
rect 34038 25346 34094 25378
rect 34128 25346 34184 25378
rect 34218 25346 34274 25378
rect 34308 25378 34316 25380
rect 34350 25380 34416 25412
rect 34350 25378 34364 25380
rect 34308 25346 34364 25378
rect 34398 25378 34416 25380
rect 34450 25380 34516 25412
rect 34550 25380 34637 25412
rect 34450 25378 34454 25380
rect 34398 25346 34454 25378
rect 34488 25378 34516 25380
rect 34488 25346 34544 25378
rect 34578 25346 34637 25380
rect 33943 25312 34637 25346
rect 33943 25290 34016 25312
rect 34050 25290 34116 25312
rect 34150 25290 34216 25312
rect 34250 25290 34316 25312
rect 33943 25256 34004 25290
rect 34050 25278 34094 25290
rect 34150 25278 34184 25290
rect 34250 25278 34274 25290
rect 34038 25256 34094 25278
rect 34128 25256 34184 25278
rect 34218 25256 34274 25278
rect 34308 25278 34316 25290
rect 34350 25290 34416 25312
rect 34350 25278 34364 25290
rect 34308 25256 34364 25278
rect 34398 25278 34416 25290
rect 34450 25290 34516 25312
rect 34550 25290 34637 25312
rect 34450 25278 34454 25290
rect 34398 25256 34454 25278
rect 34488 25278 34516 25290
rect 34488 25256 34544 25278
rect 34578 25256 34637 25290
rect 33943 25212 34637 25256
rect 33943 25200 34016 25212
rect 34050 25200 34116 25212
rect 34150 25200 34216 25212
rect 34250 25200 34316 25212
rect 33943 25166 34004 25200
rect 34050 25178 34094 25200
rect 34150 25178 34184 25200
rect 34250 25178 34274 25200
rect 34038 25166 34094 25178
rect 34128 25166 34184 25178
rect 34218 25166 34274 25178
rect 34308 25178 34316 25200
rect 34350 25200 34416 25212
rect 34350 25178 34364 25200
rect 34308 25166 34364 25178
rect 34398 25178 34416 25200
rect 34450 25200 34516 25212
rect 34550 25200 34637 25212
rect 34450 25178 34454 25200
rect 34398 25166 34454 25178
rect 34488 25178 34516 25200
rect 34488 25166 34544 25178
rect 34578 25166 34637 25200
rect 33943 25105 34637 25166
rect 34699 25748 34771 25804
rect 34699 25714 34718 25748
rect 34752 25714 34771 25748
rect 34699 25658 34771 25714
rect 34699 25624 34718 25658
rect 34752 25624 34771 25658
rect 34699 25568 34771 25624
rect 34699 25534 34718 25568
rect 34752 25534 34771 25568
rect 34699 25478 34771 25534
rect 34699 25444 34718 25478
rect 34752 25444 34771 25478
rect 34699 25388 34771 25444
rect 34699 25354 34718 25388
rect 34752 25354 34771 25388
rect 34699 25298 34771 25354
rect 34699 25264 34718 25298
rect 34752 25264 34771 25298
rect 34699 25208 34771 25264
rect 34699 25174 34718 25208
rect 34752 25174 34771 25208
rect 34699 25118 34771 25174
rect 33809 25043 33881 25103
rect 34699 25084 34718 25118
rect 34752 25084 34771 25118
rect 34699 25043 34771 25084
rect 33809 25024 34771 25043
rect 33809 24990 33906 25024
rect 33940 24990 33996 25024
rect 34030 24990 34086 25024
rect 34120 24990 34176 25024
rect 34210 24990 34266 25024
rect 34300 24990 34356 25024
rect 34390 24990 34446 25024
rect 34480 24990 34536 25024
rect 34570 24990 34626 25024
rect 34660 24990 34771 25024
rect 33809 24971 34771 24990
rect 34835 25914 34867 25948
rect 34901 25914 35020 25948
rect 35054 25914 35085 25948
rect 36175 25948 36425 25997
rect 34835 25858 35085 25914
rect 34835 25824 34867 25858
rect 34901 25824 35020 25858
rect 35054 25824 35085 25858
rect 34835 25768 35085 25824
rect 34835 25734 34867 25768
rect 34901 25734 35020 25768
rect 35054 25734 35085 25768
rect 34835 25678 35085 25734
rect 34835 25644 34867 25678
rect 34901 25644 35020 25678
rect 35054 25644 35085 25678
rect 34835 25588 35085 25644
rect 34835 25554 34867 25588
rect 34901 25554 35020 25588
rect 35054 25554 35085 25588
rect 34835 25498 35085 25554
rect 34835 25464 34867 25498
rect 34901 25464 35020 25498
rect 35054 25464 35085 25498
rect 34835 25408 35085 25464
rect 34835 25374 34867 25408
rect 34901 25374 35020 25408
rect 35054 25374 35085 25408
rect 34835 25318 35085 25374
rect 34835 25284 34867 25318
rect 34901 25284 35020 25318
rect 35054 25284 35085 25318
rect 34835 25228 35085 25284
rect 34835 25194 34867 25228
rect 34901 25194 35020 25228
rect 35054 25194 35085 25228
rect 34835 25138 35085 25194
rect 34835 25104 34867 25138
rect 34901 25104 35020 25138
rect 35054 25104 35085 25138
rect 34835 25048 35085 25104
rect 34835 25014 34867 25048
rect 34901 25014 35020 25048
rect 35054 25014 35085 25048
rect 33495 24924 33527 24958
rect 33561 24924 33680 24958
rect 33714 24924 33745 24958
rect 33495 24907 33745 24924
rect 34835 24958 35085 25014
rect 35149 25916 36111 25933
rect 35149 25882 35170 25916
rect 35204 25882 35260 25916
rect 35294 25914 35350 25916
rect 35384 25914 35440 25916
rect 35474 25914 35530 25916
rect 35564 25914 35620 25916
rect 35654 25914 35710 25916
rect 35744 25914 35800 25916
rect 35834 25914 35890 25916
rect 35924 25914 35980 25916
rect 36014 25914 36070 25916
rect 35314 25882 35350 25914
rect 35404 25882 35440 25914
rect 35494 25882 35530 25914
rect 35584 25882 35620 25914
rect 35674 25882 35710 25914
rect 35764 25882 35800 25914
rect 35854 25882 35890 25914
rect 35944 25882 35980 25914
rect 36034 25882 36070 25914
rect 36104 25882 36111 25916
rect 35149 25880 35280 25882
rect 35314 25880 35370 25882
rect 35404 25880 35460 25882
rect 35494 25880 35550 25882
rect 35584 25880 35640 25882
rect 35674 25880 35730 25882
rect 35764 25880 35820 25882
rect 35854 25880 35910 25882
rect 35944 25880 36000 25882
rect 36034 25880 36111 25882
rect 35149 25861 36111 25880
rect 35149 25857 35221 25861
rect 35149 25823 35168 25857
rect 35202 25823 35221 25857
rect 35149 25767 35221 25823
rect 36039 25838 36111 25861
rect 36039 25804 36058 25838
rect 36092 25804 36111 25838
rect 35149 25733 35168 25767
rect 35202 25733 35221 25767
rect 35149 25677 35221 25733
rect 35149 25643 35168 25677
rect 35202 25643 35221 25677
rect 35149 25587 35221 25643
rect 35149 25553 35168 25587
rect 35202 25553 35221 25587
rect 35149 25497 35221 25553
rect 35149 25463 35168 25497
rect 35202 25463 35221 25497
rect 35149 25407 35221 25463
rect 35149 25373 35168 25407
rect 35202 25373 35221 25407
rect 35149 25317 35221 25373
rect 35149 25283 35168 25317
rect 35202 25283 35221 25317
rect 35149 25227 35221 25283
rect 35149 25193 35168 25227
rect 35202 25193 35221 25227
rect 35149 25137 35221 25193
rect 35149 25103 35168 25137
rect 35202 25103 35221 25137
rect 35283 25740 35977 25799
rect 35283 25706 35344 25740
rect 35378 25712 35434 25740
rect 35468 25712 35524 25740
rect 35558 25712 35614 25740
rect 35390 25706 35434 25712
rect 35490 25706 35524 25712
rect 35590 25706 35614 25712
rect 35648 25712 35704 25740
rect 35648 25706 35656 25712
rect 35283 25678 35356 25706
rect 35390 25678 35456 25706
rect 35490 25678 35556 25706
rect 35590 25678 35656 25706
rect 35690 25706 35704 25712
rect 35738 25712 35794 25740
rect 35738 25706 35756 25712
rect 35690 25678 35756 25706
rect 35790 25706 35794 25712
rect 35828 25712 35884 25740
rect 35828 25706 35856 25712
rect 35918 25706 35977 25740
rect 35790 25678 35856 25706
rect 35890 25678 35977 25706
rect 35283 25650 35977 25678
rect 35283 25616 35344 25650
rect 35378 25616 35434 25650
rect 35468 25616 35524 25650
rect 35558 25616 35614 25650
rect 35648 25616 35704 25650
rect 35738 25616 35794 25650
rect 35828 25616 35884 25650
rect 35918 25616 35977 25650
rect 35283 25612 35977 25616
rect 35283 25578 35356 25612
rect 35390 25578 35456 25612
rect 35490 25578 35556 25612
rect 35590 25578 35656 25612
rect 35690 25578 35756 25612
rect 35790 25578 35856 25612
rect 35890 25578 35977 25612
rect 35283 25560 35977 25578
rect 35283 25526 35344 25560
rect 35378 25526 35434 25560
rect 35468 25526 35524 25560
rect 35558 25526 35614 25560
rect 35648 25526 35704 25560
rect 35738 25526 35794 25560
rect 35828 25526 35884 25560
rect 35918 25526 35977 25560
rect 35283 25512 35977 25526
rect 35283 25478 35356 25512
rect 35390 25478 35456 25512
rect 35490 25478 35556 25512
rect 35590 25478 35656 25512
rect 35690 25478 35756 25512
rect 35790 25478 35856 25512
rect 35890 25478 35977 25512
rect 35283 25470 35977 25478
rect 35283 25436 35344 25470
rect 35378 25436 35434 25470
rect 35468 25436 35524 25470
rect 35558 25436 35614 25470
rect 35648 25436 35704 25470
rect 35738 25436 35794 25470
rect 35828 25436 35884 25470
rect 35918 25436 35977 25470
rect 35283 25412 35977 25436
rect 35283 25380 35356 25412
rect 35390 25380 35456 25412
rect 35490 25380 35556 25412
rect 35590 25380 35656 25412
rect 35283 25346 35344 25380
rect 35390 25378 35434 25380
rect 35490 25378 35524 25380
rect 35590 25378 35614 25380
rect 35378 25346 35434 25378
rect 35468 25346 35524 25378
rect 35558 25346 35614 25378
rect 35648 25378 35656 25380
rect 35690 25380 35756 25412
rect 35690 25378 35704 25380
rect 35648 25346 35704 25378
rect 35738 25378 35756 25380
rect 35790 25380 35856 25412
rect 35890 25380 35977 25412
rect 35790 25378 35794 25380
rect 35738 25346 35794 25378
rect 35828 25378 35856 25380
rect 35828 25346 35884 25378
rect 35918 25346 35977 25380
rect 35283 25312 35977 25346
rect 35283 25290 35356 25312
rect 35390 25290 35456 25312
rect 35490 25290 35556 25312
rect 35590 25290 35656 25312
rect 35283 25256 35344 25290
rect 35390 25278 35434 25290
rect 35490 25278 35524 25290
rect 35590 25278 35614 25290
rect 35378 25256 35434 25278
rect 35468 25256 35524 25278
rect 35558 25256 35614 25278
rect 35648 25278 35656 25290
rect 35690 25290 35756 25312
rect 35690 25278 35704 25290
rect 35648 25256 35704 25278
rect 35738 25278 35756 25290
rect 35790 25290 35856 25312
rect 35890 25290 35977 25312
rect 35790 25278 35794 25290
rect 35738 25256 35794 25278
rect 35828 25278 35856 25290
rect 35828 25256 35884 25278
rect 35918 25256 35977 25290
rect 35283 25212 35977 25256
rect 35283 25200 35356 25212
rect 35390 25200 35456 25212
rect 35490 25200 35556 25212
rect 35590 25200 35656 25212
rect 35283 25166 35344 25200
rect 35390 25178 35434 25200
rect 35490 25178 35524 25200
rect 35590 25178 35614 25200
rect 35378 25166 35434 25178
rect 35468 25166 35524 25178
rect 35558 25166 35614 25178
rect 35648 25178 35656 25200
rect 35690 25200 35756 25212
rect 35690 25178 35704 25200
rect 35648 25166 35704 25178
rect 35738 25178 35756 25200
rect 35790 25200 35856 25212
rect 35890 25200 35977 25212
rect 35790 25178 35794 25200
rect 35738 25166 35794 25178
rect 35828 25178 35856 25200
rect 35828 25166 35884 25178
rect 35918 25166 35977 25200
rect 35283 25105 35977 25166
rect 36039 25748 36111 25804
rect 36039 25714 36058 25748
rect 36092 25714 36111 25748
rect 36039 25658 36111 25714
rect 36039 25624 36058 25658
rect 36092 25624 36111 25658
rect 36039 25568 36111 25624
rect 36039 25534 36058 25568
rect 36092 25534 36111 25568
rect 36039 25478 36111 25534
rect 36039 25444 36058 25478
rect 36092 25444 36111 25478
rect 36039 25388 36111 25444
rect 36039 25354 36058 25388
rect 36092 25354 36111 25388
rect 36039 25298 36111 25354
rect 36039 25264 36058 25298
rect 36092 25264 36111 25298
rect 36039 25208 36111 25264
rect 36039 25174 36058 25208
rect 36092 25174 36111 25208
rect 36039 25118 36111 25174
rect 35149 25043 35221 25103
rect 36039 25084 36058 25118
rect 36092 25084 36111 25118
rect 36039 25043 36111 25084
rect 35149 25024 36111 25043
rect 35149 24990 35246 25024
rect 35280 24990 35336 25024
rect 35370 24990 35426 25024
rect 35460 24990 35516 25024
rect 35550 24990 35606 25024
rect 35640 24990 35696 25024
rect 35730 24990 35786 25024
rect 35820 24990 35876 25024
rect 35910 24990 35966 25024
rect 36000 24990 36111 25024
rect 35149 24971 36111 24990
rect 36175 25914 36207 25948
rect 36241 25914 36360 25948
rect 36394 25914 36425 25948
rect 37515 25948 37765 25997
rect 36175 25858 36425 25914
rect 36175 25824 36207 25858
rect 36241 25824 36360 25858
rect 36394 25824 36425 25858
rect 36175 25768 36425 25824
rect 36175 25734 36207 25768
rect 36241 25734 36360 25768
rect 36394 25734 36425 25768
rect 36175 25678 36425 25734
rect 36175 25644 36207 25678
rect 36241 25644 36360 25678
rect 36394 25644 36425 25678
rect 36175 25588 36425 25644
rect 36175 25554 36207 25588
rect 36241 25554 36360 25588
rect 36394 25554 36425 25588
rect 36175 25498 36425 25554
rect 36175 25464 36207 25498
rect 36241 25464 36360 25498
rect 36394 25464 36425 25498
rect 36175 25408 36425 25464
rect 36175 25374 36207 25408
rect 36241 25374 36360 25408
rect 36394 25374 36425 25408
rect 36175 25318 36425 25374
rect 36175 25284 36207 25318
rect 36241 25284 36360 25318
rect 36394 25284 36425 25318
rect 36175 25228 36425 25284
rect 36175 25194 36207 25228
rect 36241 25194 36360 25228
rect 36394 25194 36425 25228
rect 36175 25138 36425 25194
rect 36175 25104 36207 25138
rect 36241 25104 36360 25138
rect 36394 25104 36425 25138
rect 36175 25048 36425 25104
rect 36175 25014 36207 25048
rect 36241 25014 36360 25048
rect 36394 25014 36425 25048
rect 34835 24924 34867 24958
rect 34901 24924 35020 24958
rect 35054 24924 35085 24958
rect 34835 24907 35085 24924
rect 36175 24958 36425 25014
rect 36489 25916 37451 25933
rect 36489 25882 36510 25916
rect 36544 25882 36600 25916
rect 36634 25914 36690 25916
rect 36724 25914 36780 25916
rect 36814 25914 36870 25916
rect 36904 25914 36960 25916
rect 36994 25914 37050 25916
rect 37084 25914 37140 25916
rect 37174 25914 37230 25916
rect 37264 25914 37320 25916
rect 37354 25914 37410 25916
rect 36654 25882 36690 25914
rect 36744 25882 36780 25914
rect 36834 25882 36870 25914
rect 36924 25882 36960 25914
rect 37014 25882 37050 25914
rect 37104 25882 37140 25914
rect 37194 25882 37230 25914
rect 37284 25882 37320 25914
rect 37374 25882 37410 25914
rect 37444 25882 37451 25916
rect 36489 25880 36620 25882
rect 36654 25880 36710 25882
rect 36744 25880 36800 25882
rect 36834 25880 36890 25882
rect 36924 25880 36980 25882
rect 37014 25880 37070 25882
rect 37104 25880 37160 25882
rect 37194 25880 37250 25882
rect 37284 25880 37340 25882
rect 37374 25880 37451 25882
rect 36489 25861 37451 25880
rect 36489 25857 36561 25861
rect 36489 25823 36508 25857
rect 36542 25823 36561 25857
rect 36489 25767 36561 25823
rect 37379 25838 37451 25861
rect 37379 25804 37398 25838
rect 37432 25804 37451 25838
rect 36489 25733 36508 25767
rect 36542 25733 36561 25767
rect 36489 25677 36561 25733
rect 36489 25643 36508 25677
rect 36542 25643 36561 25677
rect 36489 25587 36561 25643
rect 36489 25553 36508 25587
rect 36542 25553 36561 25587
rect 36489 25497 36561 25553
rect 36489 25463 36508 25497
rect 36542 25463 36561 25497
rect 36489 25407 36561 25463
rect 36489 25373 36508 25407
rect 36542 25373 36561 25407
rect 36489 25317 36561 25373
rect 36489 25283 36508 25317
rect 36542 25283 36561 25317
rect 36489 25227 36561 25283
rect 36489 25193 36508 25227
rect 36542 25193 36561 25227
rect 36489 25137 36561 25193
rect 36489 25103 36508 25137
rect 36542 25103 36561 25137
rect 36623 25740 37317 25799
rect 36623 25706 36684 25740
rect 36718 25712 36774 25740
rect 36808 25712 36864 25740
rect 36898 25712 36954 25740
rect 36730 25706 36774 25712
rect 36830 25706 36864 25712
rect 36930 25706 36954 25712
rect 36988 25712 37044 25740
rect 36988 25706 36996 25712
rect 36623 25678 36696 25706
rect 36730 25678 36796 25706
rect 36830 25678 36896 25706
rect 36930 25678 36996 25706
rect 37030 25706 37044 25712
rect 37078 25712 37134 25740
rect 37078 25706 37096 25712
rect 37030 25678 37096 25706
rect 37130 25706 37134 25712
rect 37168 25712 37224 25740
rect 37168 25706 37196 25712
rect 37258 25706 37317 25740
rect 37130 25678 37196 25706
rect 37230 25678 37317 25706
rect 36623 25650 37317 25678
rect 36623 25616 36684 25650
rect 36718 25616 36774 25650
rect 36808 25616 36864 25650
rect 36898 25616 36954 25650
rect 36988 25616 37044 25650
rect 37078 25616 37134 25650
rect 37168 25616 37224 25650
rect 37258 25616 37317 25650
rect 36623 25612 37317 25616
rect 36623 25578 36696 25612
rect 36730 25578 36796 25612
rect 36830 25578 36896 25612
rect 36930 25578 36996 25612
rect 37030 25578 37096 25612
rect 37130 25578 37196 25612
rect 37230 25578 37317 25612
rect 36623 25560 37317 25578
rect 36623 25526 36684 25560
rect 36718 25526 36774 25560
rect 36808 25526 36864 25560
rect 36898 25526 36954 25560
rect 36988 25526 37044 25560
rect 37078 25526 37134 25560
rect 37168 25526 37224 25560
rect 37258 25526 37317 25560
rect 36623 25512 37317 25526
rect 36623 25478 36696 25512
rect 36730 25478 36796 25512
rect 36830 25478 36896 25512
rect 36930 25478 36996 25512
rect 37030 25478 37096 25512
rect 37130 25478 37196 25512
rect 37230 25478 37317 25512
rect 36623 25470 37317 25478
rect 36623 25436 36684 25470
rect 36718 25436 36774 25470
rect 36808 25436 36864 25470
rect 36898 25436 36954 25470
rect 36988 25436 37044 25470
rect 37078 25436 37134 25470
rect 37168 25436 37224 25470
rect 37258 25436 37317 25470
rect 36623 25412 37317 25436
rect 36623 25380 36696 25412
rect 36730 25380 36796 25412
rect 36830 25380 36896 25412
rect 36930 25380 36996 25412
rect 36623 25346 36684 25380
rect 36730 25378 36774 25380
rect 36830 25378 36864 25380
rect 36930 25378 36954 25380
rect 36718 25346 36774 25378
rect 36808 25346 36864 25378
rect 36898 25346 36954 25378
rect 36988 25378 36996 25380
rect 37030 25380 37096 25412
rect 37030 25378 37044 25380
rect 36988 25346 37044 25378
rect 37078 25378 37096 25380
rect 37130 25380 37196 25412
rect 37230 25380 37317 25412
rect 37130 25378 37134 25380
rect 37078 25346 37134 25378
rect 37168 25378 37196 25380
rect 37168 25346 37224 25378
rect 37258 25346 37317 25380
rect 36623 25312 37317 25346
rect 36623 25290 36696 25312
rect 36730 25290 36796 25312
rect 36830 25290 36896 25312
rect 36930 25290 36996 25312
rect 36623 25256 36684 25290
rect 36730 25278 36774 25290
rect 36830 25278 36864 25290
rect 36930 25278 36954 25290
rect 36718 25256 36774 25278
rect 36808 25256 36864 25278
rect 36898 25256 36954 25278
rect 36988 25278 36996 25290
rect 37030 25290 37096 25312
rect 37030 25278 37044 25290
rect 36988 25256 37044 25278
rect 37078 25278 37096 25290
rect 37130 25290 37196 25312
rect 37230 25290 37317 25312
rect 37130 25278 37134 25290
rect 37078 25256 37134 25278
rect 37168 25278 37196 25290
rect 37168 25256 37224 25278
rect 37258 25256 37317 25290
rect 36623 25212 37317 25256
rect 36623 25200 36696 25212
rect 36730 25200 36796 25212
rect 36830 25200 36896 25212
rect 36930 25200 36996 25212
rect 36623 25166 36684 25200
rect 36730 25178 36774 25200
rect 36830 25178 36864 25200
rect 36930 25178 36954 25200
rect 36718 25166 36774 25178
rect 36808 25166 36864 25178
rect 36898 25166 36954 25178
rect 36988 25178 36996 25200
rect 37030 25200 37096 25212
rect 37030 25178 37044 25200
rect 36988 25166 37044 25178
rect 37078 25178 37096 25200
rect 37130 25200 37196 25212
rect 37230 25200 37317 25212
rect 37130 25178 37134 25200
rect 37078 25166 37134 25178
rect 37168 25178 37196 25200
rect 37168 25166 37224 25178
rect 37258 25166 37317 25200
rect 36623 25105 37317 25166
rect 37379 25748 37451 25804
rect 37379 25714 37398 25748
rect 37432 25714 37451 25748
rect 37379 25658 37451 25714
rect 37379 25624 37398 25658
rect 37432 25624 37451 25658
rect 37379 25568 37451 25624
rect 37379 25534 37398 25568
rect 37432 25534 37451 25568
rect 37379 25478 37451 25534
rect 37379 25444 37398 25478
rect 37432 25444 37451 25478
rect 37379 25388 37451 25444
rect 37379 25354 37398 25388
rect 37432 25354 37451 25388
rect 37379 25298 37451 25354
rect 37379 25264 37398 25298
rect 37432 25264 37451 25298
rect 37379 25208 37451 25264
rect 37379 25174 37398 25208
rect 37432 25174 37451 25208
rect 37379 25118 37451 25174
rect 36489 25043 36561 25103
rect 37379 25084 37398 25118
rect 37432 25084 37451 25118
rect 37379 25043 37451 25084
rect 36489 25024 37451 25043
rect 36489 24990 36586 25024
rect 36620 24990 36676 25024
rect 36710 24990 36766 25024
rect 36800 24990 36856 25024
rect 36890 24990 36946 25024
rect 36980 24990 37036 25024
rect 37070 24990 37126 25024
rect 37160 24990 37216 25024
rect 37250 24990 37306 25024
rect 37340 24990 37451 25024
rect 36489 24971 37451 24990
rect 37515 25914 37547 25948
rect 37581 25914 37700 25948
rect 37734 25914 37765 25948
rect 38855 25948 38954 25997
rect 37515 25858 37765 25914
rect 37515 25824 37547 25858
rect 37581 25824 37700 25858
rect 37734 25824 37765 25858
rect 37515 25768 37765 25824
rect 37515 25734 37547 25768
rect 37581 25734 37700 25768
rect 37734 25734 37765 25768
rect 37515 25678 37765 25734
rect 37515 25644 37547 25678
rect 37581 25644 37700 25678
rect 37734 25644 37765 25678
rect 37515 25588 37765 25644
rect 37515 25554 37547 25588
rect 37581 25554 37700 25588
rect 37734 25554 37765 25588
rect 37515 25498 37765 25554
rect 37515 25464 37547 25498
rect 37581 25464 37700 25498
rect 37734 25464 37765 25498
rect 37515 25408 37765 25464
rect 37515 25374 37547 25408
rect 37581 25374 37700 25408
rect 37734 25374 37765 25408
rect 37515 25318 37765 25374
rect 37515 25284 37547 25318
rect 37581 25284 37700 25318
rect 37734 25284 37765 25318
rect 37515 25228 37765 25284
rect 37515 25194 37547 25228
rect 37581 25194 37700 25228
rect 37734 25194 37765 25228
rect 37515 25138 37765 25194
rect 37515 25104 37547 25138
rect 37581 25104 37700 25138
rect 37734 25104 37765 25138
rect 37515 25048 37765 25104
rect 37515 25014 37547 25048
rect 37581 25014 37700 25048
rect 37734 25014 37765 25048
rect 36175 24924 36207 24958
rect 36241 24924 36360 24958
rect 36394 24924 36425 24958
rect 36175 24907 36425 24924
rect 37515 24958 37765 25014
rect 37829 25916 38791 25933
rect 37829 25882 37850 25916
rect 37884 25882 37940 25916
rect 37974 25914 38030 25916
rect 38064 25914 38120 25916
rect 38154 25914 38210 25916
rect 38244 25914 38300 25916
rect 38334 25914 38390 25916
rect 38424 25914 38480 25916
rect 38514 25914 38570 25916
rect 38604 25914 38660 25916
rect 38694 25914 38750 25916
rect 37994 25882 38030 25914
rect 38084 25882 38120 25914
rect 38174 25882 38210 25914
rect 38264 25882 38300 25914
rect 38354 25882 38390 25914
rect 38444 25882 38480 25914
rect 38534 25882 38570 25914
rect 38624 25882 38660 25914
rect 38714 25882 38750 25914
rect 38784 25882 38791 25916
rect 37829 25880 37960 25882
rect 37994 25880 38050 25882
rect 38084 25880 38140 25882
rect 38174 25880 38230 25882
rect 38264 25880 38320 25882
rect 38354 25880 38410 25882
rect 38444 25880 38500 25882
rect 38534 25880 38590 25882
rect 38624 25880 38680 25882
rect 38714 25880 38791 25882
rect 37829 25861 38791 25880
rect 37829 25857 37901 25861
rect 37829 25823 37848 25857
rect 37882 25823 37901 25857
rect 37829 25767 37901 25823
rect 38719 25838 38791 25861
rect 38719 25804 38738 25838
rect 38772 25804 38791 25838
rect 37829 25733 37848 25767
rect 37882 25733 37901 25767
rect 37829 25677 37901 25733
rect 37829 25643 37848 25677
rect 37882 25643 37901 25677
rect 37829 25587 37901 25643
rect 37829 25553 37848 25587
rect 37882 25553 37901 25587
rect 37829 25497 37901 25553
rect 37829 25463 37848 25497
rect 37882 25463 37901 25497
rect 37829 25407 37901 25463
rect 37829 25373 37848 25407
rect 37882 25373 37901 25407
rect 37829 25317 37901 25373
rect 37829 25283 37848 25317
rect 37882 25283 37901 25317
rect 37829 25227 37901 25283
rect 37829 25193 37848 25227
rect 37882 25193 37901 25227
rect 37829 25137 37901 25193
rect 37829 25103 37848 25137
rect 37882 25103 37901 25137
rect 37963 25740 38657 25799
rect 37963 25706 38024 25740
rect 38058 25712 38114 25740
rect 38148 25712 38204 25740
rect 38238 25712 38294 25740
rect 38070 25706 38114 25712
rect 38170 25706 38204 25712
rect 38270 25706 38294 25712
rect 38328 25712 38384 25740
rect 38328 25706 38336 25712
rect 37963 25678 38036 25706
rect 38070 25678 38136 25706
rect 38170 25678 38236 25706
rect 38270 25678 38336 25706
rect 38370 25706 38384 25712
rect 38418 25712 38474 25740
rect 38418 25706 38436 25712
rect 38370 25678 38436 25706
rect 38470 25706 38474 25712
rect 38508 25712 38564 25740
rect 38508 25706 38536 25712
rect 38598 25706 38657 25740
rect 38470 25678 38536 25706
rect 38570 25678 38657 25706
rect 37963 25650 38657 25678
rect 37963 25616 38024 25650
rect 38058 25616 38114 25650
rect 38148 25616 38204 25650
rect 38238 25616 38294 25650
rect 38328 25616 38384 25650
rect 38418 25616 38474 25650
rect 38508 25616 38564 25650
rect 38598 25616 38657 25650
rect 37963 25612 38657 25616
rect 37963 25578 38036 25612
rect 38070 25578 38136 25612
rect 38170 25578 38236 25612
rect 38270 25578 38336 25612
rect 38370 25578 38436 25612
rect 38470 25578 38536 25612
rect 38570 25578 38657 25612
rect 37963 25560 38657 25578
rect 37963 25526 38024 25560
rect 38058 25526 38114 25560
rect 38148 25526 38204 25560
rect 38238 25526 38294 25560
rect 38328 25526 38384 25560
rect 38418 25526 38474 25560
rect 38508 25526 38564 25560
rect 38598 25526 38657 25560
rect 37963 25512 38657 25526
rect 37963 25478 38036 25512
rect 38070 25478 38136 25512
rect 38170 25478 38236 25512
rect 38270 25478 38336 25512
rect 38370 25478 38436 25512
rect 38470 25478 38536 25512
rect 38570 25478 38657 25512
rect 37963 25470 38657 25478
rect 37963 25436 38024 25470
rect 38058 25436 38114 25470
rect 38148 25436 38204 25470
rect 38238 25436 38294 25470
rect 38328 25436 38384 25470
rect 38418 25436 38474 25470
rect 38508 25436 38564 25470
rect 38598 25436 38657 25470
rect 37963 25412 38657 25436
rect 37963 25380 38036 25412
rect 38070 25380 38136 25412
rect 38170 25380 38236 25412
rect 38270 25380 38336 25412
rect 37963 25346 38024 25380
rect 38070 25378 38114 25380
rect 38170 25378 38204 25380
rect 38270 25378 38294 25380
rect 38058 25346 38114 25378
rect 38148 25346 38204 25378
rect 38238 25346 38294 25378
rect 38328 25378 38336 25380
rect 38370 25380 38436 25412
rect 38370 25378 38384 25380
rect 38328 25346 38384 25378
rect 38418 25378 38436 25380
rect 38470 25380 38536 25412
rect 38570 25380 38657 25412
rect 38470 25378 38474 25380
rect 38418 25346 38474 25378
rect 38508 25378 38536 25380
rect 38508 25346 38564 25378
rect 38598 25346 38657 25380
rect 37963 25312 38657 25346
rect 37963 25290 38036 25312
rect 38070 25290 38136 25312
rect 38170 25290 38236 25312
rect 38270 25290 38336 25312
rect 37963 25256 38024 25290
rect 38070 25278 38114 25290
rect 38170 25278 38204 25290
rect 38270 25278 38294 25290
rect 38058 25256 38114 25278
rect 38148 25256 38204 25278
rect 38238 25256 38294 25278
rect 38328 25278 38336 25290
rect 38370 25290 38436 25312
rect 38370 25278 38384 25290
rect 38328 25256 38384 25278
rect 38418 25278 38436 25290
rect 38470 25290 38536 25312
rect 38570 25290 38657 25312
rect 38470 25278 38474 25290
rect 38418 25256 38474 25278
rect 38508 25278 38536 25290
rect 38508 25256 38564 25278
rect 38598 25256 38657 25290
rect 37963 25212 38657 25256
rect 37963 25200 38036 25212
rect 38070 25200 38136 25212
rect 38170 25200 38236 25212
rect 38270 25200 38336 25212
rect 37963 25166 38024 25200
rect 38070 25178 38114 25200
rect 38170 25178 38204 25200
rect 38270 25178 38294 25200
rect 38058 25166 38114 25178
rect 38148 25166 38204 25178
rect 38238 25166 38294 25178
rect 38328 25178 38336 25200
rect 38370 25200 38436 25212
rect 38370 25178 38384 25200
rect 38328 25166 38384 25178
rect 38418 25178 38436 25200
rect 38470 25200 38536 25212
rect 38570 25200 38657 25212
rect 38470 25178 38474 25200
rect 38418 25166 38474 25178
rect 38508 25178 38536 25200
rect 38508 25166 38564 25178
rect 38598 25166 38657 25200
rect 37963 25105 38657 25166
rect 38719 25748 38791 25804
rect 38719 25714 38738 25748
rect 38772 25714 38791 25748
rect 38719 25658 38791 25714
rect 38719 25624 38738 25658
rect 38772 25624 38791 25658
rect 38719 25568 38791 25624
rect 38719 25534 38738 25568
rect 38772 25534 38791 25568
rect 38719 25478 38791 25534
rect 38719 25444 38738 25478
rect 38772 25444 38791 25478
rect 38719 25388 38791 25444
rect 38719 25354 38738 25388
rect 38772 25354 38791 25388
rect 38719 25298 38791 25354
rect 38719 25264 38738 25298
rect 38772 25264 38791 25298
rect 38719 25208 38791 25264
rect 38719 25174 38738 25208
rect 38772 25174 38791 25208
rect 38719 25118 38791 25174
rect 37829 25043 37901 25103
rect 38719 25084 38738 25118
rect 38772 25084 38791 25118
rect 38719 25043 38791 25084
rect 37829 25024 38791 25043
rect 37829 24990 37926 25024
rect 37960 24990 38016 25024
rect 38050 24990 38106 25024
rect 38140 24990 38196 25024
rect 38230 24990 38286 25024
rect 38320 24990 38376 25024
rect 38410 24990 38466 25024
rect 38500 24990 38556 25024
rect 38590 24990 38646 25024
rect 38680 24990 38791 25024
rect 37829 24971 38791 24990
rect 38855 25914 38887 25948
rect 38921 25914 38954 25948
rect 38855 25858 38954 25914
rect 38855 25824 38887 25858
rect 38921 25824 38954 25858
rect 38855 25768 38954 25824
rect 38855 25734 38887 25768
rect 38921 25734 38954 25768
rect 38855 25678 38954 25734
rect 38855 25644 38887 25678
rect 38921 25644 38954 25678
rect 38855 25588 38954 25644
rect 38855 25554 38887 25588
rect 38921 25554 38954 25588
rect 38855 25498 38954 25554
rect 38855 25464 38887 25498
rect 38921 25464 38954 25498
rect 38855 25408 38954 25464
rect 38855 25374 38887 25408
rect 38921 25374 38954 25408
rect 38855 25318 38954 25374
rect 38855 25284 38887 25318
rect 38921 25284 38954 25318
rect 38855 25228 38954 25284
rect 38855 25194 38887 25228
rect 38921 25194 38954 25228
rect 40658 25443 41274 25482
rect 40658 25341 40745 25443
rect 41187 25341 41274 25443
rect 38855 25138 38954 25194
rect 38855 25104 38887 25138
rect 38921 25104 38954 25138
rect 38855 25048 38954 25104
rect 38855 25014 38887 25048
rect 38921 25014 38954 25048
rect 37515 24924 37547 24958
rect 37581 24924 37700 24958
rect 37734 24924 37765 24958
rect 37515 24907 37765 24924
rect 38855 24958 38954 25014
rect 38855 24924 38887 24958
rect 38921 24924 38954 24958
rect 38855 24907 38954 24924
rect 23048 24871 27148 24876
rect 23048 24863 23305 24871
rect 23048 24829 23151 24863
rect 23185 24837 23305 24863
rect 23339 24863 27148 24871
rect 23339 24837 23551 24863
rect 23185 24829 23551 24837
rect 23585 24829 23951 24863
rect 23985 24829 24351 24863
rect 24385 24829 24751 24863
rect 24785 24829 25151 24863
rect 25185 24829 25551 24863
rect 25585 24829 25951 24863
rect 25985 24829 26351 24863
rect 26385 24829 26751 24863
rect 26785 24829 27148 24863
rect 23048 24816 27148 24829
rect 28286 24874 38954 24907
rect 28286 24840 28416 24874
rect 28450 24840 28506 24874
rect 28540 24840 28596 24874
rect 28630 24840 28686 24874
rect 28720 24840 28776 24874
rect 28810 24840 28866 24874
rect 28900 24840 28956 24874
rect 28990 24840 29046 24874
rect 29080 24840 29136 24874
rect 29170 24840 29226 24874
rect 29260 24840 29316 24874
rect 29350 24840 29406 24874
rect 29440 24840 29756 24874
rect 29790 24840 29846 24874
rect 29880 24840 29936 24874
rect 29970 24840 30026 24874
rect 30060 24840 30116 24874
rect 30150 24840 30206 24874
rect 30240 24840 30296 24874
rect 30330 24840 30386 24874
rect 30420 24840 30476 24874
rect 30510 24840 30566 24874
rect 30600 24840 30656 24874
rect 30690 24840 30746 24874
rect 30780 24840 31096 24874
rect 31130 24840 31186 24874
rect 31220 24840 31276 24874
rect 31310 24840 31366 24874
rect 31400 24840 31456 24874
rect 31490 24840 31546 24874
rect 31580 24840 31636 24874
rect 31670 24840 31726 24874
rect 31760 24840 31816 24874
rect 31850 24840 31906 24874
rect 31940 24840 31996 24874
rect 32030 24840 32086 24874
rect 32120 24840 32436 24874
rect 32470 24840 32526 24874
rect 32560 24840 32616 24874
rect 32650 24840 32706 24874
rect 32740 24840 32796 24874
rect 32830 24840 32886 24874
rect 32920 24840 32976 24874
rect 33010 24840 33066 24874
rect 33100 24840 33156 24874
rect 33190 24840 33246 24874
rect 33280 24840 33336 24874
rect 33370 24840 33426 24874
rect 33460 24840 33776 24874
rect 33810 24840 33866 24874
rect 33900 24840 33956 24874
rect 33990 24840 34046 24874
rect 34080 24840 34136 24874
rect 34170 24840 34226 24874
rect 34260 24840 34316 24874
rect 34350 24840 34406 24874
rect 34440 24840 34496 24874
rect 34530 24840 34586 24874
rect 34620 24840 34676 24874
rect 34710 24840 34766 24874
rect 34800 24840 35116 24874
rect 35150 24840 35206 24874
rect 35240 24840 35296 24874
rect 35330 24840 35386 24874
rect 35420 24840 35476 24874
rect 35510 24840 35566 24874
rect 35600 24840 35656 24874
rect 35690 24840 35746 24874
rect 35780 24840 35836 24874
rect 35870 24840 35926 24874
rect 35960 24840 36016 24874
rect 36050 24840 36106 24874
rect 36140 24840 36456 24874
rect 36490 24840 36546 24874
rect 36580 24840 36636 24874
rect 36670 24840 36726 24874
rect 36760 24840 36816 24874
rect 36850 24840 36906 24874
rect 36940 24840 36996 24874
rect 37030 24840 37086 24874
rect 37120 24840 37176 24874
rect 37210 24840 37266 24874
rect 37300 24840 37356 24874
rect 37390 24840 37446 24874
rect 37480 24840 37796 24874
rect 37830 24840 37886 24874
rect 37920 24840 37976 24874
rect 38010 24840 38066 24874
rect 38100 24840 38156 24874
rect 38190 24840 38246 24874
rect 38280 24840 38336 24874
rect 38370 24840 38426 24874
rect 38460 24840 38516 24874
rect 38550 24840 38606 24874
rect 38640 24840 38696 24874
rect 38730 24840 38786 24874
rect 38820 24840 38954 24874
rect 28286 24808 38954 24840
rect 9542 24722 15166 24782
rect 9542 24667 15166 24676
rect 9542 24633 9689 24667
rect 9723 24663 12541 24667
rect 12575 24663 15166 24667
rect 9723 24633 9725 24663
rect 9542 24629 9725 24633
rect 9759 24629 10125 24663
rect 10159 24629 10525 24663
rect 10559 24629 10925 24663
rect 10959 24629 11325 24663
rect 11359 24629 11725 24663
rect 11759 24629 12125 24663
rect 12159 24629 12525 24663
rect 12575 24633 12925 24663
rect 12559 24629 12925 24633
rect 12959 24629 13325 24663
rect 13359 24629 13725 24663
rect 13759 24629 14125 24663
rect 14159 24629 14525 24663
rect 14559 24629 14925 24663
rect 14959 24629 15166 24663
rect 9542 24616 15166 24629
rect 22898 24669 22958 24752
rect 22898 24635 22911 24669
rect 22945 24635 22958 24669
rect 22898 24542 22958 24635
rect 23948 24639 24108 24662
rect 23948 24605 24013 24639
rect 24047 24605 24108 24639
rect 23948 24542 24108 24605
rect 25248 24639 25408 24662
rect 25248 24605 25313 24639
rect 25347 24605 25408 24639
rect 25248 24542 25408 24605
rect 40658 24542 41274 25341
rect 41754 25197 42186 25587
rect 6720 24529 9160 24542
rect 6720 24495 6903 24529
rect 6937 24495 7103 24529
rect 7137 24495 7303 24529
rect 7337 24495 7503 24529
rect 7537 24495 7703 24529
rect 7737 24495 7903 24529
rect 7937 24495 8103 24529
rect 8137 24495 8303 24529
rect 8337 24495 8503 24529
rect 8537 24495 8703 24529
rect 8737 24495 8903 24529
rect 8937 24495 9160 24529
rect 6720 24482 9160 24495
rect 9444 24529 15166 24542
rect 9444 24495 9725 24529
rect 9759 24495 10125 24529
rect 10159 24495 10525 24529
rect 10559 24495 10925 24529
rect 10959 24495 11325 24529
rect 11359 24495 11725 24529
rect 11759 24495 12125 24529
rect 12159 24495 12525 24529
rect 12559 24495 12925 24529
rect 12959 24495 13325 24529
rect 13359 24495 13725 24529
rect 13759 24495 14125 24529
rect 14159 24495 14525 24529
rect 14559 24495 14925 24529
rect 14959 24495 15166 24529
rect 9444 24482 15166 24495
rect 15424 24529 22592 24542
rect 15424 24495 15607 24529
rect 15641 24495 16007 24529
rect 16041 24495 16407 24529
rect 16441 24495 16807 24529
rect 16841 24495 17207 24529
rect 17241 24495 17607 24529
rect 17641 24495 18007 24529
rect 18041 24495 18407 24529
rect 18441 24495 18807 24529
rect 18841 24495 19207 24529
rect 19241 24495 19607 24529
rect 19641 24495 20007 24529
rect 20041 24495 20407 24529
rect 20441 24495 20807 24529
rect 20841 24495 21207 24529
rect 21241 24495 21607 24529
rect 21641 24495 22007 24529
rect 22041 24495 22407 24529
rect 22441 24495 22592 24529
rect 15424 24482 22592 24495
rect 22870 24529 27148 24542
rect 22870 24495 23151 24529
rect 23185 24495 23551 24529
rect 23585 24495 23951 24529
rect 23985 24495 24351 24529
rect 24385 24495 24751 24529
rect 24785 24495 25151 24529
rect 25185 24495 25551 24529
rect 25585 24495 25951 24529
rect 25985 24495 26351 24529
rect 26385 24495 26751 24529
rect 26785 24495 27148 24529
rect 22870 24482 27148 24495
rect 28260 24529 38980 24542
rect 28260 24495 28443 24529
rect 28477 24495 28643 24529
rect 28677 24495 28843 24529
rect 28877 24495 29043 24529
rect 29077 24495 29243 24529
rect 29277 24495 29443 24529
rect 29477 24495 29643 24529
rect 29677 24495 29843 24529
rect 29877 24495 30043 24529
rect 30077 24495 30243 24529
rect 30277 24495 30443 24529
rect 30477 24495 30643 24529
rect 30677 24495 30843 24529
rect 30877 24495 31043 24529
rect 31077 24495 31243 24529
rect 31277 24495 31443 24529
rect 31477 24495 31643 24529
rect 31677 24495 31843 24529
rect 31877 24495 32043 24529
rect 32077 24495 32243 24529
rect 32277 24495 32443 24529
rect 32477 24495 32643 24529
rect 32677 24495 32843 24529
rect 32877 24495 33043 24529
rect 33077 24495 33243 24529
rect 33277 24495 33443 24529
rect 33477 24495 33643 24529
rect 33677 24495 33843 24529
rect 33877 24495 34043 24529
rect 34077 24495 34243 24529
rect 34277 24495 34443 24529
rect 34477 24495 34643 24529
rect 34677 24495 34843 24529
rect 34877 24495 35043 24529
rect 35077 24495 35243 24529
rect 35277 24495 35443 24529
rect 35477 24495 35643 24529
rect 35677 24495 35843 24529
rect 35877 24495 36043 24529
rect 36077 24495 36243 24529
rect 36277 24495 36443 24529
rect 36477 24495 36643 24529
rect 36677 24495 36843 24529
rect 36877 24495 37043 24529
rect 37077 24495 37243 24529
rect 37277 24495 37443 24529
rect 37477 24495 37643 24529
rect 37677 24495 37843 24529
rect 37877 24495 38043 24529
rect 38077 24495 38243 24529
rect 38277 24495 38443 24529
rect 38477 24495 38643 24529
rect 38677 24495 38843 24529
rect 38877 24495 38980 24529
rect 28260 24482 38980 24495
rect 39746 24529 42186 24542
rect 39746 24495 39929 24529
rect 39963 24495 40129 24529
rect 40163 24495 40329 24529
rect 40363 24495 40529 24529
rect 40563 24495 40729 24529
rect 40763 24495 40929 24529
rect 40963 24495 41129 24529
rect 41163 24495 41329 24529
rect 41363 24495 41529 24529
rect 41563 24495 41729 24529
rect 41763 24495 41929 24529
rect 41963 24495 42186 24529
rect 39746 24482 42186 24495
rect 7582 22649 13304 22662
rect 7582 22615 7863 22649
rect 7897 22615 8263 22649
rect 8297 22615 8663 22649
rect 8697 22615 9063 22649
rect 9097 22615 9463 22649
rect 9497 22615 9863 22649
rect 9897 22615 10263 22649
rect 10297 22615 10663 22649
rect 10697 22615 11063 22649
rect 11097 22615 11463 22649
rect 11497 22615 11863 22649
rect 11897 22615 12263 22649
rect 12297 22615 12663 22649
rect 12697 22615 13063 22649
rect 13097 22615 13304 22649
rect 7582 22602 13304 22615
rect 13562 22649 20730 22662
rect 13562 22615 13745 22649
rect 13779 22615 14145 22649
rect 14179 22615 14545 22649
rect 14579 22615 14945 22649
rect 14979 22615 15345 22649
rect 15379 22615 15745 22649
rect 15779 22615 16145 22649
rect 16179 22615 16545 22649
rect 16579 22615 16945 22649
rect 16979 22615 17345 22649
rect 17379 22615 17745 22649
rect 17779 22615 18145 22649
rect 18179 22615 18545 22649
rect 18579 22615 18945 22649
rect 18979 22615 19345 22649
rect 19379 22615 19745 22649
rect 19779 22615 20145 22649
rect 20179 22615 20545 22649
rect 20579 22615 20730 22649
rect 13562 22602 20730 22615
rect 21008 22649 22348 22662
rect 21008 22615 21191 22649
rect 21225 22615 21391 22649
rect 21425 22615 21591 22649
rect 21625 22615 21791 22649
rect 21825 22615 21991 22649
rect 22025 22615 22191 22649
rect 22225 22615 22348 22649
rect 21008 22602 22348 22615
rect 22870 22649 27148 22662
rect 22870 22615 23151 22649
rect 23185 22615 23551 22649
rect 23585 22615 23951 22649
rect 23985 22615 24351 22649
rect 24385 22615 24751 22649
rect 24785 22615 25151 22649
rect 25185 22615 25551 22649
rect 25585 22615 25951 22649
rect 25985 22615 26351 22649
rect 26385 22615 26751 22649
rect 26785 22615 27148 22649
rect 22870 22602 27148 22615
rect 28260 22649 38980 22662
rect 28260 22615 28443 22649
rect 28477 22615 28643 22649
rect 28677 22615 28843 22649
rect 28877 22615 29043 22649
rect 29077 22615 29243 22649
rect 29277 22615 29443 22649
rect 29477 22615 29643 22649
rect 29677 22615 29843 22649
rect 29877 22615 30043 22649
rect 30077 22615 30243 22649
rect 30277 22615 30443 22649
rect 30477 22615 30643 22649
rect 30677 22615 30843 22649
rect 30877 22615 31043 22649
rect 31077 22615 31243 22649
rect 31277 22615 31443 22649
rect 31477 22615 31643 22649
rect 31677 22615 31843 22649
rect 31877 22615 32043 22649
rect 32077 22615 32243 22649
rect 32277 22615 32443 22649
rect 32477 22615 32643 22649
rect 32677 22615 32843 22649
rect 32877 22615 33043 22649
rect 33077 22615 33243 22649
rect 33277 22615 33443 22649
rect 33477 22615 33643 22649
rect 33677 22615 33843 22649
rect 33877 22615 34043 22649
rect 34077 22615 34243 22649
rect 34277 22615 34443 22649
rect 34477 22615 34643 22649
rect 34677 22615 34843 22649
rect 34877 22615 35043 22649
rect 35077 22615 35243 22649
rect 35277 22615 35443 22649
rect 35477 22615 35643 22649
rect 35677 22615 35843 22649
rect 35877 22615 36043 22649
rect 36077 22615 36243 22649
rect 36277 22615 36443 22649
rect 36477 22615 36643 22649
rect 36677 22615 36843 22649
rect 36877 22615 37043 22649
rect 37077 22615 37243 22649
rect 37277 22615 37443 22649
rect 37477 22615 37643 22649
rect 37677 22615 37843 22649
rect 37877 22615 38043 22649
rect 38077 22615 38243 22649
rect 38277 22615 38443 22649
rect 38477 22615 38643 22649
rect 38677 22615 38843 22649
rect 38877 22615 38980 22649
rect 28260 22602 38980 22615
rect 39746 22649 42186 22662
rect 39746 22615 39929 22649
rect 39963 22615 40129 22649
rect 40163 22615 40329 22649
rect 40363 22615 40529 22649
rect 40563 22615 40729 22649
rect 40763 22615 40929 22649
rect 40963 22615 41129 22649
rect 41163 22615 41329 22649
rect 41363 22615 41529 22649
rect 41563 22615 41729 22649
rect 41763 22615 41929 22649
rect 41963 22615 42186 22649
rect 39746 22602 42186 22615
rect 7610 22509 7670 22602
rect 8658 22559 8818 22602
rect 8658 22525 8723 22559
rect 8757 22525 8818 22559
rect 8658 22522 8818 22525
rect 9958 22559 10118 22602
rect 9958 22525 10023 22559
rect 10057 22525 10118 22559
rect 9958 22522 10118 22525
rect 11258 22559 11418 22602
rect 11258 22525 11323 22559
rect 11357 22525 11418 22559
rect 11258 22522 11418 22525
rect 7610 22475 7623 22509
rect 7657 22475 7670 22509
rect 22968 22491 27148 22502
rect 7610 22392 7670 22475
rect 7740 22457 8309 22482
rect 8343 22457 13304 22482
rect 7740 22442 13304 22457
rect 22968 22457 26433 22491
rect 26467 22457 27148 22491
rect 22968 22442 27148 22457
rect 7727 22381 7761 22401
rect 7727 22313 7761 22347
rect 7727 22245 7761 22275
rect 7727 22177 7761 22203
rect 7727 22109 7761 22131
rect 7727 22041 7761 22059
rect 7727 21973 7761 21987
rect 7727 21905 7761 21915
rect 7727 21837 7761 21843
rect 7727 21769 7761 21771
rect 7727 21733 7761 21735
rect 7727 21661 7761 21667
rect 7727 21589 7761 21599
rect 7727 21517 7761 21531
rect 7727 21445 7761 21463
rect 7727 21373 7761 21395
rect 7727 21301 7761 21327
rect 7727 21229 7761 21259
rect 7727 21157 7761 21191
rect 7727 21022 7761 21123
rect 8185 22381 8219 22442
rect 8185 22313 8219 22347
rect 8185 22245 8219 22275
rect 8185 22177 8219 22203
rect 8185 22109 8219 22131
rect 8185 22041 8219 22059
rect 8185 21973 8219 21987
rect 8185 21905 8219 21915
rect 8185 21837 8219 21843
rect 8185 21769 8219 21771
rect 8185 21733 8219 21735
rect 8185 21661 8219 21667
rect 8185 21589 8219 21599
rect 8185 21517 8219 21531
rect 8185 21445 8219 21463
rect 8185 21373 8219 21395
rect 8185 21301 8219 21327
rect 8185 21229 8219 21259
rect 8185 21157 8219 21191
rect 8185 21103 8219 21123
rect 8643 22381 8677 22401
rect 8643 22313 8677 22347
rect 8643 22245 8677 22275
rect 8643 22177 8677 22203
rect 8643 22109 8677 22131
rect 8643 22041 8677 22059
rect 8643 21973 8677 21987
rect 8643 21905 8677 21915
rect 8643 21837 8677 21843
rect 8643 21769 8677 21771
rect 8643 21733 8677 21735
rect 8643 21661 8677 21667
rect 8643 21589 8677 21599
rect 8643 21517 8677 21531
rect 8643 21445 8677 21463
rect 8643 21373 8677 21395
rect 8643 21301 8677 21327
rect 8643 21229 8677 21259
rect 8643 21157 8677 21191
rect 8643 21022 8677 21123
rect 9101 22381 9135 22442
rect 9101 22313 9135 22347
rect 9101 22245 9135 22275
rect 9101 22177 9135 22203
rect 9101 22109 9135 22131
rect 9101 22041 9135 22059
rect 9101 21973 9135 21987
rect 9101 21905 9135 21915
rect 9101 21837 9135 21843
rect 9101 21769 9135 21771
rect 9101 21733 9135 21735
rect 9101 21661 9135 21667
rect 9101 21589 9135 21599
rect 9101 21517 9135 21531
rect 9101 21445 9135 21463
rect 9101 21373 9135 21395
rect 9101 21301 9135 21327
rect 9101 21229 9135 21259
rect 9101 21157 9135 21191
rect 9101 21103 9135 21123
rect 9559 22381 9593 22401
rect 9559 22313 9593 22347
rect 9559 22245 9593 22275
rect 9559 22177 9593 22203
rect 9559 22109 9593 22131
rect 9559 22041 9593 22059
rect 9559 21973 9593 21987
rect 9559 21905 9593 21915
rect 9559 21837 9593 21843
rect 9559 21769 9593 21771
rect 9559 21733 9593 21735
rect 9559 21661 9593 21667
rect 9559 21589 9593 21599
rect 9559 21517 9593 21531
rect 9559 21445 9593 21463
rect 9559 21373 9593 21395
rect 9559 21301 9593 21327
rect 9559 21229 9593 21259
rect 9559 21157 9593 21191
rect 9559 21022 9593 21123
rect 10017 22381 10051 22442
rect 10017 22313 10051 22347
rect 10017 22245 10051 22275
rect 10017 22177 10051 22203
rect 10017 22109 10051 22131
rect 10017 22041 10051 22059
rect 10017 21973 10051 21987
rect 10017 21905 10051 21915
rect 10017 21837 10051 21843
rect 10017 21769 10051 21771
rect 10017 21733 10051 21735
rect 10017 21661 10051 21667
rect 10017 21589 10051 21599
rect 10017 21517 10051 21531
rect 10017 21445 10051 21463
rect 10017 21373 10051 21395
rect 10017 21301 10051 21327
rect 10017 21229 10051 21259
rect 10017 21157 10051 21191
rect 10017 21103 10051 21123
rect 10475 22381 10509 22401
rect 10475 22313 10509 22347
rect 10475 22245 10509 22275
rect 10475 22177 10509 22203
rect 10475 22109 10509 22131
rect 10475 22041 10509 22059
rect 10475 21973 10509 21987
rect 10475 21905 10509 21915
rect 10475 21837 10509 21843
rect 10475 21769 10509 21771
rect 10475 21733 10509 21735
rect 10475 21661 10509 21667
rect 10475 21589 10509 21599
rect 10475 21517 10509 21531
rect 10475 21445 10509 21463
rect 10475 21373 10509 21395
rect 10475 21301 10509 21327
rect 10475 21229 10509 21259
rect 10475 21157 10509 21191
rect 10475 21022 10509 21123
rect 10933 22381 10967 22442
rect 10933 22313 10967 22347
rect 10933 22245 10967 22275
rect 10933 22177 10967 22203
rect 10933 22109 10967 22131
rect 10933 22041 10967 22059
rect 10933 21973 10967 21987
rect 10933 21905 10967 21915
rect 10933 21837 10967 21843
rect 10933 21769 10967 21771
rect 10933 21733 10967 21735
rect 10933 21661 10967 21667
rect 10933 21589 10967 21599
rect 10933 21517 10967 21531
rect 10933 21445 10967 21463
rect 10933 21373 10967 21395
rect 10933 21301 10967 21327
rect 10933 21229 10967 21259
rect 10933 21157 10967 21191
rect 10933 21103 10967 21123
rect 11391 22381 11425 22401
rect 11391 22313 11425 22347
rect 11391 22245 11425 22275
rect 11391 22177 11425 22203
rect 11391 22109 11425 22131
rect 11391 22041 11425 22059
rect 11391 21973 11425 21987
rect 11391 21905 11425 21915
rect 11391 21837 11425 21843
rect 11391 21769 11425 21771
rect 11391 21733 11425 21735
rect 11391 21661 11425 21667
rect 11391 21589 11425 21599
rect 11391 21517 11425 21531
rect 11391 21445 11425 21463
rect 11391 21373 11425 21395
rect 11391 21301 11425 21327
rect 11391 21229 11425 21259
rect 11391 21157 11425 21191
rect 11391 21022 11425 21123
rect 11849 22381 11883 22442
rect 11849 22313 11883 22347
rect 11849 22245 11883 22275
rect 11849 22177 11883 22203
rect 11849 22109 11883 22131
rect 11849 22041 11883 22059
rect 11849 21973 11883 21987
rect 11849 21905 11883 21915
rect 11849 21837 11883 21843
rect 11849 21769 11883 21771
rect 11849 21733 11883 21735
rect 11849 21661 11883 21667
rect 11849 21589 11883 21599
rect 11849 21517 11883 21531
rect 11849 21445 11883 21463
rect 11849 21373 11883 21395
rect 11849 21301 11883 21327
rect 11849 21229 11883 21259
rect 11849 21157 11883 21191
rect 11849 21103 11883 21123
rect 12307 22381 12341 22401
rect 12307 22313 12341 22347
rect 12307 22245 12341 22275
rect 12307 22177 12341 22203
rect 12307 22109 12341 22131
rect 12307 22041 12341 22059
rect 12307 21973 12341 21987
rect 12307 21905 12341 21915
rect 12307 21837 12341 21843
rect 12307 21769 12341 21771
rect 12307 21733 12341 21735
rect 12307 21661 12341 21667
rect 12307 21589 12341 21599
rect 12307 21517 12341 21531
rect 12307 21445 12341 21463
rect 12307 21373 12341 21395
rect 12307 21301 12341 21327
rect 12307 21229 12341 21259
rect 12307 21157 12341 21191
rect 12307 21022 12341 21123
rect 12765 22381 12799 22442
rect 12765 22313 12799 22347
rect 12765 22245 12799 22275
rect 12765 22177 12799 22203
rect 12765 22109 12799 22131
rect 12765 22041 12799 22059
rect 12765 21973 12799 21987
rect 12765 21905 12799 21915
rect 12765 21837 12799 21843
rect 12765 21769 12799 21771
rect 12765 21733 12799 21735
rect 12765 21661 12799 21667
rect 12765 21589 12799 21599
rect 12765 21517 12799 21531
rect 12765 21445 12799 21463
rect 12765 21373 12799 21395
rect 12765 21301 12799 21327
rect 12765 21229 12799 21259
rect 12765 21157 12799 21191
rect 12765 21103 12799 21123
rect 13223 22381 13257 22401
rect 13223 22313 13257 22347
rect 13223 22245 13257 22275
rect 13223 22177 13257 22203
rect 13223 22109 13257 22131
rect 13223 22041 13257 22059
rect 13223 21973 13257 21987
rect 13223 21905 13257 21915
rect 13223 21837 13257 21843
rect 13223 21769 13257 21771
rect 13223 21733 13257 21735
rect 13223 21661 13257 21667
rect 13223 21589 13257 21599
rect 13223 21517 13257 21531
rect 13223 21445 13257 21463
rect 13223 21373 13257 21395
rect 13223 21301 13257 21327
rect 13223 21229 13257 21259
rect 13223 21157 13257 21191
rect 13223 21022 13257 21123
rect 21034 22301 22322 22336
rect 21034 22278 21164 22301
rect 21034 22244 21068 22278
rect 21102 22267 21164 22278
rect 21198 22267 21254 22301
rect 21288 22267 21344 22301
rect 21378 22267 21434 22301
rect 21468 22267 21524 22301
rect 21558 22267 21614 22301
rect 21648 22267 21704 22301
rect 21738 22267 21794 22301
rect 21828 22267 21884 22301
rect 21918 22267 21974 22301
rect 22008 22267 22064 22301
rect 22098 22267 22154 22301
rect 22188 22278 22322 22301
rect 22188 22267 22255 22278
rect 21102 22244 22255 22267
rect 22289 22244 22322 22278
rect 21034 22237 22322 22244
rect 21034 22188 21133 22237
rect 21034 22154 21068 22188
rect 21102 22154 21133 22188
rect 22223 22188 22322 22237
rect 21034 22098 21133 22154
rect 21034 22064 21068 22098
rect 21102 22064 21133 22098
rect 21034 22008 21133 22064
rect 21034 21974 21068 22008
rect 21102 21974 21133 22008
rect 21034 21918 21133 21974
rect 21034 21884 21068 21918
rect 21102 21884 21133 21918
rect 21034 21828 21133 21884
rect 21034 21794 21068 21828
rect 21102 21794 21133 21828
rect 21034 21738 21133 21794
rect 21034 21704 21068 21738
rect 21102 21704 21133 21738
rect 21034 21648 21133 21704
rect 21034 21614 21068 21648
rect 21102 21614 21133 21648
rect 21034 21558 21133 21614
rect 21034 21524 21068 21558
rect 21102 21524 21133 21558
rect 21034 21468 21133 21524
rect 21034 21434 21068 21468
rect 21102 21434 21133 21468
rect 21034 21378 21133 21434
rect 21034 21344 21068 21378
rect 21102 21344 21133 21378
rect 21034 21288 21133 21344
rect 21034 21254 21068 21288
rect 21102 21254 21133 21288
rect 21197 22154 22159 22173
rect 21197 22120 21328 22154
rect 21362 22120 21418 22154
rect 21452 22120 21508 22154
rect 21542 22120 21598 22154
rect 21632 22120 21688 22154
rect 21722 22120 21778 22154
rect 21812 22120 21868 22154
rect 21902 22120 21958 22154
rect 21992 22120 22048 22154
rect 22082 22120 22159 22154
rect 21197 22101 22159 22120
rect 21197 22097 21269 22101
rect 21197 22063 21216 22097
rect 21250 22063 21269 22097
rect 21197 22007 21269 22063
rect 22087 22078 22159 22101
rect 22087 22044 22106 22078
rect 22140 22044 22159 22078
rect 21197 21973 21216 22007
rect 21250 21973 21269 22007
rect 21197 21917 21269 21973
rect 21197 21883 21216 21917
rect 21250 21883 21269 21917
rect 21197 21827 21269 21883
rect 21197 21793 21216 21827
rect 21250 21793 21269 21827
rect 21197 21737 21269 21793
rect 21197 21703 21216 21737
rect 21250 21703 21269 21737
rect 21197 21647 21269 21703
rect 21197 21613 21216 21647
rect 21250 21613 21269 21647
rect 21197 21557 21269 21613
rect 21197 21523 21216 21557
rect 21250 21523 21269 21557
rect 21197 21467 21269 21523
rect 21197 21433 21216 21467
rect 21250 21433 21269 21467
rect 21197 21377 21269 21433
rect 21197 21343 21216 21377
rect 21250 21343 21269 21377
rect 21331 21980 22025 22039
rect 21331 21946 21392 21980
rect 21426 21952 21482 21980
rect 21516 21952 21572 21980
rect 21606 21952 21662 21980
rect 21438 21946 21482 21952
rect 21538 21946 21572 21952
rect 21638 21946 21662 21952
rect 21696 21952 21752 21980
rect 21696 21946 21704 21952
rect 21331 21918 21404 21946
rect 21438 21918 21504 21946
rect 21538 21918 21604 21946
rect 21638 21918 21704 21946
rect 21738 21946 21752 21952
rect 21786 21952 21842 21980
rect 21786 21946 21804 21952
rect 21738 21918 21804 21946
rect 21838 21946 21842 21952
rect 21876 21952 21932 21980
rect 21876 21946 21904 21952
rect 21966 21946 22025 21980
rect 21838 21918 21904 21946
rect 21938 21918 22025 21946
rect 21331 21890 22025 21918
rect 21331 21856 21392 21890
rect 21426 21856 21482 21890
rect 21516 21856 21572 21890
rect 21606 21856 21662 21890
rect 21696 21856 21752 21890
rect 21786 21856 21842 21890
rect 21876 21856 21932 21890
rect 21966 21856 22025 21890
rect 21331 21852 22025 21856
rect 21331 21818 21404 21852
rect 21438 21818 21504 21852
rect 21538 21818 21604 21852
rect 21638 21818 21704 21852
rect 21738 21818 21804 21852
rect 21838 21818 21904 21852
rect 21938 21818 22025 21852
rect 21331 21800 22025 21818
rect 21331 21766 21392 21800
rect 21426 21766 21482 21800
rect 21516 21766 21572 21800
rect 21606 21766 21662 21800
rect 21696 21766 21752 21800
rect 21786 21766 21842 21800
rect 21876 21766 21932 21800
rect 21966 21766 22025 21800
rect 21331 21752 22025 21766
rect 21331 21718 21404 21752
rect 21438 21718 21504 21752
rect 21538 21718 21604 21752
rect 21638 21718 21704 21752
rect 21738 21718 21804 21752
rect 21838 21718 21904 21752
rect 21938 21718 22025 21752
rect 21331 21710 22025 21718
rect 21331 21676 21392 21710
rect 21426 21676 21482 21710
rect 21516 21676 21572 21710
rect 21606 21676 21662 21710
rect 21696 21676 21752 21710
rect 21786 21676 21842 21710
rect 21876 21676 21932 21710
rect 21966 21676 22025 21710
rect 21331 21652 22025 21676
rect 21331 21620 21404 21652
rect 21438 21620 21504 21652
rect 21538 21620 21604 21652
rect 21638 21620 21704 21652
rect 21331 21586 21392 21620
rect 21438 21618 21482 21620
rect 21538 21618 21572 21620
rect 21638 21618 21662 21620
rect 21426 21586 21482 21618
rect 21516 21586 21572 21618
rect 21606 21586 21662 21618
rect 21696 21618 21704 21620
rect 21738 21620 21804 21652
rect 21738 21618 21752 21620
rect 21696 21586 21752 21618
rect 21786 21618 21804 21620
rect 21838 21620 21904 21652
rect 21938 21620 22025 21652
rect 21838 21618 21842 21620
rect 21786 21586 21842 21618
rect 21876 21618 21904 21620
rect 21876 21586 21932 21618
rect 21966 21586 22025 21620
rect 21331 21552 22025 21586
rect 21331 21530 21404 21552
rect 21438 21530 21504 21552
rect 21538 21530 21604 21552
rect 21638 21530 21704 21552
rect 21331 21496 21392 21530
rect 21438 21518 21482 21530
rect 21538 21518 21572 21530
rect 21638 21518 21662 21530
rect 21426 21496 21482 21518
rect 21516 21496 21572 21518
rect 21606 21496 21662 21518
rect 21696 21518 21704 21530
rect 21738 21530 21804 21552
rect 21738 21518 21752 21530
rect 21696 21496 21752 21518
rect 21786 21518 21804 21530
rect 21838 21530 21904 21552
rect 21938 21530 22025 21552
rect 21838 21518 21842 21530
rect 21786 21496 21842 21518
rect 21876 21518 21904 21530
rect 21876 21496 21932 21518
rect 21966 21496 22025 21530
rect 21331 21452 22025 21496
rect 21331 21440 21404 21452
rect 21438 21440 21504 21452
rect 21538 21440 21604 21452
rect 21638 21440 21704 21452
rect 21331 21406 21392 21440
rect 21438 21418 21482 21440
rect 21538 21418 21572 21440
rect 21638 21418 21662 21440
rect 21426 21406 21482 21418
rect 21516 21406 21572 21418
rect 21606 21406 21662 21418
rect 21696 21418 21704 21440
rect 21738 21440 21804 21452
rect 21738 21418 21752 21440
rect 21696 21406 21752 21418
rect 21786 21418 21804 21440
rect 21838 21440 21904 21452
rect 21938 21440 22025 21452
rect 21838 21418 21842 21440
rect 21786 21406 21842 21418
rect 21876 21418 21904 21440
rect 21876 21406 21932 21418
rect 21966 21406 22025 21440
rect 21331 21345 22025 21406
rect 22087 21988 22159 22044
rect 22087 21954 22106 21988
rect 22140 21954 22159 21988
rect 22087 21898 22159 21954
rect 22087 21864 22106 21898
rect 22140 21864 22159 21898
rect 22087 21808 22159 21864
rect 22087 21774 22106 21808
rect 22140 21774 22159 21808
rect 22087 21718 22159 21774
rect 22087 21684 22106 21718
rect 22140 21684 22159 21718
rect 22087 21628 22159 21684
rect 22087 21594 22106 21628
rect 22140 21594 22159 21628
rect 22087 21538 22159 21594
rect 22087 21504 22106 21538
rect 22140 21504 22159 21538
rect 22087 21448 22159 21504
rect 22087 21414 22106 21448
rect 22140 21414 22159 21448
rect 22087 21358 22159 21414
rect 21197 21283 21269 21343
rect 22087 21324 22106 21358
rect 22140 21324 22159 21358
rect 22087 21283 22159 21324
rect 21197 21267 22159 21283
rect 21034 21198 21133 21254
rect 21223 21264 22159 21267
rect 21223 21233 21294 21264
rect 21197 21230 21294 21233
rect 21328 21230 21384 21264
rect 21418 21230 21474 21264
rect 21508 21230 21564 21264
rect 21598 21230 21654 21264
rect 21688 21230 21744 21264
rect 21778 21230 21834 21264
rect 21868 21230 21924 21264
rect 21958 21230 22014 21264
rect 22048 21230 22159 21264
rect 21197 21211 22159 21230
rect 22223 22154 22255 22188
rect 22289 22154 22322 22188
rect 23437 22156 23471 22442
rect 24353 22156 24387 22442
rect 25269 22156 25303 22442
rect 26185 22156 26219 22442
rect 27101 22156 27135 22442
rect 28286 22316 38954 22336
rect 28286 22282 28306 22316
rect 28340 22282 28396 22316
rect 28430 22301 28486 22316
rect 28520 22301 28576 22316
rect 28610 22301 28666 22316
rect 28700 22301 28756 22316
rect 28790 22301 28846 22316
rect 28880 22301 28936 22316
rect 28970 22301 29026 22316
rect 29060 22301 29116 22316
rect 29150 22301 29206 22316
rect 29240 22301 29296 22316
rect 29330 22301 29386 22316
rect 29420 22301 29476 22316
rect 28450 22282 28486 22301
rect 28540 22282 28576 22301
rect 28630 22282 28666 22301
rect 28720 22282 28756 22301
rect 28810 22282 28846 22301
rect 28900 22282 28936 22301
rect 28990 22282 29026 22301
rect 29080 22282 29116 22301
rect 29170 22282 29206 22301
rect 29260 22282 29296 22301
rect 29350 22282 29386 22301
rect 29440 22282 29476 22301
rect 29510 22282 29646 22316
rect 29680 22282 29736 22316
rect 29770 22301 29826 22316
rect 29860 22301 29916 22316
rect 29950 22301 30006 22316
rect 30040 22301 30096 22316
rect 30130 22301 30186 22316
rect 30220 22301 30276 22316
rect 30310 22301 30366 22316
rect 30400 22301 30456 22316
rect 30490 22301 30546 22316
rect 30580 22301 30636 22316
rect 30670 22301 30726 22316
rect 30760 22301 30816 22316
rect 29790 22282 29826 22301
rect 29880 22282 29916 22301
rect 29970 22282 30006 22301
rect 30060 22282 30096 22301
rect 30150 22282 30186 22301
rect 30240 22282 30276 22301
rect 30330 22282 30366 22301
rect 30420 22282 30456 22301
rect 30510 22282 30546 22301
rect 30600 22282 30636 22301
rect 30690 22282 30726 22301
rect 30780 22282 30816 22301
rect 30850 22282 30986 22316
rect 31020 22282 31076 22316
rect 31110 22301 31166 22316
rect 31200 22301 31256 22316
rect 31290 22301 31346 22316
rect 31380 22301 31436 22316
rect 31470 22301 31526 22316
rect 31560 22301 31616 22316
rect 31650 22301 31706 22316
rect 31740 22301 31796 22316
rect 31830 22301 31886 22316
rect 31920 22301 31976 22316
rect 32010 22301 32066 22316
rect 32100 22301 32156 22316
rect 31130 22282 31166 22301
rect 31220 22282 31256 22301
rect 31310 22282 31346 22301
rect 31400 22282 31436 22301
rect 31490 22282 31526 22301
rect 31580 22282 31616 22301
rect 31670 22282 31706 22301
rect 31760 22282 31796 22301
rect 31850 22282 31886 22301
rect 31940 22282 31976 22301
rect 32030 22282 32066 22301
rect 32120 22282 32156 22301
rect 32190 22282 32326 22316
rect 32360 22282 32416 22316
rect 32450 22301 32506 22316
rect 32540 22301 32596 22316
rect 32630 22301 32686 22316
rect 32720 22301 32776 22316
rect 32810 22301 32866 22316
rect 32900 22301 32956 22316
rect 32990 22301 33046 22316
rect 33080 22301 33136 22316
rect 33170 22301 33226 22316
rect 33260 22301 33316 22316
rect 33350 22301 33406 22316
rect 33440 22301 33496 22316
rect 32470 22282 32506 22301
rect 32560 22282 32596 22301
rect 32650 22282 32686 22301
rect 32740 22282 32776 22301
rect 32830 22282 32866 22301
rect 32920 22282 32956 22301
rect 33010 22282 33046 22301
rect 33100 22282 33136 22301
rect 33190 22282 33226 22301
rect 33280 22282 33316 22301
rect 33370 22282 33406 22301
rect 33460 22282 33496 22301
rect 33530 22282 33666 22316
rect 33700 22282 33756 22316
rect 33790 22301 33846 22316
rect 33880 22301 33936 22316
rect 33970 22301 34026 22316
rect 34060 22301 34116 22316
rect 34150 22301 34206 22316
rect 34240 22301 34296 22316
rect 34330 22301 34386 22316
rect 34420 22301 34476 22316
rect 34510 22301 34566 22316
rect 34600 22301 34656 22316
rect 34690 22301 34746 22316
rect 34780 22301 34836 22316
rect 33810 22282 33846 22301
rect 33900 22282 33936 22301
rect 33990 22282 34026 22301
rect 34080 22282 34116 22301
rect 34170 22282 34206 22301
rect 34260 22282 34296 22301
rect 34350 22282 34386 22301
rect 34440 22282 34476 22301
rect 34530 22282 34566 22301
rect 34620 22282 34656 22301
rect 34710 22282 34746 22301
rect 34800 22282 34836 22301
rect 34870 22282 35006 22316
rect 35040 22282 35096 22316
rect 35130 22301 35186 22316
rect 35220 22301 35276 22316
rect 35310 22301 35366 22316
rect 35400 22301 35456 22316
rect 35490 22301 35546 22316
rect 35580 22301 35636 22316
rect 35670 22301 35726 22316
rect 35760 22301 35816 22316
rect 35850 22301 35906 22316
rect 35940 22301 35996 22316
rect 36030 22301 36086 22316
rect 36120 22301 36176 22316
rect 35150 22282 35186 22301
rect 35240 22282 35276 22301
rect 35330 22282 35366 22301
rect 35420 22282 35456 22301
rect 35510 22282 35546 22301
rect 35600 22282 35636 22301
rect 35690 22282 35726 22301
rect 35780 22282 35816 22301
rect 35870 22282 35906 22301
rect 35960 22282 35996 22301
rect 36050 22282 36086 22301
rect 36140 22282 36176 22301
rect 36210 22282 36346 22316
rect 36380 22282 36436 22316
rect 36470 22301 36526 22316
rect 36560 22301 36616 22316
rect 36650 22301 36706 22316
rect 36740 22301 36796 22316
rect 36830 22301 36886 22316
rect 36920 22301 36976 22316
rect 37010 22301 37066 22316
rect 37100 22301 37156 22316
rect 37190 22301 37246 22316
rect 37280 22301 37336 22316
rect 37370 22301 37426 22316
rect 37460 22301 37516 22316
rect 36490 22282 36526 22301
rect 36580 22282 36616 22301
rect 36670 22282 36706 22301
rect 36760 22282 36796 22301
rect 36850 22282 36886 22301
rect 36940 22282 36976 22301
rect 37030 22282 37066 22301
rect 37120 22282 37156 22301
rect 37210 22282 37246 22301
rect 37300 22282 37336 22301
rect 37390 22282 37426 22301
rect 37480 22282 37516 22301
rect 37550 22282 37686 22316
rect 37720 22282 37776 22316
rect 37810 22301 37866 22316
rect 37900 22301 37956 22316
rect 37990 22301 38046 22316
rect 38080 22301 38136 22316
rect 38170 22301 38226 22316
rect 38260 22301 38316 22316
rect 38350 22301 38406 22316
rect 38440 22301 38496 22316
rect 38530 22301 38586 22316
rect 38620 22301 38676 22316
rect 38710 22301 38766 22316
rect 38800 22301 38856 22316
rect 37830 22282 37866 22301
rect 37920 22282 37956 22301
rect 38010 22282 38046 22301
rect 38100 22282 38136 22301
rect 38190 22282 38226 22301
rect 38280 22282 38316 22301
rect 38370 22282 38406 22301
rect 38460 22282 38496 22301
rect 38550 22282 38586 22301
rect 38640 22282 38676 22301
rect 38730 22282 38766 22301
rect 38820 22282 38856 22301
rect 38890 22282 38954 22316
rect 28286 22278 28416 22282
rect 28286 22244 28320 22278
rect 28354 22267 28416 22278
rect 28450 22267 28506 22282
rect 28540 22267 28596 22282
rect 28630 22267 28686 22282
rect 28720 22267 28776 22282
rect 28810 22267 28866 22282
rect 28900 22267 28956 22282
rect 28990 22267 29046 22282
rect 29080 22267 29136 22282
rect 29170 22267 29226 22282
rect 29260 22267 29316 22282
rect 29350 22267 29406 22282
rect 29440 22278 29756 22282
rect 29440 22267 29507 22278
rect 28354 22244 29507 22267
rect 29541 22244 29660 22278
rect 29694 22267 29756 22278
rect 29790 22267 29846 22282
rect 29880 22267 29936 22282
rect 29970 22267 30026 22282
rect 30060 22267 30116 22282
rect 30150 22267 30206 22282
rect 30240 22267 30296 22282
rect 30330 22267 30386 22282
rect 30420 22267 30476 22282
rect 30510 22267 30566 22282
rect 30600 22267 30656 22282
rect 30690 22267 30746 22282
rect 30780 22278 31096 22282
rect 30780 22267 30847 22278
rect 29694 22244 30847 22267
rect 30881 22244 31000 22278
rect 31034 22267 31096 22278
rect 31130 22267 31186 22282
rect 31220 22267 31276 22282
rect 31310 22267 31366 22282
rect 31400 22267 31456 22282
rect 31490 22267 31546 22282
rect 31580 22267 31636 22282
rect 31670 22267 31726 22282
rect 31760 22267 31816 22282
rect 31850 22267 31906 22282
rect 31940 22267 31996 22282
rect 32030 22267 32086 22282
rect 32120 22278 32436 22282
rect 32120 22267 32187 22278
rect 31034 22244 32187 22267
rect 32221 22244 32340 22278
rect 32374 22267 32436 22278
rect 32470 22267 32526 22282
rect 32560 22267 32616 22282
rect 32650 22267 32706 22282
rect 32740 22267 32796 22282
rect 32830 22267 32886 22282
rect 32920 22267 32976 22282
rect 33010 22267 33066 22282
rect 33100 22267 33156 22282
rect 33190 22267 33246 22282
rect 33280 22267 33336 22282
rect 33370 22267 33426 22282
rect 33460 22278 33776 22282
rect 33460 22267 33527 22278
rect 32374 22244 33527 22267
rect 33561 22244 33680 22278
rect 33714 22267 33776 22278
rect 33810 22267 33866 22282
rect 33900 22267 33956 22282
rect 33990 22267 34046 22282
rect 34080 22267 34136 22282
rect 34170 22267 34226 22282
rect 34260 22267 34316 22282
rect 34350 22267 34406 22282
rect 34440 22267 34496 22282
rect 34530 22267 34586 22282
rect 34620 22267 34676 22282
rect 34710 22267 34766 22282
rect 34800 22278 35116 22282
rect 34800 22267 34867 22278
rect 33714 22244 34867 22267
rect 34901 22244 35020 22278
rect 35054 22267 35116 22278
rect 35150 22267 35206 22282
rect 35240 22267 35296 22282
rect 35330 22267 35386 22282
rect 35420 22267 35476 22282
rect 35510 22267 35566 22282
rect 35600 22267 35656 22282
rect 35690 22267 35746 22282
rect 35780 22267 35836 22282
rect 35870 22267 35926 22282
rect 35960 22267 36016 22282
rect 36050 22267 36106 22282
rect 36140 22278 36456 22282
rect 36140 22267 36207 22278
rect 35054 22244 36207 22267
rect 36241 22244 36360 22278
rect 36394 22267 36456 22278
rect 36490 22267 36546 22282
rect 36580 22267 36636 22282
rect 36670 22267 36726 22282
rect 36760 22267 36816 22282
rect 36850 22267 36906 22282
rect 36940 22267 36996 22282
rect 37030 22267 37086 22282
rect 37120 22267 37176 22282
rect 37210 22267 37266 22282
rect 37300 22267 37356 22282
rect 37390 22267 37446 22282
rect 37480 22278 37796 22282
rect 37480 22267 37547 22278
rect 36394 22244 37547 22267
rect 37581 22244 37700 22278
rect 37734 22267 37796 22278
rect 37830 22267 37886 22282
rect 37920 22267 37976 22282
rect 38010 22267 38066 22282
rect 38100 22267 38156 22282
rect 38190 22267 38246 22282
rect 38280 22267 38336 22282
rect 38370 22267 38426 22282
rect 38460 22267 38516 22282
rect 38550 22267 38606 22282
rect 38640 22267 38696 22282
rect 38730 22267 38786 22282
rect 38820 22278 38954 22282
rect 38820 22267 38887 22278
rect 37734 22244 38887 22267
rect 38921 22244 38954 22278
rect 28286 22237 38954 22244
rect 28286 22188 28385 22237
rect 22223 22098 22322 22154
rect 22223 22064 22255 22098
rect 22289 22064 22322 22098
rect 22223 22008 22322 22064
rect 22223 21974 22255 22008
rect 22289 21974 22322 22008
rect 22223 21918 22322 21974
rect 22223 21884 22255 21918
rect 22289 21884 22322 21918
rect 22223 21828 22322 21884
rect 22223 21794 22255 21828
rect 22289 21794 22322 21828
rect 22223 21738 22322 21794
rect 22223 21704 22255 21738
rect 22289 21704 22322 21738
rect 22223 21648 22322 21704
rect 22223 21614 22255 21648
rect 22289 21614 22322 21648
rect 22223 21558 22322 21614
rect 22223 21524 22255 21558
rect 22289 21524 22322 21558
rect 22223 21468 22322 21524
rect 22223 21434 22255 21468
rect 22289 21434 22322 21468
rect 22223 21378 22322 21434
rect 22980 22129 23014 22156
rect 23437 22138 23472 22156
rect 22980 22057 23014 22075
rect 22980 21985 23014 22007
rect 22980 21913 23014 21939
rect 22980 21841 23014 21871
rect 22980 21769 23014 21803
rect 22980 21701 23014 21735
rect 22980 21633 23014 21663
rect 22980 21565 23014 21591
rect 22980 21497 23014 21519
rect 22980 21429 23014 21447
rect 22223 21344 22255 21378
rect 22289 21344 22322 21378
rect 22223 21288 22322 21344
rect 22223 21254 22255 21288
rect 22289 21254 22322 21288
rect 22979 21375 22980 21406
rect 22979 21348 23014 21375
rect 23438 22129 23472 22138
rect 23438 22057 23472 22075
rect 23438 21985 23472 22007
rect 23438 21913 23472 21939
rect 23438 21841 23472 21871
rect 23438 21769 23472 21803
rect 23438 21701 23472 21735
rect 23438 21633 23472 21663
rect 23438 21565 23472 21591
rect 23438 21497 23472 21519
rect 23438 21429 23472 21447
rect 23896 22129 23930 22156
rect 24353 22138 24388 22156
rect 23896 22057 23930 22075
rect 23896 21985 23930 22007
rect 23896 21913 23930 21939
rect 23896 21841 23930 21871
rect 23896 21769 23930 21803
rect 23896 21701 23930 21735
rect 23896 21633 23930 21663
rect 23896 21565 23930 21591
rect 23896 21497 23930 21519
rect 23896 21429 23930 21447
rect 23438 21348 23472 21375
rect 23895 21375 23896 21406
rect 23895 21348 23930 21375
rect 24354 22129 24388 22138
rect 24354 22057 24388 22075
rect 24354 21985 24388 22007
rect 24354 21913 24388 21939
rect 24354 21841 24388 21871
rect 24354 21769 24388 21803
rect 24354 21701 24388 21735
rect 24354 21633 24388 21663
rect 24354 21565 24388 21591
rect 24354 21497 24388 21519
rect 24354 21429 24388 21447
rect 24812 22129 24846 22156
rect 25269 22138 25304 22156
rect 24812 22057 24846 22075
rect 24812 21985 24846 22007
rect 24812 21913 24846 21939
rect 24812 21841 24846 21871
rect 24812 21769 24846 21803
rect 24812 21701 24846 21735
rect 24812 21633 24846 21663
rect 24812 21565 24846 21591
rect 24812 21497 24846 21519
rect 24812 21429 24846 21447
rect 24354 21348 24388 21375
rect 24811 21375 24812 21406
rect 24811 21348 24846 21375
rect 25270 22129 25304 22138
rect 25270 22057 25304 22075
rect 25270 21985 25304 22007
rect 25270 21913 25304 21939
rect 25270 21841 25304 21871
rect 25270 21769 25304 21803
rect 25270 21701 25304 21735
rect 25270 21633 25304 21663
rect 25270 21565 25304 21591
rect 25270 21497 25304 21519
rect 25270 21429 25304 21447
rect 25728 22129 25762 22156
rect 26185 22138 26220 22156
rect 25728 22057 25762 22075
rect 25728 21985 25762 22007
rect 25728 21913 25762 21939
rect 25728 21841 25762 21871
rect 25728 21769 25762 21803
rect 25728 21701 25762 21735
rect 25728 21633 25762 21663
rect 25728 21565 25762 21591
rect 25728 21497 25762 21519
rect 25728 21429 25762 21447
rect 25270 21348 25304 21375
rect 25727 21375 25728 21406
rect 25727 21348 25762 21375
rect 26186 22129 26220 22138
rect 26186 22057 26220 22075
rect 26186 21985 26220 22007
rect 26186 21913 26220 21939
rect 26186 21841 26220 21871
rect 26186 21769 26220 21803
rect 26186 21701 26220 21735
rect 26186 21633 26220 21663
rect 26186 21565 26220 21591
rect 26186 21497 26220 21519
rect 26186 21429 26220 21447
rect 26644 22129 26678 22156
rect 27101 22138 27136 22156
rect 26644 22057 26678 22075
rect 26644 21985 26678 22007
rect 26644 21913 26678 21939
rect 26644 21841 26678 21871
rect 26644 21769 26678 21803
rect 26644 21701 26678 21735
rect 26644 21633 26678 21663
rect 26644 21565 26678 21591
rect 26644 21497 26678 21519
rect 26644 21429 26678 21447
rect 26186 21348 26220 21375
rect 26643 21375 26644 21406
rect 26643 21348 26678 21375
rect 27102 22129 27136 22138
rect 27102 22057 27136 22075
rect 27102 21985 27136 22007
rect 27102 21913 27136 21939
rect 27102 21841 27136 21871
rect 27102 21769 27136 21803
rect 27102 21701 27136 21735
rect 27102 21633 27136 21663
rect 27102 21565 27136 21591
rect 27102 21497 27136 21519
rect 27102 21429 27136 21447
rect 27102 21348 27136 21375
rect 28286 22154 28320 22188
rect 28354 22154 28385 22188
rect 29475 22188 29725 22237
rect 28286 22098 28385 22154
rect 28286 22064 28320 22098
rect 28354 22064 28385 22098
rect 28286 22008 28385 22064
rect 28286 21974 28320 22008
rect 28354 21974 28385 22008
rect 28286 21918 28385 21974
rect 28286 21884 28320 21918
rect 28354 21884 28385 21918
rect 28286 21828 28385 21884
rect 28286 21794 28320 21828
rect 28354 21794 28385 21828
rect 28286 21738 28385 21794
rect 28286 21704 28320 21738
rect 28354 21704 28385 21738
rect 28286 21648 28385 21704
rect 28286 21614 28320 21648
rect 28354 21614 28385 21648
rect 28286 21558 28385 21614
rect 28286 21524 28320 21558
rect 28354 21524 28385 21558
rect 28286 21468 28385 21524
rect 28286 21434 28320 21468
rect 28354 21434 28385 21468
rect 28286 21378 28385 21434
rect 22979 21282 23013 21348
rect 23895 21282 23929 21348
rect 24811 21282 24845 21348
rect 25727 21282 25761 21348
rect 26643 21282 26677 21348
rect 28286 21344 28320 21378
rect 28354 21344 28385 21378
rect 28286 21288 28385 21344
rect 21034 21164 21068 21198
rect 21102 21164 21133 21198
rect 21034 21147 21133 21164
rect 22223 21198 22322 21254
rect 22968 21267 27148 21282
rect 22968 21233 26525 21267
rect 26559 21233 27148 21267
rect 22968 21222 27148 21233
rect 28286 21254 28320 21288
rect 28354 21254 28385 21288
rect 22223 21164 22255 21198
rect 22289 21164 22322 21198
rect 22223 21147 22322 21164
rect 21034 21131 22322 21147
rect 28286 21198 28385 21254
rect 28449 22156 29411 22173
rect 28449 22122 28470 22156
rect 28504 22122 28560 22156
rect 28594 22154 28650 22156
rect 28684 22154 28740 22156
rect 28774 22154 28830 22156
rect 28864 22154 28920 22156
rect 28954 22154 29010 22156
rect 29044 22154 29100 22156
rect 29134 22154 29190 22156
rect 29224 22154 29280 22156
rect 29314 22154 29370 22156
rect 28614 22122 28650 22154
rect 28704 22122 28740 22154
rect 28794 22122 28830 22154
rect 28884 22122 28920 22154
rect 28974 22122 29010 22154
rect 29064 22122 29100 22154
rect 29154 22122 29190 22154
rect 29244 22122 29280 22154
rect 29334 22122 29370 22154
rect 29404 22122 29411 22156
rect 28449 22120 28580 22122
rect 28614 22120 28670 22122
rect 28704 22120 28760 22122
rect 28794 22120 28850 22122
rect 28884 22120 28940 22122
rect 28974 22120 29030 22122
rect 29064 22120 29120 22122
rect 29154 22120 29210 22122
rect 29244 22120 29300 22122
rect 29334 22120 29411 22122
rect 28449 22101 29411 22120
rect 28449 22097 28521 22101
rect 28449 22063 28468 22097
rect 28502 22063 28521 22097
rect 28449 22007 28521 22063
rect 29339 22078 29411 22101
rect 29339 22044 29358 22078
rect 29392 22044 29411 22078
rect 28449 21973 28468 22007
rect 28502 21973 28521 22007
rect 28449 21917 28521 21973
rect 28449 21883 28468 21917
rect 28502 21883 28521 21917
rect 28449 21827 28521 21883
rect 28449 21793 28468 21827
rect 28502 21793 28521 21827
rect 28449 21737 28521 21793
rect 28449 21703 28468 21737
rect 28502 21703 28521 21737
rect 28449 21647 28521 21703
rect 28449 21613 28468 21647
rect 28502 21613 28521 21647
rect 28449 21557 28521 21613
rect 28449 21523 28468 21557
rect 28502 21523 28521 21557
rect 28449 21467 28521 21523
rect 28449 21433 28468 21467
rect 28502 21433 28521 21467
rect 28449 21377 28521 21433
rect 28449 21343 28468 21377
rect 28502 21343 28521 21377
rect 28583 21980 29277 22039
rect 28583 21946 28644 21980
rect 28678 21952 28734 21980
rect 28768 21952 28824 21980
rect 28858 21952 28914 21980
rect 28690 21946 28734 21952
rect 28790 21946 28824 21952
rect 28890 21946 28914 21952
rect 28948 21952 29004 21980
rect 28948 21946 28956 21952
rect 28583 21918 28656 21946
rect 28690 21918 28756 21946
rect 28790 21918 28856 21946
rect 28890 21918 28956 21946
rect 28990 21946 29004 21952
rect 29038 21952 29094 21980
rect 29038 21946 29056 21952
rect 28990 21918 29056 21946
rect 29090 21946 29094 21952
rect 29128 21952 29184 21980
rect 29128 21946 29156 21952
rect 29218 21946 29277 21980
rect 29090 21918 29156 21946
rect 29190 21918 29277 21946
rect 28583 21890 29277 21918
rect 28583 21856 28644 21890
rect 28678 21856 28734 21890
rect 28768 21856 28824 21890
rect 28858 21856 28914 21890
rect 28948 21856 29004 21890
rect 29038 21856 29094 21890
rect 29128 21856 29184 21890
rect 29218 21856 29277 21890
rect 28583 21852 29277 21856
rect 28583 21818 28656 21852
rect 28690 21818 28756 21852
rect 28790 21818 28856 21852
rect 28890 21818 28956 21852
rect 28990 21818 29056 21852
rect 29090 21818 29156 21852
rect 29190 21818 29277 21852
rect 28583 21800 29277 21818
rect 28583 21766 28644 21800
rect 28678 21766 28734 21800
rect 28768 21766 28824 21800
rect 28858 21766 28914 21800
rect 28948 21766 29004 21800
rect 29038 21766 29094 21800
rect 29128 21766 29184 21800
rect 29218 21766 29277 21800
rect 28583 21752 29277 21766
rect 28583 21718 28656 21752
rect 28690 21718 28756 21752
rect 28790 21718 28856 21752
rect 28890 21718 28956 21752
rect 28990 21718 29056 21752
rect 29090 21718 29156 21752
rect 29190 21718 29277 21752
rect 28583 21710 29277 21718
rect 28583 21676 28644 21710
rect 28678 21676 28734 21710
rect 28768 21676 28824 21710
rect 28858 21676 28914 21710
rect 28948 21676 29004 21710
rect 29038 21676 29094 21710
rect 29128 21676 29184 21710
rect 29218 21676 29277 21710
rect 28583 21652 29277 21676
rect 28583 21620 28656 21652
rect 28690 21620 28756 21652
rect 28790 21620 28856 21652
rect 28890 21620 28956 21652
rect 28583 21586 28644 21620
rect 28690 21618 28734 21620
rect 28790 21618 28824 21620
rect 28890 21618 28914 21620
rect 28678 21586 28734 21618
rect 28768 21586 28824 21618
rect 28858 21586 28914 21618
rect 28948 21618 28956 21620
rect 28990 21620 29056 21652
rect 28990 21618 29004 21620
rect 28948 21586 29004 21618
rect 29038 21618 29056 21620
rect 29090 21620 29156 21652
rect 29190 21620 29277 21652
rect 29090 21618 29094 21620
rect 29038 21586 29094 21618
rect 29128 21618 29156 21620
rect 29128 21586 29184 21618
rect 29218 21586 29277 21620
rect 28583 21552 29277 21586
rect 28583 21530 28656 21552
rect 28690 21530 28756 21552
rect 28790 21530 28856 21552
rect 28890 21530 28956 21552
rect 28583 21496 28644 21530
rect 28690 21518 28734 21530
rect 28790 21518 28824 21530
rect 28890 21518 28914 21530
rect 28678 21496 28734 21518
rect 28768 21496 28824 21518
rect 28858 21496 28914 21518
rect 28948 21518 28956 21530
rect 28990 21530 29056 21552
rect 28990 21518 29004 21530
rect 28948 21496 29004 21518
rect 29038 21518 29056 21530
rect 29090 21530 29156 21552
rect 29190 21530 29277 21552
rect 29090 21518 29094 21530
rect 29038 21496 29094 21518
rect 29128 21518 29156 21530
rect 29128 21496 29184 21518
rect 29218 21496 29277 21530
rect 28583 21452 29277 21496
rect 28583 21440 28656 21452
rect 28690 21440 28756 21452
rect 28790 21440 28856 21452
rect 28890 21440 28956 21452
rect 28583 21406 28644 21440
rect 28690 21418 28734 21440
rect 28790 21418 28824 21440
rect 28890 21418 28914 21440
rect 28678 21406 28734 21418
rect 28768 21406 28824 21418
rect 28858 21406 28914 21418
rect 28948 21418 28956 21440
rect 28990 21440 29056 21452
rect 28990 21418 29004 21440
rect 28948 21406 29004 21418
rect 29038 21418 29056 21440
rect 29090 21440 29156 21452
rect 29190 21440 29277 21452
rect 29090 21418 29094 21440
rect 29038 21406 29094 21418
rect 29128 21418 29156 21440
rect 29128 21406 29184 21418
rect 29218 21406 29277 21440
rect 28583 21345 29277 21406
rect 29339 21988 29411 22044
rect 29339 21954 29358 21988
rect 29392 21954 29411 21988
rect 29339 21898 29411 21954
rect 29339 21864 29358 21898
rect 29392 21864 29411 21898
rect 29339 21808 29411 21864
rect 29339 21774 29358 21808
rect 29392 21774 29411 21808
rect 29339 21718 29411 21774
rect 29339 21684 29358 21718
rect 29392 21684 29411 21718
rect 29339 21628 29411 21684
rect 29339 21594 29358 21628
rect 29392 21594 29411 21628
rect 29339 21538 29411 21594
rect 29339 21504 29358 21538
rect 29392 21504 29411 21538
rect 29339 21448 29411 21504
rect 29339 21414 29358 21448
rect 29392 21414 29411 21448
rect 29339 21358 29411 21414
rect 28449 21283 28521 21343
rect 29339 21324 29358 21358
rect 29392 21324 29411 21358
rect 29339 21283 29411 21324
rect 28449 21264 29411 21283
rect 28449 21230 28546 21264
rect 28580 21230 28636 21264
rect 28670 21230 28726 21264
rect 28760 21230 28816 21264
rect 28850 21230 28906 21264
rect 28940 21230 28996 21264
rect 29030 21230 29086 21264
rect 29120 21230 29176 21264
rect 29210 21230 29266 21264
rect 29300 21230 29411 21264
rect 28449 21211 29411 21230
rect 29475 22154 29507 22188
rect 29541 22154 29660 22188
rect 29694 22154 29725 22188
rect 30815 22188 31065 22237
rect 29475 22098 29725 22154
rect 29475 22064 29507 22098
rect 29541 22064 29660 22098
rect 29694 22064 29725 22098
rect 29475 22008 29725 22064
rect 29475 21974 29507 22008
rect 29541 21974 29660 22008
rect 29694 21974 29725 22008
rect 29475 21918 29725 21974
rect 29475 21884 29507 21918
rect 29541 21884 29660 21918
rect 29694 21884 29725 21918
rect 29475 21828 29725 21884
rect 29475 21794 29507 21828
rect 29541 21794 29660 21828
rect 29694 21794 29725 21828
rect 29475 21738 29725 21794
rect 29475 21704 29507 21738
rect 29541 21704 29660 21738
rect 29694 21704 29725 21738
rect 29475 21648 29725 21704
rect 29475 21614 29507 21648
rect 29541 21614 29660 21648
rect 29694 21614 29725 21648
rect 29475 21558 29725 21614
rect 29475 21524 29507 21558
rect 29541 21524 29660 21558
rect 29694 21524 29725 21558
rect 29475 21468 29725 21524
rect 29475 21434 29507 21468
rect 29541 21434 29660 21468
rect 29694 21434 29725 21468
rect 29475 21378 29725 21434
rect 29475 21344 29507 21378
rect 29541 21344 29660 21378
rect 29694 21344 29725 21378
rect 29475 21288 29725 21344
rect 29475 21254 29507 21288
rect 29541 21254 29660 21288
rect 29694 21254 29725 21288
rect 28286 21164 28320 21198
rect 28354 21164 28385 21198
rect 28286 21147 28385 21164
rect 29475 21198 29725 21254
rect 29789 22156 30751 22173
rect 29789 22122 29810 22156
rect 29844 22122 29900 22156
rect 29934 22154 29990 22156
rect 30024 22154 30080 22156
rect 30114 22154 30170 22156
rect 30204 22154 30260 22156
rect 30294 22154 30350 22156
rect 30384 22154 30440 22156
rect 30474 22154 30530 22156
rect 30564 22154 30620 22156
rect 30654 22154 30710 22156
rect 29954 22122 29990 22154
rect 30044 22122 30080 22154
rect 30134 22122 30170 22154
rect 30224 22122 30260 22154
rect 30314 22122 30350 22154
rect 30404 22122 30440 22154
rect 30494 22122 30530 22154
rect 30584 22122 30620 22154
rect 30674 22122 30710 22154
rect 30744 22122 30751 22156
rect 29789 22120 29920 22122
rect 29954 22120 30010 22122
rect 30044 22120 30100 22122
rect 30134 22120 30190 22122
rect 30224 22120 30280 22122
rect 30314 22120 30370 22122
rect 30404 22120 30460 22122
rect 30494 22120 30550 22122
rect 30584 22120 30640 22122
rect 30674 22120 30751 22122
rect 29789 22101 30751 22120
rect 29789 22097 29861 22101
rect 29789 22063 29808 22097
rect 29842 22063 29861 22097
rect 29789 22007 29861 22063
rect 30679 22078 30751 22101
rect 30679 22044 30698 22078
rect 30732 22044 30751 22078
rect 29789 21973 29808 22007
rect 29842 21973 29861 22007
rect 29789 21917 29861 21973
rect 29789 21883 29808 21917
rect 29842 21883 29861 21917
rect 29789 21827 29861 21883
rect 29789 21793 29808 21827
rect 29842 21793 29861 21827
rect 29789 21737 29861 21793
rect 29789 21703 29808 21737
rect 29842 21703 29861 21737
rect 29789 21647 29861 21703
rect 29789 21613 29808 21647
rect 29842 21613 29861 21647
rect 29789 21557 29861 21613
rect 29789 21523 29808 21557
rect 29842 21523 29861 21557
rect 29789 21467 29861 21523
rect 29789 21433 29808 21467
rect 29842 21433 29861 21467
rect 29789 21377 29861 21433
rect 29789 21343 29808 21377
rect 29842 21343 29861 21377
rect 29923 21980 30617 22039
rect 29923 21946 29984 21980
rect 30018 21952 30074 21980
rect 30108 21952 30164 21980
rect 30198 21952 30254 21980
rect 30030 21946 30074 21952
rect 30130 21946 30164 21952
rect 30230 21946 30254 21952
rect 30288 21952 30344 21980
rect 30288 21946 30296 21952
rect 29923 21918 29996 21946
rect 30030 21918 30096 21946
rect 30130 21918 30196 21946
rect 30230 21918 30296 21946
rect 30330 21946 30344 21952
rect 30378 21952 30434 21980
rect 30378 21946 30396 21952
rect 30330 21918 30396 21946
rect 30430 21946 30434 21952
rect 30468 21952 30524 21980
rect 30468 21946 30496 21952
rect 30558 21946 30617 21980
rect 30430 21918 30496 21946
rect 30530 21918 30617 21946
rect 29923 21890 30617 21918
rect 29923 21856 29984 21890
rect 30018 21856 30074 21890
rect 30108 21856 30164 21890
rect 30198 21856 30254 21890
rect 30288 21856 30344 21890
rect 30378 21856 30434 21890
rect 30468 21856 30524 21890
rect 30558 21856 30617 21890
rect 29923 21852 30617 21856
rect 29923 21818 29996 21852
rect 30030 21818 30096 21852
rect 30130 21818 30196 21852
rect 30230 21818 30296 21852
rect 30330 21818 30396 21852
rect 30430 21818 30496 21852
rect 30530 21818 30617 21852
rect 29923 21800 30617 21818
rect 29923 21766 29984 21800
rect 30018 21766 30074 21800
rect 30108 21766 30164 21800
rect 30198 21766 30254 21800
rect 30288 21766 30344 21800
rect 30378 21766 30434 21800
rect 30468 21766 30524 21800
rect 30558 21766 30617 21800
rect 29923 21752 30617 21766
rect 29923 21718 29996 21752
rect 30030 21718 30096 21752
rect 30130 21718 30196 21752
rect 30230 21718 30296 21752
rect 30330 21718 30396 21752
rect 30430 21718 30496 21752
rect 30530 21718 30617 21752
rect 29923 21710 30617 21718
rect 29923 21676 29984 21710
rect 30018 21676 30074 21710
rect 30108 21676 30164 21710
rect 30198 21676 30254 21710
rect 30288 21676 30344 21710
rect 30378 21676 30434 21710
rect 30468 21676 30524 21710
rect 30558 21676 30617 21710
rect 29923 21652 30617 21676
rect 29923 21620 29996 21652
rect 30030 21620 30096 21652
rect 30130 21620 30196 21652
rect 30230 21620 30296 21652
rect 29923 21586 29984 21620
rect 30030 21618 30074 21620
rect 30130 21618 30164 21620
rect 30230 21618 30254 21620
rect 30018 21586 30074 21618
rect 30108 21586 30164 21618
rect 30198 21586 30254 21618
rect 30288 21618 30296 21620
rect 30330 21620 30396 21652
rect 30330 21618 30344 21620
rect 30288 21586 30344 21618
rect 30378 21618 30396 21620
rect 30430 21620 30496 21652
rect 30530 21620 30617 21652
rect 30430 21618 30434 21620
rect 30378 21586 30434 21618
rect 30468 21618 30496 21620
rect 30468 21586 30524 21618
rect 30558 21586 30617 21620
rect 29923 21552 30617 21586
rect 29923 21530 29996 21552
rect 30030 21530 30096 21552
rect 30130 21530 30196 21552
rect 30230 21530 30296 21552
rect 29923 21496 29984 21530
rect 30030 21518 30074 21530
rect 30130 21518 30164 21530
rect 30230 21518 30254 21530
rect 30018 21496 30074 21518
rect 30108 21496 30164 21518
rect 30198 21496 30254 21518
rect 30288 21518 30296 21530
rect 30330 21530 30396 21552
rect 30330 21518 30344 21530
rect 30288 21496 30344 21518
rect 30378 21518 30396 21530
rect 30430 21530 30496 21552
rect 30530 21530 30617 21552
rect 30430 21518 30434 21530
rect 30378 21496 30434 21518
rect 30468 21518 30496 21530
rect 30468 21496 30524 21518
rect 30558 21496 30617 21530
rect 29923 21452 30617 21496
rect 29923 21440 29996 21452
rect 30030 21440 30096 21452
rect 30130 21440 30196 21452
rect 30230 21440 30296 21452
rect 29923 21406 29984 21440
rect 30030 21418 30074 21440
rect 30130 21418 30164 21440
rect 30230 21418 30254 21440
rect 30018 21406 30074 21418
rect 30108 21406 30164 21418
rect 30198 21406 30254 21418
rect 30288 21418 30296 21440
rect 30330 21440 30396 21452
rect 30330 21418 30344 21440
rect 30288 21406 30344 21418
rect 30378 21418 30396 21440
rect 30430 21440 30496 21452
rect 30530 21440 30617 21452
rect 30430 21418 30434 21440
rect 30378 21406 30434 21418
rect 30468 21418 30496 21440
rect 30468 21406 30524 21418
rect 30558 21406 30617 21440
rect 29923 21345 30617 21406
rect 30679 21988 30751 22044
rect 30679 21954 30698 21988
rect 30732 21954 30751 21988
rect 30679 21898 30751 21954
rect 30679 21864 30698 21898
rect 30732 21864 30751 21898
rect 30679 21808 30751 21864
rect 30679 21774 30698 21808
rect 30732 21774 30751 21808
rect 30679 21718 30751 21774
rect 30679 21684 30698 21718
rect 30732 21684 30751 21718
rect 30679 21628 30751 21684
rect 30679 21594 30698 21628
rect 30732 21594 30751 21628
rect 30679 21538 30751 21594
rect 30679 21504 30698 21538
rect 30732 21504 30751 21538
rect 30679 21448 30751 21504
rect 30679 21414 30698 21448
rect 30732 21414 30751 21448
rect 30679 21358 30751 21414
rect 29789 21283 29861 21343
rect 30679 21324 30698 21358
rect 30732 21324 30751 21358
rect 30679 21283 30751 21324
rect 29789 21264 30751 21283
rect 29789 21230 29886 21264
rect 29920 21230 29976 21264
rect 30010 21230 30066 21264
rect 30100 21230 30156 21264
rect 30190 21230 30246 21264
rect 30280 21230 30336 21264
rect 30370 21230 30426 21264
rect 30460 21230 30516 21264
rect 30550 21230 30606 21264
rect 30640 21230 30751 21264
rect 29789 21211 30751 21230
rect 30815 22154 30847 22188
rect 30881 22154 31000 22188
rect 31034 22154 31065 22188
rect 32155 22188 32405 22237
rect 30815 22098 31065 22154
rect 30815 22064 30847 22098
rect 30881 22064 31000 22098
rect 31034 22064 31065 22098
rect 30815 22008 31065 22064
rect 30815 21974 30847 22008
rect 30881 21974 31000 22008
rect 31034 21974 31065 22008
rect 30815 21918 31065 21974
rect 30815 21884 30847 21918
rect 30881 21884 31000 21918
rect 31034 21884 31065 21918
rect 30815 21828 31065 21884
rect 30815 21794 30847 21828
rect 30881 21794 31000 21828
rect 31034 21794 31065 21828
rect 30815 21738 31065 21794
rect 30815 21704 30847 21738
rect 30881 21704 31000 21738
rect 31034 21704 31065 21738
rect 30815 21648 31065 21704
rect 30815 21614 30847 21648
rect 30881 21614 31000 21648
rect 31034 21614 31065 21648
rect 30815 21558 31065 21614
rect 30815 21524 30847 21558
rect 30881 21524 31000 21558
rect 31034 21524 31065 21558
rect 30815 21468 31065 21524
rect 30815 21434 30847 21468
rect 30881 21434 31000 21468
rect 31034 21434 31065 21468
rect 30815 21378 31065 21434
rect 30815 21344 30847 21378
rect 30881 21344 31000 21378
rect 31034 21344 31065 21378
rect 30815 21288 31065 21344
rect 30815 21254 30847 21288
rect 30881 21254 31000 21288
rect 31034 21254 31065 21288
rect 29475 21164 29507 21198
rect 29541 21164 29660 21198
rect 29694 21164 29725 21198
rect 29475 21147 29725 21164
rect 30815 21198 31065 21254
rect 31129 22156 32091 22173
rect 31129 22122 31150 22156
rect 31184 22122 31240 22156
rect 31274 22154 31330 22156
rect 31364 22154 31420 22156
rect 31454 22154 31510 22156
rect 31544 22154 31600 22156
rect 31634 22154 31690 22156
rect 31724 22154 31780 22156
rect 31814 22154 31870 22156
rect 31904 22154 31960 22156
rect 31994 22154 32050 22156
rect 31294 22122 31330 22154
rect 31384 22122 31420 22154
rect 31474 22122 31510 22154
rect 31564 22122 31600 22154
rect 31654 22122 31690 22154
rect 31744 22122 31780 22154
rect 31834 22122 31870 22154
rect 31924 22122 31960 22154
rect 32014 22122 32050 22154
rect 32084 22122 32091 22156
rect 31129 22120 31260 22122
rect 31294 22120 31350 22122
rect 31384 22120 31440 22122
rect 31474 22120 31530 22122
rect 31564 22120 31620 22122
rect 31654 22120 31710 22122
rect 31744 22120 31800 22122
rect 31834 22120 31890 22122
rect 31924 22120 31980 22122
rect 32014 22120 32091 22122
rect 31129 22101 32091 22120
rect 31129 22097 31201 22101
rect 31129 22063 31148 22097
rect 31182 22063 31201 22097
rect 31129 22007 31201 22063
rect 32019 22078 32091 22101
rect 32019 22044 32038 22078
rect 32072 22044 32091 22078
rect 31129 21973 31148 22007
rect 31182 21973 31201 22007
rect 31129 21917 31201 21973
rect 31129 21883 31148 21917
rect 31182 21883 31201 21917
rect 31129 21827 31201 21883
rect 31129 21793 31148 21827
rect 31182 21793 31201 21827
rect 31129 21737 31201 21793
rect 31129 21703 31148 21737
rect 31182 21703 31201 21737
rect 31129 21647 31201 21703
rect 31129 21613 31148 21647
rect 31182 21613 31201 21647
rect 31129 21557 31201 21613
rect 31129 21523 31148 21557
rect 31182 21523 31201 21557
rect 31129 21467 31201 21523
rect 31129 21433 31148 21467
rect 31182 21433 31201 21467
rect 31129 21377 31201 21433
rect 31129 21343 31148 21377
rect 31182 21343 31201 21377
rect 31263 21980 31957 22039
rect 31263 21946 31324 21980
rect 31358 21952 31414 21980
rect 31448 21952 31504 21980
rect 31538 21952 31594 21980
rect 31370 21946 31414 21952
rect 31470 21946 31504 21952
rect 31570 21946 31594 21952
rect 31628 21952 31684 21980
rect 31628 21946 31636 21952
rect 31263 21918 31336 21946
rect 31370 21918 31436 21946
rect 31470 21918 31536 21946
rect 31570 21918 31636 21946
rect 31670 21946 31684 21952
rect 31718 21952 31774 21980
rect 31718 21946 31736 21952
rect 31670 21918 31736 21946
rect 31770 21946 31774 21952
rect 31808 21952 31864 21980
rect 31808 21946 31836 21952
rect 31898 21946 31957 21980
rect 31770 21918 31836 21946
rect 31870 21918 31957 21946
rect 31263 21890 31957 21918
rect 31263 21856 31324 21890
rect 31358 21856 31414 21890
rect 31448 21856 31504 21890
rect 31538 21856 31594 21890
rect 31628 21856 31684 21890
rect 31718 21856 31774 21890
rect 31808 21856 31864 21890
rect 31898 21856 31957 21890
rect 31263 21852 31957 21856
rect 31263 21818 31336 21852
rect 31370 21818 31436 21852
rect 31470 21818 31536 21852
rect 31570 21818 31636 21852
rect 31670 21818 31736 21852
rect 31770 21818 31836 21852
rect 31870 21818 31957 21852
rect 31263 21800 31957 21818
rect 31263 21766 31324 21800
rect 31358 21766 31414 21800
rect 31448 21766 31504 21800
rect 31538 21766 31594 21800
rect 31628 21766 31684 21800
rect 31718 21766 31774 21800
rect 31808 21766 31864 21800
rect 31898 21766 31957 21800
rect 31263 21752 31957 21766
rect 31263 21718 31336 21752
rect 31370 21718 31436 21752
rect 31470 21718 31536 21752
rect 31570 21718 31636 21752
rect 31670 21718 31736 21752
rect 31770 21718 31836 21752
rect 31870 21718 31957 21752
rect 31263 21710 31957 21718
rect 31263 21676 31324 21710
rect 31358 21676 31414 21710
rect 31448 21676 31504 21710
rect 31538 21676 31594 21710
rect 31628 21676 31684 21710
rect 31718 21676 31774 21710
rect 31808 21676 31864 21710
rect 31898 21676 31957 21710
rect 31263 21652 31957 21676
rect 31263 21620 31336 21652
rect 31370 21620 31436 21652
rect 31470 21620 31536 21652
rect 31570 21620 31636 21652
rect 31263 21586 31324 21620
rect 31370 21618 31414 21620
rect 31470 21618 31504 21620
rect 31570 21618 31594 21620
rect 31358 21586 31414 21618
rect 31448 21586 31504 21618
rect 31538 21586 31594 21618
rect 31628 21618 31636 21620
rect 31670 21620 31736 21652
rect 31670 21618 31684 21620
rect 31628 21586 31684 21618
rect 31718 21618 31736 21620
rect 31770 21620 31836 21652
rect 31870 21620 31957 21652
rect 31770 21618 31774 21620
rect 31718 21586 31774 21618
rect 31808 21618 31836 21620
rect 31808 21586 31864 21618
rect 31898 21586 31957 21620
rect 31263 21552 31957 21586
rect 31263 21530 31336 21552
rect 31370 21530 31436 21552
rect 31470 21530 31536 21552
rect 31570 21530 31636 21552
rect 31263 21496 31324 21530
rect 31370 21518 31414 21530
rect 31470 21518 31504 21530
rect 31570 21518 31594 21530
rect 31358 21496 31414 21518
rect 31448 21496 31504 21518
rect 31538 21496 31594 21518
rect 31628 21518 31636 21530
rect 31670 21530 31736 21552
rect 31670 21518 31684 21530
rect 31628 21496 31684 21518
rect 31718 21518 31736 21530
rect 31770 21530 31836 21552
rect 31870 21530 31957 21552
rect 31770 21518 31774 21530
rect 31718 21496 31774 21518
rect 31808 21518 31836 21530
rect 31808 21496 31864 21518
rect 31898 21496 31957 21530
rect 31263 21452 31957 21496
rect 31263 21440 31336 21452
rect 31370 21440 31436 21452
rect 31470 21440 31536 21452
rect 31570 21440 31636 21452
rect 31263 21406 31324 21440
rect 31370 21418 31414 21440
rect 31470 21418 31504 21440
rect 31570 21418 31594 21440
rect 31358 21406 31414 21418
rect 31448 21406 31504 21418
rect 31538 21406 31594 21418
rect 31628 21418 31636 21440
rect 31670 21440 31736 21452
rect 31670 21418 31684 21440
rect 31628 21406 31684 21418
rect 31718 21418 31736 21440
rect 31770 21440 31836 21452
rect 31870 21440 31957 21452
rect 31770 21418 31774 21440
rect 31718 21406 31774 21418
rect 31808 21418 31836 21440
rect 31808 21406 31864 21418
rect 31898 21406 31957 21440
rect 31263 21345 31957 21406
rect 32019 21988 32091 22044
rect 32019 21954 32038 21988
rect 32072 21954 32091 21988
rect 32019 21898 32091 21954
rect 32019 21864 32038 21898
rect 32072 21864 32091 21898
rect 32019 21808 32091 21864
rect 32019 21774 32038 21808
rect 32072 21774 32091 21808
rect 32019 21718 32091 21774
rect 32019 21684 32038 21718
rect 32072 21684 32091 21718
rect 32019 21628 32091 21684
rect 32019 21594 32038 21628
rect 32072 21594 32091 21628
rect 32019 21538 32091 21594
rect 32019 21504 32038 21538
rect 32072 21504 32091 21538
rect 32019 21448 32091 21504
rect 32019 21414 32038 21448
rect 32072 21414 32091 21448
rect 32019 21358 32091 21414
rect 31129 21283 31201 21343
rect 32019 21324 32038 21358
rect 32072 21324 32091 21358
rect 32019 21283 32091 21324
rect 31129 21264 32091 21283
rect 31129 21230 31226 21264
rect 31260 21230 31316 21264
rect 31350 21230 31406 21264
rect 31440 21230 31496 21264
rect 31530 21230 31586 21264
rect 31620 21230 31676 21264
rect 31710 21230 31766 21264
rect 31800 21230 31856 21264
rect 31890 21230 31946 21264
rect 31980 21230 32091 21264
rect 31129 21211 32091 21230
rect 32155 22154 32187 22188
rect 32221 22154 32340 22188
rect 32374 22154 32405 22188
rect 33495 22188 33745 22237
rect 32155 22098 32405 22154
rect 32155 22064 32187 22098
rect 32221 22064 32340 22098
rect 32374 22064 32405 22098
rect 32155 22008 32405 22064
rect 32155 21974 32187 22008
rect 32221 21974 32340 22008
rect 32374 21974 32405 22008
rect 32155 21918 32405 21974
rect 32155 21884 32187 21918
rect 32221 21884 32340 21918
rect 32374 21884 32405 21918
rect 32155 21828 32405 21884
rect 32155 21794 32187 21828
rect 32221 21794 32340 21828
rect 32374 21794 32405 21828
rect 32155 21738 32405 21794
rect 32155 21704 32187 21738
rect 32221 21704 32340 21738
rect 32374 21704 32405 21738
rect 32155 21648 32405 21704
rect 32155 21614 32187 21648
rect 32221 21614 32340 21648
rect 32374 21614 32405 21648
rect 32155 21558 32405 21614
rect 32155 21524 32187 21558
rect 32221 21524 32340 21558
rect 32374 21524 32405 21558
rect 32155 21468 32405 21524
rect 32155 21434 32187 21468
rect 32221 21434 32340 21468
rect 32374 21434 32405 21468
rect 32155 21378 32405 21434
rect 32155 21344 32187 21378
rect 32221 21344 32340 21378
rect 32374 21344 32405 21378
rect 32155 21288 32405 21344
rect 32155 21254 32187 21288
rect 32221 21254 32340 21288
rect 32374 21254 32405 21288
rect 30815 21164 30847 21198
rect 30881 21164 31000 21198
rect 31034 21164 31065 21198
rect 30815 21147 31065 21164
rect 32155 21198 32405 21254
rect 32469 22156 33431 22173
rect 32469 22122 32490 22156
rect 32524 22122 32580 22156
rect 32614 22154 32670 22156
rect 32704 22154 32760 22156
rect 32794 22154 32850 22156
rect 32884 22154 32940 22156
rect 32974 22154 33030 22156
rect 33064 22154 33120 22156
rect 33154 22154 33210 22156
rect 33244 22154 33300 22156
rect 33334 22154 33390 22156
rect 32634 22122 32670 22154
rect 32724 22122 32760 22154
rect 32814 22122 32850 22154
rect 32904 22122 32940 22154
rect 32994 22122 33030 22154
rect 33084 22122 33120 22154
rect 33174 22122 33210 22154
rect 33264 22122 33300 22154
rect 33354 22122 33390 22154
rect 33424 22122 33431 22156
rect 32469 22120 32600 22122
rect 32634 22120 32690 22122
rect 32724 22120 32780 22122
rect 32814 22120 32870 22122
rect 32904 22120 32960 22122
rect 32994 22120 33050 22122
rect 33084 22120 33140 22122
rect 33174 22120 33230 22122
rect 33264 22120 33320 22122
rect 33354 22120 33431 22122
rect 32469 22101 33431 22120
rect 32469 22097 32541 22101
rect 32469 22063 32488 22097
rect 32522 22063 32541 22097
rect 32469 22007 32541 22063
rect 33359 22078 33431 22101
rect 33359 22044 33378 22078
rect 33412 22044 33431 22078
rect 32469 21973 32488 22007
rect 32522 21973 32541 22007
rect 32469 21917 32541 21973
rect 32469 21883 32488 21917
rect 32522 21883 32541 21917
rect 32469 21827 32541 21883
rect 32469 21793 32488 21827
rect 32522 21793 32541 21827
rect 32469 21737 32541 21793
rect 32469 21703 32488 21737
rect 32522 21703 32541 21737
rect 32469 21647 32541 21703
rect 32469 21613 32488 21647
rect 32522 21613 32541 21647
rect 32469 21557 32541 21613
rect 32469 21523 32488 21557
rect 32522 21523 32541 21557
rect 32469 21467 32541 21523
rect 32469 21433 32488 21467
rect 32522 21433 32541 21467
rect 32469 21377 32541 21433
rect 32469 21343 32488 21377
rect 32522 21343 32541 21377
rect 32603 21980 33297 22039
rect 32603 21946 32664 21980
rect 32698 21952 32754 21980
rect 32788 21952 32844 21980
rect 32878 21952 32934 21980
rect 32710 21946 32754 21952
rect 32810 21946 32844 21952
rect 32910 21946 32934 21952
rect 32968 21952 33024 21980
rect 32968 21946 32976 21952
rect 32603 21918 32676 21946
rect 32710 21918 32776 21946
rect 32810 21918 32876 21946
rect 32910 21918 32976 21946
rect 33010 21946 33024 21952
rect 33058 21952 33114 21980
rect 33058 21946 33076 21952
rect 33010 21918 33076 21946
rect 33110 21946 33114 21952
rect 33148 21952 33204 21980
rect 33148 21946 33176 21952
rect 33238 21946 33297 21980
rect 33110 21918 33176 21946
rect 33210 21918 33297 21946
rect 32603 21890 33297 21918
rect 32603 21856 32664 21890
rect 32698 21856 32754 21890
rect 32788 21856 32844 21890
rect 32878 21856 32934 21890
rect 32968 21856 33024 21890
rect 33058 21856 33114 21890
rect 33148 21856 33204 21890
rect 33238 21856 33297 21890
rect 32603 21852 33297 21856
rect 32603 21818 32676 21852
rect 32710 21818 32776 21852
rect 32810 21818 32876 21852
rect 32910 21818 32976 21852
rect 33010 21818 33076 21852
rect 33110 21818 33176 21852
rect 33210 21818 33297 21852
rect 32603 21800 33297 21818
rect 32603 21766 32664 21800
rect 32698 21766 32754 21800
rect 32788 21766 32844 21800
rect 32878 21766 32934 21800
rect 32968 21766 33024 21800
rect 33058 21766 33114 21800
rect 33148 21766 33204 21800
rect 33238 21766 33297 21800
rect 32603 21752 33297 21766
rect 32603 21718 32676 21752
rect 32710 21718 32776 21752
rect 32810 21718 32876 21752
rect 32910 21718 32976 21752
rect 33010 21718 33076 21752
rect 33110 21718 33176 21752
rect 33210 21718 33297 21752
rect 32603 21710 33297 21718
rect 32603 21676 32664 21710
rect 32698 21676 32754 21710
rect 32788 21676 32844 21710
rect 32878 21676 32934 21710
rect 32968 21676 33024 21710
rect 33058 21676 33114 21710
rect 33148 21676 33204 21710
rect 33238 21676 33297 21710
rect 32603 21652 33297 21676
rect 32603 21620 32676 21652
rect 32710 21620 32776 21652
rect 32810 21620 32876 21652
rect 32910 21620 32976 21652
rect 32603 21586 32664 21620
rect 32710 21618 32754 21620
rect 32810 21618 32844 21620
rect 32910 21618 32934 21620
rect 32698 21586 32754 21618
rect 32788 21586 32844 21618
rect 32878 21586 32934 21618
rect 32968 21618 32976 21620
rect 33010 21620 33076 21652
rect 33010 21618 33024 21620
rect 32968 21586 33024 21618
rect 33058 21618 33076 21620
rect 33110 21620 33176 21652
rect 33210 21620 33297 21652
rect 33110 21618 33114 21620
rect 33058 21586 33114 21618
rect 33148 21618 33176 21620
rect 33148 21586 33204 21618
rect 33238 21586 33297 21620
rect 32603 21552 33297 21586
rect 32603 21530 32676 21552
rect 32710 21530 32776 21552
rect 32810 21530 32876 21552
rect 32910 21530 32976 21552
rect 32603 21496 32664 21530
rect 32710 21518 32754 21530
rect 32810 21518 32844 21530
rect 32910 21518 32934 21530
rect 32698 21496 32754 21518
rect 32788 21496 32844 21518
rect 32878 21496 32934 21518
rect 32968 21518 32976 21530
rect 33010 21530 33076 21552
rect 33010 21518 33024 21530
rect 32968 21496 33024 21518
rect 33058 21518 33076 21530
rect 33110 21530 33176 21552
rect 33210 21530 33297 21552
rect 33110 21518 33114 21530
rect 33058 21496 33114 21518
rect 33148 21518 33176 21530
rect 33148 21496 33204 21518
rect 33238 21496 33297 21530
rect 32603 21452 33297 21496
rect 32603 21440 32676 21452
rect 32710 21440 32776 21452
rect 32810 21440 32876 21452
rect 32910 21440 32976 21452
rect 32603 21406 32664 21440
rect 32710 21418 32754 21440
rect 32810 21418 32844 21440
rect 32910 21418 32934 21440
rect 32698 21406 32754 21418
rect 32788 21406 32844 21418
rect 32878 21406 32934 21418
rect 32968 21418 32976 21440
rect 33010 21440 33076 21452
rect 33010 21418 33024 21440
rect 32968 21406 33024 21418
rect 33058 21418 33076 21440
rect 33110 21440 33176 21452
rect 33210 21440 33297 21452
rect 33110 21418 33114 21440
rect 33058 21406 33114 21418
rect 33148 21418 33176 21440
rect 33148 21406 33204 21418
rect 33238 21406 33297 21440
rect 32603 21345 33297 21406
rect 33359 21988 33431 22044
rect 33359 21954 33378 21988
rect 33412 21954 33431 21988
rect 33359 21898 33431 21954
rect 33359 21864 33378 21898
rect 33412 21864 33431 21898
rect 33359 21808 33431 21864
rect 33359 21774 33378 21808
rect 33412 21774 33431 21808
rect 33359 21718 33431 21774
rect 33359 21684 33378 21718
rect 33412 21684 33431 21718
rect 33359 21628 33431 21684
rect 33359 21594 33378 21628
rect 33412 21594 33431 21628
rect 33359 21538 33431 21594
rect 33359 21504 33378 21538
rect 33412 21504 33431 21538
rect 33359 21448 33431 21504
rect 33359 21414 33378 21448
rect 33412 21414 33431 21448
rect 33359 21358 33431 21414
rect 32469 21283 32541 21343
rect 33359 21324 33378 21358
rect 33412 21324 33431 21358
rect 33359 21283 33431 21324
rect 32469 21264 33431 21283
rect 32469 21230 32566 21264
rect 32600 21230 32656 21264
rect 32690 21230 32746 21264
rect 32780 21230 32836 21264
rect 32870 21230 32926 21264
rect 32960 21230 33016 21264
rect 33050 21230 33106 21264
rect 33140 21230 33196 21264
rect 33230 21230 33286 21264
rect 33320 21230 33431 21264
rect 32469 21211 33431 21230
rect 33495 22154 33527 22188
rect 33561 22154 33680 22188
rect 33714 22154 33745 22188
rect 34835 22188 35085 22237
rect 33495 22098 33745 22154
rect 33495 22064 33527 22098
rect 33561 22064 33680 22098
rect 33714 22064 33745 22098
rect 33495 22008 33745 22064
rect 33495 21974 33527 22008
rect 33561 21974 33680 22008
rect 33714 21974 33745 22008
rect 33495 21918 33745 21974
rect 33495 21884 33527 21918
rect 33561 21884 33680 21918
rect 33714 21884 33745 21918
rect 33495 21828 33745 21884
rect 33495 21794 33527 21828
rect 33561 21794 33680 21828
rect 33714 21794 33745 21828
rect 33495 21738 33745 21794
rect 33495 21704 33527 21738
rect 33561 21704 33680 21738
rect 33714 21704 33745 21738
rect 33495 21648 33745 21704
rect 33495 21614 33527 21648
rect 33561 21614 33680 21648
rect 33714 21614 33745 21648
rect 33495 21558 33745 21614
rect 33495 21524 33527 21558
rect 33561 21524 33680 21558
rect 33714 21524 33745 21558
rect 33495 21468 33745 21524
rect 33495 21434 33527 21468
rect 33561 21434 33680 21468
rect 33714 21434 33745 21468
rect 33495 21378 33745 21434
rect 33495 21344 33527 21378
rect 33561 21344 33680 21378
rect 33714 21344 33745 21378
rect 33495 21288 33745 21344
rect 33495 21254 33527 21288
rect 33561 21254 33680 21288
rect 33714 21254 33745 21288
rect 32155 21164 32187 21198
rect 32221 21164 32340 21198
rect 32374 21164 32405 21198
rect 32155 21147 32405 21164
rect 33495 21198 33745 21254
rect 33809 22156 34771 22173
rect 33809 22122 33830 22156
rect 33864 22122 33920 22156
rect 33954 22154 34010 22156
rect 34044 22154 34100 22156
rect 34134 22154 34190 22156
rect 34224 22154 34280 22156
rect 34314 22154 34370 22156
rect 34404 22154 34460 22156
rect 34494 22154 34550 22156
rect 34584 22154 34640 22156
rect 34674 22154 34730 22156
rect 33974 22122 34010 22154
rect 34064 22122 34100 22154
rect 34154 22122 34190 22154
rect 34244 22122 34280 22154
rect 34334 22122 34370 22154
rect 34424 22122 34460 22154
rect 34514 22122 34550 22154
rect 34604 22122 34640 22154
rect 34694 22122 34730 22154
rect 34764 22122 34771 22156
rect 33809 22120 33940 22122
rect 33974 22120 34030 22122
rect 34064 22120 34120 22122
rect 34154 22120 34210 22122
rect 34244 22120 34300 22122
rect 34334 22120 34390 22122
rect 34424 22120 34480 22122
rect 34514 22120 34570 22122
rect 34604 22120 34660 22122
rect 34694 22120 34771 22122
rect 33809 22101 34771 22120
rect 33809 22097 33881 22101
rect 33809 22063 33828 22097
rect 33862 22063 33881 22097
rect 33809 22007 33881 22063
rect 34699 22078 34771 22101
rect 34699 22044 34718 22078
rect 34752 22044 34771 22078
rect 33809 21973 33828 22007
rect 33862 21973 33881 22007
rect 33809 21917 33881 21973
rect 33809 21883 33828 21917
rect 33862 21883 33881 21917
rect 33809 21827 33881 21883
rect 33809 21793 33828 21827
rect 33862 21793 33881 21827
rect 33809 21737 33881 21793
rect 33809 21703 33828 21737
rect 33862 21703 33881 21737
rect 33809 21647 33881 21703
rect 33809 21613 33828 21647
rect 33862 21613 33881 21647
rect 33809 21557 33881 21613
rect 33809 21523 33828 21557
rect 33862 21523 33881 21557
rect 33809 21467 33881 21523
rect 33809 21433 33828 21467
rect 33862 21433 33881 21467
rect 33809 21377 33881 21433
rect 33809 21343 33828 21377
rect 33862 21343 33881 21377
rect 33943 21980 34637 22039
rect 33943 21946 34004 21980
rect 34038 21952 34094 21980
rect 34128 21952 34184 21980
rect 34218 21952 34274 21980
rect 34050 21946 34094 21952
rect 34150 21946 34184 21952
rect 34250 21946 34274 21952
rect 34308 21952 34364 21980
rect 34308 21946 34316 21952
rect 33943 21918 34016 21946
rect 34050 21918 34116 21946
rect 34150 21918 34216 21946
rect 34250 21918 34316 21946
rect 34350 21946 34364 21952
rect 34398 21952 34454 21980
rect 34398 21946 34416 21952
rect 34350 21918 34416 21946
rect 34450 21946 34454 21952
rect 34488 21952 34544 21980
rect 34488 21946 34516 21952
rect 34578 21946 34637 21980
rect 34450 21918 34516 21946
rect 34550 21918 34637 21946
rect 33943 21890 34637 21918
rect 33943 21856 34004 21890
rect 34038 21856 34094 21890
rect 34128 21856 34184 21890
rect 34218 21856 34274 21890
rect 34308 21856 34364 21890
rect 34398 21856 34454 21890
rect 34488 21856 34544 21890
rect 34578 21856 34637 21890
rect 33943 21852 34637 21856
rect 33943 21818 34016 21852
rect 34050 21818 34116 21852
rect 34150 21818 34216 21852
rect 34250 21818 34316 21852
rect 34350 21818 34416 21852
rect 34450 21818 34516 21852
rect 34550 21818 34637 21852
rect 33943 21800 34637 21818
rect 33943 21766 34004 21800
rect 34038 21766 34094 21800
rect 34128 21766 34184 21800
rect 34218 21766 34274 21800
rect 34308 21766 34364 21800
rect 34398 21766 34454 21800
rect 34488 21766 34544 21800
rect 34578 21766 34637 21800
rect 33943 21752 34637 21766
rect 33943 21718 34016 21752
rect 34050 21718 34116 21752
rect 34150 21718 34216 21752
rect 34250 21718 34316 21752
rect 34350 21718 34416 21752
rect 34450 21718 34516 21752
rect 34550 21718 34637 21752
rect 33943 21710 34637 21718
rect 33943 21676 34004 21710
rect 34038 21676 34094 21710
rect 34128 21676 34184 21710
rect 34218 21676 34274 21710
rect 34308 21676 34364 21710
rect 34398 21676 34454 21710
rect 34488 21676 34544 21710
rect 34578 21676 34637 21710
rect 33943 21652 34637 21676
rect 33943 21620 34016 21652
rect 34050 21620 34116 21652
rect 34150 21620 34216 21652
rect 34250 21620 34316 21652
rect 33943 21586 34004 21620
rect 34050 21618 34094 21620
rect 34150 21618 34184 21620
rect 34250 21618 34274 21620
rect 34038 21586 34094 21618
rect 34128 21586 34184 21618
rect 34218 21586 34274 21618
rect 34308 21618 34316 21620
rect 34350 21620 34416 21652
rect 34350 21618 34364 21620
rect 34308 21586 34364 21618
rect 34398 21618 34416 21620
rect 34450 21620 34516 21652
rect 34550 21620 34637 21652
rect 34450 21618 34454 21620
rect 34398 21586 34454 21618
rect 34488 21618 34516 21620
rect 34488 21586 34544 21618
rect 34578 21586 34637 21620
rect 33943 21552 34637 21586
rect 33943 21530 34016 21552
rect 34050 21530 34116 21552
rect 34150 21530 34216 21552
rect 34250 21530 34316 21552
rect 33943 21496 34004 21530
rect 34050 21518 34094 21530
rect 34150 21518 34184 21530
rect 34250 21518 34274 21530
rect 34038 21496 34094 21518
rect 34128 21496 34184 21518
rect 34218 21496 34274 21518
rect 34308 21518 34316 21530
rect 34350 21530 34416 21552
rect 34350 21518 34364 21530
rect 34308 21496 34364 21518
rect 34398 21518 34416 21530
rect 34450 21530 34516 21552
rect 34550 21530 34637 21552
rect 34450 21518 34454 21530
rect 34398 21496 34454 21518
rect 34488 21518 34516 21530
rect 34488 21496 34544 21518
rect 34578 21496 34637 21530
rect 33943 21452 34637 21496
rect 33943 21440 34016 21452
rect 34050 21440 34116 21452
rect 34150 21440 34216 21452
rect 34250 21440 34316 21452
rect 33943 21406 34004 21440
rect 34050 21418 34094 21440
rect 34150 21418 34184 21440
rect 34250 21418 34274 21440
rect 34038 21406 34094 21418
rect 34128 21406 34184 21418
rect 34218 21406 34274 21418
rect 34308 21418 34316 21440
rect 34350 21440 34416 21452
rect 34350 21418 34364 21440
rect 34308 21406 34364 21418
rect 34398 21418 34416 21440
rect 34450 21440 34516 21452
rect 34550 21440 34637 21452
rect 34450 21418 34454 21440
rect 34398 21406 34454 21418
rect 34488 21418 34516 21440
rect 34488 21406 34544 21418
rect 34578 21406 34637 21440
rect 33943 21345 34637 21406
rect 34699 21988 34771 22044
rect 34699 21954 34718 21988
rect 34752 21954 34771 21988
rect 34699 21898 34771 21954
rect 34699 21864 34718 21898
rect 34752 21864 34771 21898
rect 34699 21808 34771 21864
rect 34699 21774 34718 21808
rect 34752 21774 34771 21808
rect 34699 21718 34771 21774
rect 34699 21684 34718 21718
rect 34752 21684 34771 21718
rect 34699 21628 34771 21684
rect 34699 21594 34718 21628
rect 34752 21594 34771 21628
rect 34699 21538 34771 21594
rect 34699 21504 34718 21538
rect 34752 21504 34771 21538
rect 34699 21448 34771 21504
rect 34699 21414 34718 21448
rect 34752 21414 34771 21448
rect 34699 21358 34771 21414
rect 33809 21283 33881 21343
rect 34699 21324 34718 21358
rect 34752 21324 34771 21358
rect 34699 21283 34771 21324
rect 33809 21264 34771 21283
rect 33809 21230 33906 21264
rect 33940 21230 33996 21264
rect 34030 21230 34086 21264
rect 34120 21230 34176 21264
rect 34210 21230 34266 21264
rect 34300 21230 34356 21264
rect 34390 21230 34446 21264
rect 34480 21230 34536 21264
rect 34570 21230 34626 21264
rect 34660 21230 34771 21264
rect 33809 21211 34771 21230
rect 34835 22154 34867 22188
rect 34901 22154 35020 22188
rect 35054 22154 35085 22188
rect 36175 22188 36425 22237
rect 34835 22098 35085 22154
rect 34835 22064 34867 22098
rect 34901 22064 35020 22098
rect 35054 22064 35085 22098
rect 34835 22008 35085 22064
rect 34835 21974 34867 22008
rect 34901 21974 35020 22008
rect 35054 21974 35085 22008
rect 34835 21918 35085 21974
rect 34835 21884 34867 21918
rect 34901 21884 35020 21918
rect 35054 21884 35085 21918
rect 34835 21828 35085 21884
rect 34835 21794 34867 21828
rect 34901 21794 35020 21828
rect 35054 21794 35085 21828
rect 34835 21738 35085 21794
rect 34835 21704 34867 21738
rect 34901 21704 35020 21738
rect 35054 21704 35085 21738
rect 34835 21648 35085 21704
rect 34835 21614 34867 21648
rect 34901 21614 35020 21648
rect 35054 21614 35085 21648
rect 34835 21558 35085 21614
rect 34835 21524 34867 21558
rect 34901 21524 35020 21558
rect 35054 21524 35085 21558
rect 34835 21468 35085 21524
rect 34835 21434 34867 21468
rect 34901 21434 35020 21468
rect 35054 21434 35085 21468
rect 34835 21378 35085 21434
rect 34835 21344 34867 21378
rect 34901 21344 35020 21378
rect 35054 21344 35085 21378
rect 34835 21288 35085 21344
rect 34835 21254 34867 21288
rect 34901 21254 35020 21288
rect 35054 21254 35085 21288
rect 33495 21164 33527 21198
rect 33561 21164 33680 21198
rect 33714 21164 33745 21198
rect 33495 21147 33745 21164
rect 34835 21198 35085 21254
rect 35149 22156 36111 22173
rect 35149 22122 35170 22156
rect 35204 22122 35260 22156
rect 35294 22154 35350 22156
rect 35384 22154 35440 22156
rect 35474 22154 35530 22156
rect 35564 22154 35620 22156
rect 35654 22154 35710 22156
rect 35744 22154 35800 22156
rect 35834 22154 35890 22156
rect 35924 22154 35980 22156
rect 36014 22154 36070 22156
rect 35314 22122 35350 22154
rect 35404 22122 35440 22154
rect 35494 22122 35530 22154
rect 35584 22122 35620 22154
rect 35674 22122 35710 22154
rect 35764 22122 35800 22154
rect 35854 22122 35890 22154
rect 35944 22122 35980 22154
rect 36034 22122 36070 22154
rect 36104 22122 36111 22156
rect 35149 22120 35280 22122
rect 35314 22120 35370 22122
rect 35404 22120 35460 22122
rect 35494 22120 35550 22122
rect 35584 22120 35640 22122
rect 35674 22120 35730 22122
rect 35764 22120 35820 22122
rect 35854 22120 35910 22122
rect 35944 22120 36000 22122
rect 36034 22120 36111 22122
rect 35149 22101 36111 22120
rect 35149 22097 35221 22101
rect 35149 22063 35168 22097
rect 35202 22063 35221 22097
rect 35149 22007 35221 22063
rect 36039 22078 36111 22101
rect 36039 22044 36058 22078
rect 36092 22044 36111 22078
rect 35149 21973 35168 22007
rect 35202 21973 35221 22007
rect 35149 21917 35221 21973
rect 35149 21883 35168 21917
rect 35202 21883 35221 21917
rect 35149 21827 35221 21883
rect 35149 21793 35168 21827
rect 35202 21793 35221 21827
rect 35149 21737 35221 21793
rect 35149 21703 35168 21737
rect 35202 21703 35221 21737
rect 35149 21647 35221 21703
rect 35149 21613 35168 21647
rect 35202 21613 35221 21647
rect 35149 21557 35221 21613
rect 35149 21523 35168 21557
rect 35202 21523 35221 21557
rect 35149 21467 35221 21523
rect 35149 21433 35168 21467
rect 35202 21433 35221 21467
rect 35149 21377 35221 21433
rect 35149 21343 35168 21377
rect 35202 21343 35221 21377
rect 35283 21980 35977 22039
rect 35283 21946 35344 21980
rect 35378 21952 35434 21980
rect 35468 21952 35524 21980
rect 35558 21952 35614 21980
rect 35390 21946 35434 21952
rect 35490 21946 35524 21952
rect 35590 21946 35614 21952
rect 35648 21952 35704 21980
rect 35648 21946 35656 21952
rect 35283 21918 35356 21946
rect 35390 21918 35456 21946
rect 35490 21918 35556 21946
rect 35590 21918 35656 21946
rect 35690 21946 35704 21952
rect 35738 21952 35794 21980
rect 35738 21946 35756 21952
rect 35690 21918 35756 21946
rect 35790 21946 35794 21952
rect 35828 21952 35884 21980
rect 35828 21946 35856 21952
rect 35918 21946 35977 21980
rect 35790 21918 35856 21946
rect 35890 21918 35977 21946
rect 35283 21890 35977 21918
rect 35283 21856 35344 21890
rect 35378 21856 35434 21890
rect 35468 21856 35524 21890
rect 35558 21856 35614 21890
rect 35648 21856 35704 21890
rect 35738 21856 35794 21890
rect 35828 21856 35884 21890
rect 35918 21856 35977 21890
rect 35283 21852 35977 21856
rect 35283 21818 35356 21852
rect 35390 21818 35456 21852
rect 35490 21818 35556 21852
rect 35590 21818 35656 21852
rect 35690 21818 35756 21852
rect 35790 21818 35856 21852
rect 35890 21818 35977 21852
rect 35283 21800 35977 21818
rect 35283 21766 35344 21800
rect 35378 21766 35434 21800
rect 35468 21766 35524 21800
rect 35558 21766 35614 21800
rect 35648 21766 35704 21800
rect 35738 21766 35794 21800
rect 35828 21766 35884 21800
rect 35918 21766 35977 21800
rect 35283 21752 35977 21766
rect 35283 21718 35356 21752
rect 35390 21718 35456 21752
rect 35490 21718 35556 21752
rect 35590 21718 35656 21752
rect 35690 21718 35756 21752
rect 35790 21718 35856 21752
rect 35890 21718 35977 21752
rect 35283 21710 35977 21718
rect 35283 21676 35344 21710
rect 35378 21676 35434 21710
rect 35468 21676 35524 21710
rect 35558 21676 35614 21710
rect 35648 21676 35704 21710
rect 35738 21676 35794 21710
rect 35828 21676 35884 21710
rect 35918 21676 35977 21710
rect 35283 21652 35977 21676
rect 35283 21620 35356 21652
rect 35390 21620 35456 21652
rect 35490 21620 35556 21652
rect 35590 21620 35656 21652
rect 35283 21586 35344 21620
rect 35390 21618 35434 21620
rect 35490 21618 35524 21620
rect 35590 21618 35614 21620
rect 35378 21586 35434 21618
rect 35468 21586 35524 21618
rect 35558 21586 35614 21618
rect 35648 21618 35656 21620
rect 35690 21620 35756 21652
rect 35690 21618 35704 21620
rect 35648 21586 35704 21618
rect 35738 21618 35756 21620
rect 35790 21620 35856 21652
rect 35890 21620 35977 21652
rect 35790 21618 35794 21620
rect 35738 21586 35794 21618
rect 35828 21618 35856 21620
rect 35828 21586 35884 21618
rect 35918 21586 35977 21620
rect 35283 21552 35977 21586
rect 35283 21530 35356 21552
rect 35390 21530 35456 21552
rect 35490 21530 35556 21552
rect 35590 21530 35656 21552
rect 35283 21496 35344 21530
rect 35390 21518 35434 21530
rect 35490 21518 35524 21530
rect 35590 21518 35614 21530
rect 35378 21496 35434 21518
rect 35468 21496 35524 21518
rect 35558 21496 35614 21518
rect 35648 21518 35656 21530
rect 35690 21530 35756 21552
rect 35690 21518 35704 21530
rect 35648 21496 35704 21518
rect 35738 21518 35756 21530
rect 35790 21530 35856 21552
rect 35890 21530 35977 21552
rect 35790 21518 35794 21530
rect 35738 21496 35794 21518
rect 35828 21518 35856 21530
rect 35828 21496 35884 21518
rect 35918 21496 35977 21530
rect 35283 21452 35977 21496
rect 35283 21440 35356 21452
rect 35390 21440 35456 21452
rect 35490 21440 35556 21452
rect 35590 21440 35656 21452
rect 35283 21406 35344 21440
rect 35390 21418 35434 21440
rect 35490 21418 35524 21440
rect 35590 21418 35614 21440
rect 35378 21406 35434 21418
rect 35468 21406 35524 21418
rect 35558 21406 35614 21418
rect 35648 21418 35656 21440
rect 35690 21440 35756 21452
rect 35690 21418 35704 21440
rect 35648 21406 35704 21418
rect 35738 21418 35756 21440
rect 35790 21440 35856 21452
rect 35890 21440 35977 21452
rect 35790 21418 35794 21440
rect 35738 21406 35794 21418
rect 35828 21418 35856 21440
rect 35828 21406 35884 21418
rect 35918 21406 35977 21440
rect 35283 21345 35977 21406
rect 36039 21988 36111 22044
rect 36039 21954 36058 21988
rect 36092 21954 36111 21988
rect 36039 21898 36111 21954
rect 36039 21864 36058 21898
rect 36092 21864 36111 21898
rect 36039 21808 36111 21864
rect 36039 21774 36058 21808
rect 36092 21774 36111 21808
rect 36039 21718 36111 21774
rect 36039 21684 36058 21718
rect 36092 21684 36111 21718
rect 36039 21628 36111 21684
rect 36039 21594 36058 21628
rect 36092 21594 36111 21628
rect 36039 21538 36111 21594
rect 36039 21504 36058 21538
rect 36092 21504 36111 21538
rect 36039 21448 36111 21504
rect 36039 21414 36058 21448
rect 36092 21414 36111 21448
rect 36039 21358 36111 21414
rect 35149 21283 35221 21343
rect 36039 21324 36058 21358
rect 36092 21324 36111 21358
rect 36039 21283 36111 21324
rect 35149 21264 36111 21283
rect 35149 21230 35246 21264
rect 35280 21230 35336 21264
rect 35370 21230 35426 21264
rect 35460 21230 35516 21264
rect 35550 21230 35606 21264
rect 35640 21230 35696 21264
rect 35730 21230 35786 21264
rect 35820 21230 35876 21264
rect 35910 21230 35966 21264
rect 36000 21230 36111 21264
rect 35149 21211 36111 21230
rect 36175 22154 36207 22188
rect 36241 22154 36360 22188
rect 36394 22154 36425 22188
rect 37515 22188 37765 22237
rect 36175 22098 36425 22154
rect 36175 22064 36207 22098
rect 36241 22064 36360 22098
rect 36394 22064 36425 22098
rect 36175 22008 36425 22064
rect 36175 21974 36207 22008
rect 36241 21974 36360 22008
rect 36394 21974 36425 22008
rect 36175 21918 36425 21974
rect 36175 21884 36207 21918
rect 36241 21884 36360 21918
rect 36394 21884 36425 21918
rect 36175 21828 36425 21884
rect 36175 21794 36207 21828
rect 36241 21794 36360 21828
rect 36394 21794 36425 21828
rect 36175 21738 36425 21794
rect 36175 21704 36207 21738
rect 36241 21704 36360 21738
rect 36394 21704 36425 21738
rect 36175 21648 36425 21704
rect 36175 21614 36207 21648
rect 36241 21614 36360 21648
rect 36394 21614 36425 21648
rect 36175 21558 36425 21614
rect 36175 21524 36207 21558
rect 36241 21524 36360 21558
rect 36394 21524 36425 21558
rect 36175 21468 36425 21524
rect 36175 21434 36207 21468
rect 36241 21434 36360 21468
rect 36394 21434 36425 21468
rect 36175 21378 36425 21434
rect 36175 21344 36207 21378
rect 36241 21344 36360 21378
rect 36394 21344 36425 21378
rect 36175 21288 36425 21344
rect 36175 21254 36207 21288
rect 36241 21254 36360 21288
rect 36394 21254 36425 21288
rect 34835 21164 34867 21198
rect 34901 21164 35020 21198
rect 35054 21164 35085 21198
rect 34835 21147 35085 21164
rect 36175 21198 36425 21254
rect 36489 22156 37451 22173
rect 36489 22122 36510 22156
rect 36544 22122 36600 22156
rect 36634 22154 36690 22156
rect 36724 22154 36780 22156
rect 36814 22154 36870 22156
rect 36904 22154 36960 22156
rect 36994 22154 37050 22156
rect 37084 22154 37140 22156
rect 37174 22154 37230 22156
rect 37264 22154 37320 22156
rect 37354 22154 37410 22156
rect 36654 22122 36690 22154
rect 36744 22122 36780 22154
rect 36834 22122 36870 22154
rect 36924 22122 36960 22154
rect 37014 22122 37050 22154
rect 37104 22122 37140 22154
rect 37194 22122 37230 22154
rect 37284 22122 37320 22154
rect 37374 22122 37410 22154
rect 37444 22122 37451 22156
rect 36489 22120 36620 22122
rect 36654 22120 36710 22122
rect 36744 22120 36800 22122
rect 36834 22120 36890 22122
rect 36924 22120 36980 22122
rect 37014 22120 37070 22122
rect 37104 22120 37160 22122
rect 37194 22120 37250 22122
rect 37284 22120 37340 22122
rect 37374 22120 37451 22122
rect 36489 22101 37451 22120
rect 36489 22097 36561 22101
rect 36489 22063 36508 22097
rect 36542 22063 36561 22097
rect 36489 22007 36561 22063
rect 37379 22078 37451 22101
rect 37379 22044 37398 22078
rect 37432 22044 37451 22078
rect 36489 21973 36508 22007
rect 36542 21973 36561 22007
rect 36489 21917 36561 21973
rect 36489 21883 36508 21917
rect 36542 21883 36561 21917
rect 36489 21827 36561 21883
rect 36489 21793 36508 21827
rect 36542 21793 36561 21827
rect 36489 21737 36561 21793
rect 36489 21703 36508 21737
rect 36542 21703 36561 21737
rect 36489 21647 36561 21703
rect 36489 21613 36508 21647
rect 36542 21613 36561 21647
rect 36489 21557 36561 21613
rect 36489 21523 36508 21557
rect 36542 21523 36561 21557
rect 36489 21467 36561 21523
rect 36489 21433 36508 21467
rect 36542 21433 36561 21467
rect 36489 21377 36561 21433
rect 36489 21343 36508 21377
rect 36542 21343 36561 21377
rect 36623 21980 37317 22039
rect 36623 21946 36684 21980
rect 36718 21952 36774 21980
rect 36808 21952 36864 21980
rect 36898 21952 36954 21980
rect 36730 21946 36774 21952
rect 36830 21946 36864 21952
rect 36930 21946 36954 21952
rect 36988 21952 37044 21980
rect 36988 21946 36996 21952
rect 36623 21918 36696 21946
rect 36730 21918 36796 21946
rect 36830 21918 36896 21946
rect 36930 21918 36996 21946
rect 37030 21946 37044 21952
rect 37078 21952 37134 21980
rect 37078 21946 37096 21952
rect 37030 21918 37096 21946
rect 37130 21946 37134 21952
rect 37168 21952 37224 21980
rect 37168 21946 37196 21952
rect 37258 21946 37317 21980
rect 37130 21918 37196 21946
rect 37230 21918 37317 21946
rect 36623 21890 37317 21918
rect 36623 21856 36684 21890
rect 36718 21856 36774 21890
rect 36808 21856 36864 21890
rect 36898 21856 36954 21890
rect 36988 21856 37044 21890
rect 37078 21856 37134 21890
rect 37168 21856 37224 21890
rect 37258 21856 37317 21890
rect 36623 21852 37317 21856
rect 36623 21818 36696 21852
rect 36730 21818 36796 21852
rect 36830 21818 36896 21852
rect 36930 21818 36996 21852
rect 37030 21818 37096 21852
rect 37130 21818 37196 21852
rect 37230 21818 37317 21852
rect 36623 21800 37317 21818
rect 36623 21766 36684 21800
rect 36718 21766 36774 21800
rect 36808 21766 36864 21800
rect 36898 21766 36954 21800
rect 36988 21766 37044 21800
rect 37078 21766 37134 21800
rect 37168 21766 37224 21800
rect 37258 21766 37317 21800
rect 36623 21752 37317 21766
rect 36623 21718 36696 21752
rect 36730 21718 36796 21752
rect 36830 21718 36896 21752
rect 36930 21718 36996 21752
rect 37030 21718 37096 21752
rect 37130 21718 37196 21752
rect 37230 21718 37317 21752
rect 36623 21710 37317 21718
rect 36623 21676 36684 21710
rect 36718 21676 36774 21710
rect 36808 21676 36864 21710
rect 36898 21676 36954 21710
rect 36988 21676 37044 21710
rect 37078 21676 37134 21710
rect 37168 21676 37224 21710
rect 37258 21676 37317 21710
rect 36623 21652 37317 21676
rect 36623 21620 36696 21652
rect 36730 21620 36796 21652
rect 36830 21620 36896 21652
rect 36930 21620 36996 21652
rect 36623 21586 36684 21620
rect 36730 21618 36774 21620
rect 36830 21618 36864 21620
rect 36930 21618 36954 21620
rect 36718 21586 36774 21618
rect 36808 21586 36864 21618
rect 36898 21586 36954 21618
rect 36988 21618 36996 21620
rect 37030 21620 37096 21652
rect 37030 21618 37044 21620
rect 36988 21586 37044 21618
rect 37078 21618 37096 21620
rect 37130 21620 37196 21652
rect 37230 21620 37317 21652
rect 37130 21618 37134 21620
rect 37078 21586 37134 21618
rect 37168 21618 37196 21620
rect 37168 21586 37224 21618
rect 37258 21586 37317 21620
rect 36623 21552 37317 21586
rect 36623 21530 36696 21552
rect 36730 21530 36796 21552
rect 36830 21530 36896 21552
rect 36930 21530 36996 21552
rect 36623 21496 36684 21530
rect 36730 21518 36774 21530
rect 36830 21518 36864 21530
rect 36930 21518 36954 21530
rect 36718 21496 36774 21518
rect 36808 21496 36864 21518
rect 36898 21496 36954 21518
rect 36988 21518 36996 21530
rect 37030 21530 37096 21552
rect 37030 21518 37044 21530
rect 36988 21496 37044 21518
rect 37078 21518 37096 21530
rect 37130 21530 37196 21552
rect 37230 21530 37317 21552
rect 37130 21518 37134 21530
rect 37078 21496 37134 21518
rect 37168 21518 37196 21530
rect 37168 21496 37224 21518
rect 37258 21496 37317 21530
rect 36623 21452 37317 21496
rect 36623 21440 36696 21452
rect 36730 21440 36796 21452
rect 36830 21440 36896 21452
rect 36930 21440 36996 21452
rect 36623 21406 36684 21440
rect 36730 21418 36774 21440
rect 36830 21418 36864 21440
rect 36930 21418 36954 21440
rect 36718 21406 36774 21418
rect 36808 21406 36864 21418
rect 36898 21406 36954 21418
rect 36988 21418 36996 21440
rect 37030 21440 37096 21452
rect 37030 21418 37044 21440
rect 36988 21406 37044 21418
rect 37078 21418 37096 21440
rect 37130 21440 37196 21452
rect 37230 21440 37317 21452
rect 37130 21418 37134 21440
rect 37078 21406 37134 21418
rect 37168 21418 37196 21440
rect 37168 21406 37224 21418
rect 37258 21406 37317 21440
rect 36623 21345 37317 21406
rect 37379 21988 37451 22044
rect 37379 21954 37398 21988
rect 37432 21954 37451 21988
rect 37379 21898 37451 21954
rect 37379 21864 37398 21898
rect 37432 21864 37451 21898
rect 37379 21808 37451 21864
rect 37379 21774 37398 21808
rect 37432 21774 37451 21808
rect 37379 21718 37451 21774
rect 37379 21684 37398 21718
rect 37432 21684 37451 21718
rect 37379 21628 37451 21684
rect 37379 21594 37398 21628
rect 37432 21594 37451 21628
rect 37379 21538 37451 21594
rect 37379 21504 37398 21538
rect 37432 21504 37451 21538
rect 37379 21448 37451 21504
rect 37379 21414 37398 21448
rect 37432 21414 37451 21448
rect 37379 21358 37451 21414
rect 36489 21283 36561 21343
rect 37379 21324 37398 21358
rect 37432 21324 37451 21358
rect 37379 21283 37451 21324
rect 36489 21264 37451 21283
rect 36489 21230 36586 21264
rect 36620 21230 36676 21264
rect 36710 21230 36766 21264
rect 36800 21230 36856 21264
rect 36890 21230 36946 21264
rect 36980 21230 37036 21264
rect 37070 21230 37126 21264
rect 37160 21230 37216 21264
rect 37250 21230 37306 21264
rect 37340 21230 37451 21264
rect 36489 21211 37451 21230
rect 37515 22154 37547 22188
rect 37581 22154 37700 22188
rect 37734 22154 37765 22188
rect 38855 22188 38954 22237
rect 37515 22098 37765 22154
rect 37515 22064 37547 22098
rect 37581 22064 37700 22098
rect 37734 22064 37765 22098
rect 37515 22008 37765 22064
rect 37515 21974 37547 22008
rect 37581 21974 37700 22008
rect 37734 21974 37765 22008
rect 37515 21918 37765 21974
rect 37515 21884 37547 21918
rect 37581 21884 37700 21918
rect 37734 21884 37765 21918
rect 37515 21828 37765 21884
rect 37515 21794 37547 21828
rect 37581 21794 37700 21828
rect 37734 21794 37765 21828
rect 37515 21738 37765 21794
rect 37515 21704 37547 21738
rect 37581 21704 37700 21738
rect 37734 21704 37765 21738
rect 37515 21648 37765 21704
rect 37515 21614 37547 21648
rect 37581 21614 37700 21648
rect 37734 21614 37765 21648
rect 37515 21558 37765 21614
rect 37515 21524 37547 21558
rect 37581 21524 37700 21558
rect 37734 21524 37765 21558
rect 37515 21468 37765 21524
rect 37515 21434 37547 21468
rect 37581 21434 37700 21468
rect 37734 21434 37765 21468
rect 37515 21378 37765 21434
rect 37515 21344 37547 21378
rect 37581 21344 37700 21378
rect 37734 21344 37765 21378
rect 37515 21288 37765 21344
rect 37515 21254 37547 21288
rect 37581 21254 37700 21288
rect 37734 21254 37765 21288
rect 36175 21164 36207 21198
rect 36241 21164 36360 21198
rect 36394 21164 36425 21198
rect 36175 21147 36425 21164
rect 37515 21198 37765 21254
rect 37829 22156 38791 22173
rect 37829 22122 37850 22156
rect 37884 22122 37940 22156
rect 37974 22154 38030 22156
rect 38064 22154 38120 22156
rect 38154 22154 38210 22156
rect 38244 22154 38300 22156
rect 38334 22154 38390 22156
rect 38424 22154 38480 22156
rect 38514 22154 38570 22156
rect 38604 22154 38660 22156
rect 38694 22154 38750 22156
rect 37994 22122 38030 22154
rect 38084 22122 38120 22154
rect 38174 22122 38210 22154
rect 38264 22122 38300 22154
rect 38354 22122 38390 22154
rect 38444 22122 38480 22154
rect 38534 22122 38570 22154
rect 38624 22122 38660 22154
rect 38714 22122 38750 22154
rect 38784 22122 38791 22156
rect 37829 22120 37960 22122
rect 37994 22120 38050 22122
rect 38084 22120 38140 22122
rect 38174 22120 38230 22122
rect 38264 22120 38320 22122
rect 38354 22120 38410 22122
rect 38444 22120 38500 22122
rect 38534 22120 38590 22122
rect 38624 22120 38680 22122
rect 38714 22120 38791 22122
rect 37829 22101 38791 22120
rect 37829 22097 37901 22101
rect 37829 22063 37848 22097
rect 37882 22063 37901 22097
rect 37829 22007 37901 22063
rect 38719 22078 38791 22101
rect 38719 22044 38738 22078
rect 38772 22044 38791 22078
rect 37829 21973 37848 22007
rect 37882 21973 37901 22007
rect 37829 21917 37901 21973
rect 37829 21883 37848 21917
rect 37882 21883 37901 21917
rect 37829 21827 37901 21883
rect 37829 21793 37848 21827
rect 37882 21793 37901 21827
rect 37829 21737 37901 21793
rect 37829 21703 37848 21737
rect 37882 21703 37901 21737
rect 37829 21647 37901 21703
rect 37829 21613 37848 21647
rect 37882 21613 37901 21647
rect 37829 21557 37901 21613
rect 37829 21523 37848 21557
rect 37882 21523 37901 21557
rect 37829 21467 37901 21523
rect 37829 21433 37848 21467
rect 37882 21433 37901 21467
rect 37829 21377 37901 21433
rect 37829 21343 37848 21377
rect 37882 21343 37901 21377
rect 37963 21980 38657 22039
rect 37963 21946 38024 21980
rect 38058 21952 38114 21980
rect 38148 21952 38204 21980
rect 38238 21952 38294 21980
rect 38070 21946 38114 21952
rect 38170 21946 38204 21952
rect 38270 21946 38294 21952
rect 38328 21952 38384 21980
rect 38328 21946 38336 21952
rect 37963 21918 38036 21946
rect 38070 21918 38136 21946
rect 38170 21918 38236 21946
rect 38270 21918 38336 21946
rect 38370 21946 38384 21952
rect 38418 21952 38474 21980
rect 38418 21946 38436 21952
rect 38370 21918 38436 21946
rect 38470 21946 38474 21952
rect 38508 21952 38564 21980
rect 38508 21946 38536 21952
rect 38598 21946 38657 21980
rect 38470 21918 38536 21946
rect 38570 21918 38657 21946
rect 37963 21890 38657 21918
rect 37963 21856 38024 21890
rect 38058 21856 38114 21890
rect 38148 21856 38204 21890
rect 38238 21856 38294 21890
rect 38328 21856 38384 21890
rect 38418 21856 38474 21890
rect 38508 21856 38564 21890
rect 38598 21856 38657 21890
rect 37963 21852 38657 21856
rect 37963 21818 38036 21852
rect 38070 21818 38136 21852
rect 38170 21818 38236 21852
rect 38270 21818 38336 21852
rect 38370 21818 38436 21852
rect 38470 21818 38536 21852
rect 38570 21818 38657 21852
rect 37963 21800 38657 21818
rect 37963 21766 38024 21800
rect 38058 21766 38114 21800
rect 38148 21766 38204 21800
rect 38238 21766 38294 21800
rect 38328 21766 38384 21800
rect 38418 21766 38474 21800
rect 38508 21766 38564 21800
rect 38598 21766 38657 21800
rect 37963 21752 38657 21766
rect 37963 21718 38036 21752
rect 38070 21718 38136 21752
rect 38170 21718 38236 21752
rect 38270 21718 38336 21752
rect 38370 21718 38436 21752
rect 38470 21718 38536 21752
rect 38570 21718 38657 21752
rect 37963 21710 38657 21718
rect 37963 21676 38024 21710
rect 38058 21676 38114 21710
rect 38148 21676 38204 21710
rect 38238 21676 38294 21710
rect 38328 21676 38384 21710
rect 38418 21676 38474 21710
rect 38508 21676 38564 21710
rect 38598 21676 38657 21710
rect 37963 21652 38657 21676
rect 37963 21620 38036 21652
rect 38070 21620 38136 21652
rect 38170 21620 38236 21652
rect 38270 21620 38336 21652
rect 37963 21586 38024 21620
rect 38070 21618 38114 21620
rect 38170 21618 38204 21620
rect 38270 21618 38294 21620
rect 38058 21586 38114 21618
rect 38148 21586 38204 21618
rect 38238 21586 38294 21618
rect 38328 21618 38336 21620
rect 38370 21620 38436 21652
rect 38370 21618 38384 21620
rect 38328 21586 38384 21618
rect 38418 21618 38436 21620
rect 38470 21620 38536 21652
rect 38570 21620 38657 21652
rect 38470 21618 38474 21620
rect 38418 21586 38474 21618
rect 38508 21618 38536 21620
rect 38508 21586 38564 21618
rect 38598 21586 38657 21620
rect 37963 21552 38657 21586
rect 37963 21530 38036 21552
rect 38070 21530 38136 21552
rect 38170 21530 38236 21552
rect 38270 21530 38336 21552
rect 37963 21496 38024 21530
rect 38070 21518 38114 21530
rect 38170 21518 38204 21530
rect 38270 21518 38294 21530
rect 38058 21496 38114 21518
rect 38148 21496 38204 21518
rect 38238 21496 38294 21518
rect 38328 21518 38336 21530
rect 38370 21530 38436 21552
rect 38370 21518 38384 21530
rect 38328 21496 38384 21518
rect 38418 21518 38436 21530
rect 38470 21530 38536 21552
rect 38570 21530 38657 21552
rect 38470 21518 38474 21530
rect 38418 21496 38474 21518
rect 38508 21518 38536 21530
rect 38508 21496 38564 21518
rect 38598 21496 38657 21530
rect 37963 21452 38657 21496
rect 37963 21440 38036 21452
rect 38070 21440 38136 21452
rect 38170 21440 38236 21452
rect 38270 21440 38336 21452
rect 37963 21406 38024 21440
rect 38070 21418 38114 21440
rect 38170 21418 38204 21440
rect 38270 21418 38294 21440
rect 38058 21406 38114 21418
rect 38148 21406 38204 21418
rect 38238 21406 38294 21418
rect 38328 21418 38336 21440
rect 38370 21440 38436 21452
rect 38370 21418 38384 21440
rect 38328 21406 38384 21418
rect 38418 21418 38436 21440
rect 38470 21440 38536 21452
rect 38570 21440 38657 21452
rect 38470 21418 38474 21440
rect 38418 21406 38474 21418
rect 38508 21418 38536 21440
rect 38508 21406 38564 21418
rect 38598 21406 38657 21440
rect 37963 21345 38657 21406
rect 38719 21988 38791 22044
rect 38719 21954 38738 21988
rect 38772 21954 38791 21988
rect 38719 21898 38791 21954
rect 38719 21864 38738 21898
rect 38772 21864 38791 21898
rect 38719 21808 38791 21864
rect 38719 21774 38738 21808
rect 38772 21774 38791 21808
rect 38719 21718 38791 21774
rect 38719 21684 38738 21718
rect 38772 21684 38791 21718
rect 38719 21628 38791 21684
rect 38719 21594 38738 21628
rect 38772 21594 38791 21628
rect 38719 21538 38791 21594
rect 38719 21504 38738 21538
rect 38772 21504 38791 21538
rect 38719 21448 38791 21504
rect 38719 21414 38738 21448
rect 38772 21414 38791 21448
rect 38719 21358 38791 21414
rect 37829 21283 37901 21343
rect 38719 21324 38738 21358
rect 38772 21324 38791 21358
rect 38719 21283 38791 21324
rect 37829 21264 38791 21283
rect 37829 21230 37926 21264
rect 37960 21230 38016 21264
rect 38050 21230 38106 21264
rect 38140 21230 38196 21264
rect 38230 21230 38286 21264
rect 38320 21230 38376 21264
rect 38410 21230 38466 21264
rect 38500 21230 38556 21264
rect 38590 21230 38646 21264
rect 38680 21230 38791 21264
rect 37829 21211 38791 21230
rect 38855 22154 38887 22188
rect 38921 22154 38954 22188
rect 38855 22098 38954 22154
rect 38855 22064 38887 22098
rect 38921 22064 38954 22098
rect 38855 22008 38954 22064
rect 38855 21974 38887 22008
rect 38921 21974 38954 22008
rect 38855 21918 38954 21974
rect 38855 21884 38887 21918
rect 38921 21884 38954 21918
rect 38855 21828 38954 21884
rect 38855 21794 38887 21828
rect 38921 21794 38954 21828
rect 38855 21738 38954 21794
rect 38855 21704 38887 21738
rect 38921 21704 38954 21738
rect 38855 21648 38954 21704
rect 38855 21614 38887 21648
rect 38921 21614 38954 21648
rect 38855 21558 38954 21614
rect 38855 21524 38887 21558
rect 38921 21524 38954 21558
rect 38855 21468 38954 21524
rect 38855 21434 38887 21468
rect 38921 21434 38954 21468
rect 40658 21683 41274 21722
rect 40658 21581 40745 21683
rect 41187 21581 41274 21683
rect 38855 21378 38954 21434
rect 38855 21344 38887 21378
rect 38921 21344 38954 21378
rect 38855 21288 38954 21344
rect 38855 21254 38887 21288
rect 38921 21254 38954 21288
rect 37515 21164 37547 21198
rect 37581 21164 37700 21198
rect 37734 21164 37765 21198
rect 37515 21147 37765 21164
rect 38855 21198 38954 21254
rect 38855 21164 38887 21198
rect 38921 21164 38954 21198
rect 38855 21147 38954 21164
rect 21034 21097 21097 21131
rect 21131 21114 22322 21131
rect 21131 21097 21164 21114
rect 21034 21080 21164 21097
rect 21198 21080 21254 21114
rect 21288 21080 21344 21114
rect 21378 21080 21434 21114
rect 21468 21080 21524 21114
rect 21558 21080 21614 21114
rect 21648 21080 21704 21114
rect 21738 21080 21794 21114
rect 21828 21080 21884 21114
rect 21918 21080 21974 21114
rect 22008 21080 22064 21114
rect 22098 21080 22154 21114
rect 22188 21080 22322 21114
rect 21034 21048 22322 21080
rect 23048 21103 26893 21116
rect 23048 21069 23151 21103
rect 23185 21069 23551 21103
rect 23585 21069 23951 21103
rect 23985 21069 24351 21103
rect 24385 21069 24751 21103
rect 24785 21069 25151 21103
rect 25185 21069 25551 21103
rect 25585 21069 25951 21103
rect 25985 21069 26351 21103
rect 26385 21069 26751 21103
rect 26785 21097 26893 21103
rect 26927 21097 27148 21116
rect 26785 21069 27148 21097
rect 23048 21056 27148 21069
rect 28286 21114 38954 21147
rect 28286 21080 28416 21114
rect 28450 21080 28506 21114
rect 28540 21080 28596 21114
rect 28630 21080 28686 21114
rect 28720 21080 28776 21114
rect 28810 21080 28866 21114
rect 28900 21080 28956 21114
rect 28990 21080 29046 21114
rect 29080 21080 29136 21114
rect 29170 21080 29226 21114
rect 29260 21080 29316 21114
rect 29350 21080 29406 21114
rect 29440 21080 29756 21114
rect 29790 21080 29846 21114
rect 29880 21080 29936 21114
rect 29970 21080 30026 21114
rect 30060 21080 30116 21114
rect 30150 21080 30206 21114
rect 30240 21080 30296 21114
rect 30330 21080 30386 21114
rect 30420 21080 30476 21114
rect 30510 21080 30566 21114
rect 30600 21080 30656 21114
rect 30690 21080 30746 21114
rect 30780 21080 31096 21114
rect 31130 21080 31186 21114
rect 31220 21080 31276 21114
rect 31310 21080 31366 21114
rect 31400 21080 31456 21114
rect 31490 21080 31546 21114
rect 31580 21080 31636 21114
rect 31670 21080 31726 21114
rect 31760 21080 31816 21114
rect 31850 21080 31906 21114
rect 31940 21080 31996 21114
rect 32030 21080 32086 21114
rect 32120 21080 32436 21114
rect 32470 21080 32526 21114
rect 32560 21080 32616 21114
rect 32650 21080 32706 21114
rect 32740 21080 32796 21114
rect 32830 21080 32886 21114
rect 32920 21080 32976 21114
rect 33010 21080 33066 21114
rect 33100 21080 33156 21114
rect 33190 21080 33246 21114
rect 33280 21080 33336 21114
rect 33370 21080 33426 21114
rect 33460 21080 33776 21114
rect 33810 21080 33866 21114
rect 33900 21080 33956 21114
rect 33990 21080 34046 21114
rect 34080 21080 34136 21114
rect 34170 21080 34226 21114
rect 34260 21080 34316 21114
rect 34350 21080 34406 21114
rect 34440 21080 34496 21114
rect 34530 21080 34586 21114
rect 34620 21080 34676 21114
rect 34710 21080 34766 21114
rect 34800 21080 35116 21114
rect 35150 21080 35206 21114
rect 35240 21080 35296 21114
rect 35330 21080 35386 21114
rect 35420 21080 35476 21114
rect 35510 21080 35566 21114
rect 35600 21080 35656 21114
rect 35690 21080 35746 21114
rect 35780 21080 35836 21114
rect 35870 21080 35926 21114
rect 35960 21080 36016 21114
rect 36050 21080 36106 21114
rect 36140 21080 36456 21114
rect 36490 21080 36546 21114
rect 36580 21080 36636 21114
rect 36670 21080 36726 21114
rect 36760 21080 36816 21114
rect 36850 21080 36906 21114
rect 36940 21080 36996 21114
rect 37030 21080 37086 21114
rect 37120 21080 37176 21114
rect 37210 21080 37266 21114
rect 37300 21080 37356 21114
rect 37390 21080 37446 21114
rect 37480 21080 37796 21114
rect 37830 21080 37886 21114
rect 37920 21080 37976 21114
rect 38010 21080 38066 21114
rect 38100 21080 38156 21114
rect 38190 21080 38246 21114
rect 38280 21080 38336 21114
rect 38370 21080 38426 21114
rect 38460 21080 38516 21114
rect 38550 21080 38606 21114
rect 38640 21080 38696 21114
rect 38730 21080 38786 21114
rect 38820 21080 38954 21114
rect 28286 21048 38954 21080
rect 7680 20995 13304 21022
rect 7680 20962 13277 20995
rect 7680 20903 8309 20916
rect 7680 20869 7863 20903
rect 7897 20869 8263 20903
rect 8297 20893 8309 20903
rect 8343 20903 13304 20916
rect 8343 20893 8663 20903
rect 8297 20869 8663 20893
rect 8697 20869 9063 20903
rect 9097 20869 9463 20903
rect 9497 20869 9863 20903
rect 9897 20869 10263 20903
rect 10297 20869 10663 20903
rect 10697 20869 11063 20903
rect 11097 20869 11463 20903
rect 11497 20869 11863 20903
rect 11897 20869 12263 20903
rect 12297 20869 12663 20903
rect 12697 20869 13063 20903
rect 13097 20869 13304 20903
rect 7680 20856 13304 20869
rect 22898 20909 22958 20992
rect 22898 20875 22911 20909
rect 22945 20875 22958 20909
rect 22898 20782 22958 20875
rect 23948 20879 24108 20902
rect 23948 20845 24013 20879
rect 24047 20845 24108 20879
rect 23948 20782 24108 20845
rect 25248 20879 25408 20902
rect 25248 20845 25313 20879
rect 25347 20845 25408 20879
rect 25248 20782 25408 20845
rect 40658 20782 41274 21581
rect 41754 21437 42186 21827
rect 7582 20769 13304 20782
rect 7582 20735 7863 20769
rect 7897 20735 8263 20769
rect 8297 20735 8663 20769
rect 8697 20735 9063 20769
rect 9097 20735 9463 20769
rect 9497 20735 9863 20769
rect 9897 20735 10263 20769
rect 10297 20735 10663 20769
rect 10697 20735 11063 20769
rect 11097 20735 11463 20769
rect 11497 20735 11863 20769
rect 11897 20735 12263 20769
rect 12297 20735 12663 20769
rect 12697 20735 13063 20769
rect 13097 20735 13304 20769
rect 7582 20722 13304 20735
rect 13562 20769 20730 20782
rect 13562 20735 13745 20769
rect 13779 20735 14145 20769
rect 14179 20735 14545 20769
rect 14579 20735 14945 20769
rect 14979 20735 15345 20769
rect 15379 20735 15745 20769
rect 15779 20735 16145 20769
rect 16179 20735 16545 20769
rect 16579 20735 16945 20769
rect 16979 20735 17345 20769
rect 17379 20735 17745 20769
rect 17779 20735 18145 20769
rect 18179 20735 18545 20769
rect 18579 20735 18945 20769
rect 18979 20735 19345 20769
rect 19379 20735 19745 20769
rect 19779 20735 20145 20769
rect 20179 20735 20545 20769
rect 20579 20735 20730 20769
rect 13562 20722 20730 20735
rect 21008 20769 22348 20782
rect 21008 20735 21191 20769
rect 21225 20735 21391 20769
rect 21425 20735 21591 20769
rect 21625 20735 21791 20769
rect 21825 20735 21991 20769
rect 22025 20735 22191 20769
rect 22225 20735 22348 20769
rect 21008 20722 22348 20735
rect 22870 20769 27148 20782
rect 22870 20735 23151 20769
rect 23185 20735 23551 20769
rect 23585 20735 23951 20769
rect 23985 20735 24351 20769
rect 24385 20735 24751 20769
rect 24785 20735 25151 20769
rect 25185 20735 25551 20769
rect 25585 20735 25951 20769
rect 25985 20735 26351 20769
rect 26385 20735 26751 20769
rect 26785 20735 27148 20769
rect 22870 20722 27148 20735
rect 28260 20769 38980 20782
rect 28260 20735 28443 20769
rect 28477 20735 28643 20769
rect 28677 20735 28843 20769
rect 28877 20735 29043 20769
rect 29077 20735 29243 20769
rect 29277 20735 29443 20769
rect 29477 20735 29643 20769
rect 29677 20735 29843 20769
rect 29877 20735 30043 20769
rect 30077 20735 30243 20769
rect 30277 20735 30443 20769
rect 30477 20735 30643 20769
rect 30677 20735 30843 20769
rect 30877 20735 31043 20769
rect 31077 20735 31243 20769
rect 31277 20735 31443 20769
rect 31477 20735 31643 20769
rect 31677 20735 31843 20769
rect 31877 20735 32043 20769
rect 32077 20735 32243 20769
rect 32277 20735 32443 20769
rect 32477 20735 32643 20769
rect 32677 20735 32843 20769
rect 32877 20735 33043 20769
rect 33077 20735 33243 20769
rect 33277 20735 33443 20769
rect 33477 20735 33643 20769
rect 33677 20735 33843 20769
rect 33877 20735 34043 20769
rect 34077 20735 34243 20769
rect 34277 20735 34443 20769
rect 34477 20735 34643 20769
rect 34677 20735 34843 20769
rect 34877 20735 35043 20769
rect 35077 20735 35243 20769
rect 35277 20735 35443 20769
rect 35477 20735 35643 20769
rect 35677 20735 35843 20769
rect 35877 20735 36043 20769
rect 36077 20735 36243 20769
rect 36277 20735 36443 20769
rect 36477 20735 36643 20769
rect 36677 20735 36843 20769
rect 36877 20735 37043 20769
rect 37077 20735 37243 20769
rect 37277 20735 37443 20769
rect 37477 20735 37643 20769
rect 37677 20735 37843 20769
rect 37877 20735 38043 20769
rect 38077 20735 38243 20769
rect 38277 20735 38443 20769
rect 38477 20735 38643 20769
rect 38677 20735 38843 20769
rect 38877 20735 38980 20769
rect 28260 20722 38980 20735
rect 39746 20769 42186 20782
rect 39746 20735 39929 20769
rect 39963 20735 40129 20769
rect 40163 20735 40329 20769
rect 40363 20735 40529 20769
rect 40563 20735 40729 20769
rect 40763 20735 40929 20769
rect 40963 20735 41129 20769
rect 41163 20735 41329 20769
rect 41363 20735 41529 20769
rect 41563 20735 41729 20769
rect 41763 20735 41929 20769
rect 41963 20735 42186 20769
rect 39746 20722 42186 20735
rect 5916 18889 10194 18902
rect 5916 18855 6197 18889
rect 6231 18855 6597 18889
rect 6631 18855 6997 18889
rect 7031 18855 7397 18889
rect 7431 18855 7797 18889
rect 7831 18855 8197 18889
rect 8231 18855 8597 18889
rect 8631 18855 8997 18889
rect 9031 18855 9397 18889
rect 9431 18855 9797 18889
rect 9831 18855 10194 18889
rect 5916 18842 10194 18855
rect 10640 18889 13080 18902
rect 10640 18855 10823 18889
rect 10857 18855 11023 18889
rect 11057 18855 11223 18889
rect 11257 18855 11423 18889
rect 11457 18855 11623 18889
rect 11657 18855 11823 18889
rect 11857 18855 12023 18889
rect 12057 18855 12223 18889
rect 12257 18855 12423 18889
rect 12457 18855 12623 18889
rect 12657 18855 12823 18889
rect 12857 18855 13080 18889
rect 10640 18842 13080 18855
rect 13384 18889 15824 18902
rect 13384 18855 13567 18889
rect 13601 18855 13767 18889
rect 13801 18855 13967 18889
rect 14001 18855 14167 18889
rect 14201 18855 14367 18889
rect 14401 18855 14567 18889
rect 14601 18855 14767 18889
rect 14801 18855 14967 18889
rect 15001 18855 15167 18889
rect 15201 18855 15367 18889
rect 15401 18855 15567 18889
rect 15601 18855 15824 18889
rect 13384 18842 15824 18855
rect 16110 18889 23278 18902
rect 16110 18855 16293 18889
rect 16327 18855 16693 18889
rect 16727 18855 17093 18889
rect 17127 18855 17493 18889
rect 17527 18855 17893 18889
rect 17927 18855 18293 18889
rect 18327 18855 18693 18889
rect 18727 18855 19093 18889
rect 19127 18855 19493 18889
rect 19527 18855 19893 18889
rect 19927 18855 20293 18889
rect 20327 18855 20693 18889
rect 20727 18855 21093 18889
rect 21127 18855 21493 18889
rect 21527 18855 21893 18889
rect 21927 18855 22293 18889
rect 22327 18855 22693 18889
rect 22727 18855 23093 18889
rect 23127 18855 23278 18889
rect 16110 18842 23278 18855
rect 23850 18889 26824 18902
rect 23850 18855 24131 18889
rect 24165 18855 24531 18889
rect 24565 18855 24931 18889
rect 24965 18855 25331 18889
rect 25365 18855 25731 18889
rect 25765 18855 26131 18889
rect 26165 18855 26531 18889
rect 26565 18855 26824 18889
rect 23850 18842 26824 18855
rect 28260 18889 38980 18902
rect 28260 18855 28443 18889
rect 28477 18855 28643 18889
rect 28677 18855 28843 18889
rect 28877 18855 29043 18889
rect 29077 18855 29243 18889
rect 29277 18855 29443 18889
rect 29477 18855 29643 18889
rect 29677 18855 29843 18889
rect 29877 18855 30043 18889
rect 30077 18855 30243 18889
rect 30277 18855 30443 18889
rect 30477 18855 30643 18889
rect 30677 18855 30843 18889
rect 30877 18855 31043 18889
rect 31077 18855 31243 18889
rect 31277 18855 31443 18889
rect 31477 18855 31643 18889
rect 31677 18855 31843 18889
rect 31877 18855 32043 18889
rect 32077 18855 32243 18889
rect 32277 18855 32443 18889
rect 32477 18855 32643 18889
rect 32677 18855 32843 18889
rect 32877 18855 33043 18889
rect 33077 18855 33243 18889
rect 33277 18855 33443 18889
rect 33477 18855 33643 18889
rect 33677 18855 33843 18889
rect 33877 18855 34043 18889
rect 34077 18855 34243 18889
rect 34277 18855 34443 18889
rect 34477 18855 34643 18889
rect 34677 18855 34843 18889
rect 34877 18855 35043 18889
rect 35077 18855 35243 18889
rect 35277 18855 35443 18889
rect 35477 18855 35643 18889
rect 35677 18855 35843 18889
rect 35877 18855 36043 18889
rect 36077 18855 36243 18889
rect 36277 18855 36443 18889
rect 36477 18855 36643 18889
rect 36677 18855 36843 18889
rect 36877 18855 37043 18889
rect 37077 18855 37243 18889
rect 37277 18855 37443 18889
rect 37477 18855 37643 18889
rect 37677 18855 37843 18889
rect 37877 18855 38043 18889
rect 38077 18855 38243 18889
rect 38277 18855 38443 18889
rect 38477 18855 38643 18889
rect 38677 18855 38843 18889
rect 38877 18855 38980 18889
rect 28260 18842 38980 18855
rect 39256 18889 41696 18902
rect 39256 18855 39439 18889
rect 39473 18855 39639 18889
rect 39673 18855 39839 18889
rect 39873 18855 40039 18889
rect 40073 18855 40239 18889
rect 40273 18855 40439 18889
rect 40473 18855 40639 18889
rect 40673 18855 40839 18889
rect 40873 18855 41039 18889
rect 41073 18855 41239 18889
rect 41273 18855 41439 18889
rect 41473 18855 41696 18889
rect 39256 18842 41696 18855
rect 23878 18749 23938 18842
rect 24926 18799 25086 18842
rect 24926 18765 24991 18799
rect 25025 18765 25086 18799
rect 24926 18762 25086 18765
rect 6014 18682 10194 18742
rect 23878 18715 23891 18749
rect 23925 18715 23938 18749
rect 6483 18396 6517 18682
rect 7399 18396 7433 18682
rect 8315 18396 8349 18682
rect 9231 18396 9265 18682
rect 10147 18396 10181 18682
rect 6026 18369 6060 18396
rect 6483 18378 6518 18396
rect 6026 18297 6060 18315
rect 6026 18225 6060 18247
rect 6026 18153 6060 18179
rect 6026 18081 6060 18111
rect 6026 18009 6060 18043
rect 6026 17941 6060 17975
rect 6026 17873 6060 17903
rect 6026 17805 6060 17831
rect 6026 17737 6060 17759
rect 6026 17669 6060 17687
rect 6025 17615 6026 17646
rect 6025 17588 6060 17615
rect 6484 18369 6518 18378
rect 6484 18297 6518 18315
rect 6484 18225 6518 18247
rect 6484 18153 6518 18179
rect 6484 18081 6518 18111
rect 6484 18009 6518 18043
rect 6484 17941 6518 17975
rect 6484 17873 6518 17903
rect 6484 17805 6518 17831
rect 6484 17737 6518 17759
rect 6484 17669 6518 17687
rect 6942 18369 6976 18396
rect 7399 18378 7434 18396
rect 6942 18297 6976 18315
rect 6942 18225 6976 18247
rect 6942 18153 6976 18179
rect 6942 18081 6976 18111
rect 6942 18009 6976 18043
rect 6942 17941 6976 17975
rect 6942 17873 6976 17903
rect 6942 17805 6976 17831
rect 6942 17737 6976 17759
rect 6942 17669 6976 17687
rect 6484 17588 6518 17615
rect 6941 17615 6942 17646
rect 6941 17588 6976 17615
rect 7400 18369 7434 18378
rect 7400 18297 7434 18315
rect 7400 18225 7434 18247
rect 7400 18153 7434 18179
rect 7400 18081 7434 18111
rect 7400 18009 7434 18043
rect 7400 17941 7434 17975
rect 7400 17873 7434 17903
rect 7400 17805 7434 17831
rect 7400 17737 7434 17759
rect 7400 17669 7434 17687
rect 7858 18369 7892 18396
rect 8315 18378 8350 18396
rect 7858 18297 7892 18315
rect 7858 18225 7892 18247
rect 7858 18153 7892 18179
rect 7858 18081 7892 18111
rect 7858 18009 7892 18043
rect 7858 17941 7892 17975
rect 7858 17873 7892 17903
rect 7858 17805 7892 17831
rect 7858 17737 7892 17759
rect 7858 17669 7892 17687
rect 7400 17588 7434 17615
rect 7857 17615 7858 17646
rect 7857 17588 7892 17615
rect 8316 18369 8350 18378
rect 8316 18297 8350 18315
rect 8316 18225 8350 18247
rect 8316 18153 8350 18179
rect 8316 18081 8350 18111
rect 8316 18009 8350 18043
rect 8316 17941 8350 17975
rect 8316 17873 8350 17903
rect 8316 17805 8350 17831
rect 8316 17737 8350 17759
rect 8316 17669 8350 17687
rect 8774 18369 8808 18396
rect 9231 18378 9266 18396
rect 8774 18297 8808 18315
rect 8774 18225 8808 18247
rect 8774 18153 8808 18179
rect 8774 18081 8808 18111
rect 8774 18009 8808 18043
rect 8774 17941 8808 17975
rect 8774 17873 8808 17903
rect 8774 17805 8808 17831
rect 8774 17737 8808 17759
rect 8774 17669 8808 17687
rect 8316 17588 8350 17615
rect 8773 17615 8774 17646
rect 8773 17588 8808 17615
rect 9232 18369 9266 18378
rect 9232 18297 9266 18315
rect 9232 18225 9266 18247
rect 9232 18153 9266 18179
rect 9232 18081 9266 18111
rect 9232 18009 9266 18043
rect 9232 17941 9266 17975
rect 9232 17873 9266 17903
rect 9232 17805 9266 17831
rect 9232 17737 9266 17759
rect 9232 17669 9266 17687
rect 9690 18369 9724 18396
rect 10147 18378 10182 18396
rect 9690 18297 9724 18315
rect 9690 18225 9724 18247
rect 9690 18153 9724 18179
rect 9690 18081 9724 18111
rect 9690 18009 9724 18043
rect 9690 17941 9724 17975
rect 9690 17873 9724 17903
rect 9690 17805 9724 17831
rect 9690 17737 9724 17759
rect 9690 17669 9724 17687
rect 9232 17588 9266 17615
rect 9689 17615 9690 17646
rect 9689 17588 9724 17615
rect 10148 18369 10182 18378
rect 10148 18297 10182 18315
rect 10148 18225 10182 18247
rect 10148 18153 10182 18179
rect 10148 18081 10182 18111
rect 23878 18632 23938 18715
rect 24008 18717 26824 18722
rect 24008 18683 26157 18717
rect 26191 18683 26824 18717
rect 24008 18682 26824 18683
rect 10148 18009 10182 18043
rect 10148 17941 10182 17975
rect 10148 17873 10182 17903
rect 10148 17805 10182 17831
rect 10148 17737 10182 17759
rect 10148 17669 10182 17687
rect 11552 17923 12168 17962
rect 11552 17821 11639 17923
rect 12081 17821 12168 17923
rect 10148 17588 10182 17615
rect 6025 17522 6059 17588
rect 6941 17522 6975 17588
rect 7857 17522 7891 17588
rect 8773 17522 8807 17588
rect 9689 17522 9723 17588
rect 6014 17462 10194 17522
rect 6094 17343 10194 17356
rect 6094 17323 6197 17343
rect 6094 17296 6101 17323
rect 6135 17309 6197 17323
rect 6231 17309 6597 17343
rect 6631 17309 6997 17343
rect 7031 17309 7397 17343
rect 7431 17309 7797 17343
rect 7831 17309 8197 17343
rect 8231 17309 8597 17343
rect 8631 17309 8997 17343
rect 9031 17309 9397 17343
rect 9431 17309 9797 17343
rect 9831 17309 10194 17343
rect 6135 17296 10194 17309
rect 5944 17149 6004 17232
rect 5944 17115 5957 17149
rect 5991 17115 6004 17149
rect 5944 17022 6004 17115
rect 6994 17119 7154 17142
rect 6994 17085 7059 17119
rect 7093 17085 7154 17119
rect 6994 17022 7154 17085
rect 8294 17119 8454 17142
rect 8294 17085 8359 17119
rect 8393 17085 8454 17119
rect 8294 17022 8454 17085
rect 11552 17022 12168 17821
rect 12648 17677 13080 18067
rect 14296 17923 14912 17962
rect 14296 17821 14383 17923
rect 14825 17821 14912 17923
rect 14296 17022 14912 17821
rect 15392 17677 15824 18067
rect 23995 18621 24029 18641
rect 23995 18553 24029 18587
rect 23995 18485 24029 18515
rect 23995 18417 24029 18443
rect 23995 18349 24029 18371
rect 23995 18281 24029 18299
rect 23995 18213 24029 18227
rect 23995 18145 24029 18155
rect 23995 18077 24029 18083
rect 23995 18009 24029 18011
rect 23995 17973 24029 17975
rect 23995 17901 24029 17907
rect 23995 17829 24029 17839
rect 23995 17757 24029 17771
rect 23995 17685 24029 17703
rect 23995 17613 24029 17635
rect 23995 17541 24029 17567
rect 23995 17469 24029 17499
rect 23995 17397 24029 17431
rect 23995 17262 24029 17363
rect 24453 18621 24487 18682
rect 24453 18553 24487 18587
rect 24453 18485 24487 18515
rect 24453 18417 24487 18443
rect 24453 18349 24487 18371
rect 24453 18281 24487 18299
rect 24453 18213 24487 18227
rect 24453 18145 24487 18155
rect 24453 18077 24487 18083
rect 24453 18009 24487 18011
rect 24453 17973 24487 17975
rect 24453 17901 24487 17907
rect 24453 17829 24487 17839
rect 24453 17757 24487 17771
rect 24453 17685 24487 17703
rect 24453 17613 24487 17635
rect 24453 17541 24487 17567
rect 24453 17469 24487 17499
rect 24453 17397 24487 17431
rect 24453 17343 24487 17363
rect 24911 18621 24945 18641
rect 24911 18553 24945 18587
rect 24911 18485 24945 18515
rect 24911 18417 24945 18443
rect 24911 18349 24945 18371
rect 24911 18281 24945 18299
rect 24911 18213 24945 18227
rect 24911 18145 24945 18155
rect 24911 18077 24945 18083
rect 24911 18009 24945 18011
rect 24911 17973 24945 17975
rect 24911 17901 24945 17907
rect 24911 17829 24945 17839
rect 24911 17757 24945 17771
rect 24911 17685 24945 17703
rect 24911 17613 24945 17635
rect 24911 17541 24945 17567
rect 24911 17469 24945 17499
rect 24911 17397 24945 17431
rect 24911 17262 24945 17363
rect 25369 18621 25403 18682
rect 25369 18553 25403 18587
rect 25369 18485 25403 18515
rect 25369 18417 25403 18443
rect 25369 18349 25403 18371
rect 25369 18281 25403 18299
rect 25369 18213 25403 18227
rect 25369 18145 25403 18155
rect 25369 18077 25403 18083
rect 25369 18009 25403 18011
rect 25369 17973 25403 17975
rect 25369 17901 25403 17907
rect 25369 17829 25403 17839
rect 25369 17757 25403 17771
rect 25369 17685 25403 17703
rect 25369 17613 25403 17635
rect 25369 17541 25403 17567
rect 25369 17469 25403 17499
rect 25369 17397 25403 17431
rect 25369 17343 25403 17363
rect 25827 18621 25861 18641
rect 25827 18553 25861 18587
rect 25827 18485 25861 18515
rect 25827 18417 25861 18443
rect 25827 18349 25861 18371
rect 25827 18281 25861 18299
rect 25827 18213 25861 18227
rect 25827 18145 25861 18155
rect 25827 18077 25861 18083
rect 25827 18009 25861 18011
rect 25827 17973 25861 17975
rect 25827 17901 25861 17907
rect 25827 17829 25861 17839
rect 25827 17757 25861 17771
rect 25827 17685 25861 17703
rect 25827 17613 25861 17635
rect 25827 17541 25861 17567
rect 25827 17469 25861 17499
rect 25827 17397 25861 17431
rect 25827 17262 25861 17363
rect 26285 18621 26319 18682
rect 26285 18553 26319 18587
rect 26285 18485 26319 18515
rect 26285 18417 26319 18443
rect 26285 18349 26319 18371
rect 26285 18281 26319 18299
rect 26285 18213 26319 18227
rect 26285 18145 26319 18155
rect 26285 18077 26319 18083
rect 26285 18009 26319 18011
rect 26285 17973 26319 17975
rect 26285 17901 26319 17907
rect 26285 17829 26319 17839
rect 26285 17757 26319 17771
rect 26285 17685 26319 17703
rect 26285 17613 26319 17635
rect 26285 17541 26319 17567
rect 26285 17469 26319 17499
rect 26285 17397 26319 17431
rect 26285 17343 26319 17363
rect 26743 18621 26777 18641
rect 26743 18553 26777 18587
rect 26743 18485 26777 18515
rect 26743 18417 26777 18443
rect 26743 18349 26777 18371
rect 26743 18281 26777 18299
rect 26743 18213 26777 18227
rect 26743 18145 26777 18155
rect 26743 18077 26777 18083
rect 26743 18009 26777 18011
rect 26743 17973 26777 17975
rect 26743 17901 26777 17907
rect 26743 17829 26777 17839
rect 26743 17757 26777 17771
rect 26743 17685 26777 17703
rect 26743 17613 26777 17635
rect 26743 17541 26777 17567
rect 26743 17469 26777 17499
rect 26743 17397 26777 17431
rect 26743 17262 26777 17363
rect 28286 18556 38954 18576
rect 28286 18522 28306 18556
rect 28340 18522 28396 18556
rect 28430 18541 28486 18556
rect 28520 18541 28576 18556
rect 28610 18541 28666 18556
rect 28700 18541 28756 18556
rect 28790 18541 28846 18556
rect 28880 18541 28936 18556
rect 28970 18541 29026 18556
rect 29060 18541 29116 18556
rect 29150 18541 29206 18556
rect 29240 18541 29296 18556
rect 29330 18541 29386 18556
rect 29420 18541 29476 18556
rect 28450 18522 28486 18541
rect 28540 18522 28576 18541
rect 28630 18522 28666 18541
rect 28720 18522 28756 18541
rect 28810 18522 28846 18541
rect 28900 18522 28936 18541
rect 28990 18522 29026 18541
rect 29080 18522 29116 18541
rect 29170 18522 29206 18541
rect 29260 18522 29296 18541
rect 29350 18522 29386 18541
rect 29440 18522 29476 18541
rect 29510 18522 29646 18556
rect 29680 18522 29736 18556
rect 29770 18541 29826 18556
rect 29860 18541 29916 18556
rect 29950 18541 30006 18556
rect 30040 18541 30096 18556
rect 30130 18541 30186 18556
rect 30220 18541 30276 18556
rect 30310 18541 30366 18556
rect 30400 18541 30456 18556
rect 30490 18541 30546 18556
rect 30580 18541 30636 18556
rect 30670 18541 30726 18556
rect 30760 18541 30816 18556
rect 29790 18522 29826 18541
rect 29880 18522 29916 18541
rect 29970 18522 30006 18541
rect 30060 18522 30096 18541
rect 30150 18522 30186 18541
rect 30240 18522 30276 18541
rect 30330 18522 30366 18541
rect 30420 18522 30456 18541
rect 30510 18522 30546 18541
rect 30600 18522 30636 18541
rect 30690 18522 30726 18541
rect 30780 18522 30816 18541
rect 30850 18522 30986 18556
rect 31020 18522 31076 18556
rect 31110 18541 31166 18556
rect 31200 18541 31256 18556
rect 31290 18541 31346 18556
rect 31380 18541 31436 18556
rect 31470 18541 31526 18556
rect 31560 18541 31616 18556
rect 31650 18541 31706 18556
rect 31740 18541 31796 18556
rect 31830 18541 31886 18556
rect 31920 18541 31976 18556
rect 32010 18541 32066 18556
rect 32100 18541 32156 18556
rect 31130 18522 31166 18541
rect 31220 18522 31256 18541
rect 31310 18522 31346 18541
rect 31400 18522 31436 18541
rect 31490 18522 31526 18541
rect 31580 18522 31616 18541
rect 31670 18522 31706 18541
rect 31760 18522 31796 18541
rect 31850 18522 31886 18541
rect 31940 18522 31976 18541
rect 32030 18522 32066 18541
rect 32120 18522 32156 18541
rect 32190 18522 32326 18556
rect 32360 18522 32416 18556
rect 32450 18541 32506 18556
rect 32540 18541 32596 18556
rect 32630 18541 32686 18556
rect 32720 18541 32776 18556
rect 32810 18541 32866 18556
rect 32900 18541 32956 18556
rect 32990 18541 33046 18556
rect 33080 18541 33136 18556
rect 33170 18541 33226 18556
rect 33260 18541 33316 18556
rect 33350 18541 33406 18556
rect 33440 18541 33496 18556
rect 32470 18522 32506 18541
rect 32560 18522 32596 18541
rect 32650 18522 32686 18541
rect 32740 18522 32776 18541
rect 32830 18522 32866 18541
rect 32920 18522 32956 18541
rect 33010 18522 33046 18541
rect 33100 18522 33136 18541
rect 33190 18522 33226 18541
rect 33280 18522 33316 18541
rect 33370 18522 33406 18541
rect 33460 18522 33496 18541
rect 33530 18522 33666 18556
rect 33700 18522 33756 18556
rect 33790 18541 33846 18556
rect 33880 18541 33936 18556
rect 33970 18541 34026 18556
rect 34060 18541 34116 18556
rect 34150 18541 34206 18556
rect 34240 18541 34296 18556
rect 34330 18541 34386 18556
rect 34420 18541 34476 18556
rect 34510 18541 34566 18556
rect 34600 18541 34656 18556
rect 34690 18541 34746 18556
rect 34780 18541 34836 18556
rect 33810 18522 33846 18541
rect 33900 18522 33936 18541
rect 33990 18522 34026 18541
rect 34080 18522 34116 18541
rect 34170 18522 34206 18541
rect 34260 18522 34296 18541
rect 34350 18522 34386 18541
rect 34440 18522 34476 18541
rect 34530 18522 34566 18541
rect 34620 18522 34656 18541
rect 34710 18522 34746 18541
rect 34800 18522 34836 18541
rect 34870 18522 35006 18556
rect 35040 18522 35096 18556
rect 35130 18541 35186 18556
rect 35220 18541 35276 18556
rect 35310 18541 35366 18556
rect 35400 18541 35456 18556
rect 35490 18541 35546 18556
rect 35580 18541 35636 18556
rect 35670 18541 35726 18556
rect 35760 18541 35816 18556
rect 35850 18541 35906 18556
rect 35940 18541 35996 18556
rect 36030 18541 36086 18556
rect 36120 18541 36176 18556
rect 35150 18522 35186 18541
rect 35240 18522 35276 18541
rect 35330 18522 35366 18541
rect 35420 18522 35456 18541
rect 35510 18522 35546 18541
rect 35600 18522 35636 18541
rect 35690 18522 35726 18541
rect 35780 18522 35816 18541
rect 35870 18522 35906 18541
rect 35960 18522 35996 18541
rect 36050 18522 36086 18541
rect 36140 18522 36176 18541
rect 36210 18522 36346 18556
rect 36380 18522 36436 18556
rect 36470 18541 36526 18556
rect 36560 18541 36616 18556
rect 36650 18541 36706 18556
rect 36740 18541 36796 18556
rect 36830 18541 36886 18556
rect 36920 18541 36976 18556
rect 37010 18541 37066 18556
rect 37100 18541 37156 18556
rect 37190 18541 37246 18556
rect 37280 18541 37336 18556
rect 37370 18541 37426 18556
rect 37460 18541 37516 18556
rect 36490 18522 36526 18541
rect 36580 18522 36616 18541
rect 36670 18522 36706 18541
rect 36760 18522 36796 18541
rect 36850 18522 36886 18541
rect 36940 18522 36976 18541
rect 37030 18522 37066 18541
rect 37120 18522 37156 18541
rect 37210 18522 37246 18541
rect 37300 18522 37336 18541
rect 37390 18522 37426 18541
rect 37480 18522 37516 18541
rect 37550 18522 37686 18556
rect 37720 18522 37776 18556
rect 37810 18541 37866 18556
rect 37900 18541 37956 18556
rect 37990 18541 38046 18556
rect 38080 18541 38136 18556
rect 38170 18541 38226 18556
rect 38260 18541 38316 18556
rect 38350 18541 38406 18556
rect 38440 18541 38496 18556
rect 38530 18541 38586 18556
rect 38620 18541 38676 18556
rect 38710 18541 38766 18556
rect 38800 18541 38856 18556
rect 37830 18522 37866 18541
rect 37920 18522 37956 18541
rect 38010 18522 38046 18541
rect 38100 18522 38136 18541
rect 38190 18522 38226 18541
rect 38280 18522 38316 18541
rect 38370 18522 38406 18541
rect 38460 18522 38496 18541
rect 38550 18522 38586 18541
rect 38640 18522 38676 18541
rect 38730 18522 38766 18541
rect 38820 18522 38856 18541
rect 38890 18522 38954 18556
rect 28286 18518 28416 18522
rect 28286 18484 28320 18518
rect 28354 18507 28416 18518
rect 28450 18507 28506 18522
rect 28540 18507 28596 18522
rect 28630 18507 28686 18522
rect 28720 18507 28776 18522
rect 28810 18507 28866 18522
rect 28900 18507 28956 18522
rect 28990 18507 29046 18522
rect 29080 18507 29136 18522
rect 29170 18507 29226 18522
rect 29260 18507 29316 18522
rect 29350 18507 29406 18522
rect 29440 18518 29756 18522
rect 29440 18507 29507 18518
rect 28354 18484 29507 18507
rect 29541 18484 29660 18518
rect 29694 18507 29756 18518
rect 29790 18507 29846 18522
rect 29880 18507 29936 18522
rect 29970 18507 30026 18522
rect 30060 18507 30116 18522
rect 30150 18507 30206 18522
rect 30240 18507 30296 18522
rect 30330 18507 30386 18522
rect 30420 18507 30476 18522
rect 30510 18507 30566 18522
rect 30600 18507 30656 18522
rect 30690 18507 30746 18522
rect 30780 18518 31096 18522
rect 30780 18507 30847 18518
rect 29694 18484 30847 18507
rect 30881 18484 31000 18518
rect 31034 18507 31096 18518
rect 31130 18507 31186 18522
rect 31220 18507 31276 18522
rect 31310 18507 31366 18522
rect 31400 18507 31456 18522
rect 31490 18507 31546 18522
rect 31580 18507 31636 18522
rect 31670 18507 31726 18522
rect 31760 18507 31816 18522
rect 31850 18507 31906 18522
rect 31940 18507 31996 18522
rect 32030 18507 32086 18522
rect 32120 18518 32436 18522
rect 32120 18507 32187 18518
rect 31034 18484 32187 18507
rect 32221 18484 32340 18518
rect 32374 18507 32436 18518
rect 32470 18507 32526 18522
rect 32560 18507 32616 18522
rect 32650 18507 32706 18522
rect 32740 18507 32796 18522
rect 32830 18507 32886 18522
rect 32920 18507 32976 18522
rect 33010 18507 33066 18522
rect 33100 18507 33156 18522
rect 33190 18507 33246 18522
rect 33280 18507 33336 18522
rect 33370 18507 33426 18522
rect 33460 18518 33776 18522
rect 33460 18507 33527 18518
rect 32374 18484 33527 18507
rect 33561 18484 33680 18518
rect 33714 18507 33776 18518
rect 33810 18507 33866 18522
rect 33900 18507 33956 18522
rect 33990 18507 34046 18522
rect 34080 18507 34136 18522
rect 34170 18507 34226 18522
rect 34260 18507 34316 18522
rect 34350 18507 34406 18522
rect 34440 18507 34496 18522
rect 34530 18507 34586 18522
rect 34620 18507 34676 18522
rect 34710 18507 34766 18522
rect 34800 18518 35116 18522
rect 34800 18507 34867 18518
rect 33714 18484 34867 18507
rect 34901 18484 35020 18518
rect 35054 18507 35116 18518
rect 35150 18507 35206 18522
rect 35240 18507 35296 18522
rect 35330 18507 35386 18522
rect 35420 18507 35476 18522
rect 35510 18507 35566 18522
rect 35600 18507 35656 18522
rect 35690 18507 35746 18522
rect 35780 18507 35836 18522
rect 35870 18507 35926 18522
rect 35960 18507 36016 18522
rect 36050 18507 36106 18522
rect 36140 18518 36456 18522
rect 36140 18507 36207 18518
rect 35054 18484 36207 18507
rect 36241 18484 36360 18518
rect 36394 18507 36456 18518
rect 36490 18507 36546 18522
rect 36580 18507 36636 18522
rect 36670 18507 36726 18522
rect 36760 18507 36816 18522
rect 36850 18507 36906 18522
rect 36940 18507 36996 18522
rect 37030 18507 37086 18522
rect 37120 18507 37176 18522
rect 37210 18507 37266 18522
rect 37300 18507 37356 18522
rect 37390 18507 37446 18522
rect 37480 18518 37796 18522
rect 37480 18507 37547 18518
rect 36394 18484 37547 18507
rect 37581 18484 37700 18518
rect 37734 18507 37796 18518
rect 37830 18507 37886 18522
rect 37920 18507 37976 18522
rect 38010 18507 38066 18522
rect 38100 18507 38156 18522
rect 38190 18507 38246 18522
rect 38280 18507 38336 18522
rect 38370 18507 38426 18522
rect 38460 18507 38516 18522
rect 38550 18507 38606 18522
rect 38640 18507 38696 18522
rect 38730 18507 38786 18522
rect 38820 18518 38954 18522
rect 38820 18507 38887 18518
rect 37734 18484 38887 18507
rect 38921 18484 38954 18518
rect 28286 18477 38954 18484
rect 28286 18428 28385 18477
rect 28286 18394 28320 18428
rect 28354 18394 28385 18428
rect 29475 18428 29725 18477
rect 28286 18338 28385 18394
rect 28286 18304 28320 18338
rect 28354 18304 28385 18338
rect 28286 18248 28385 18304
rect 28286 18214 28320 18248
rect 28354 18214 28385 18248
rect 28286 18158 28385 18214
rect 28286 18124 28320 18158
rect 28354 18124 28385 18158
rect 28286 18068 28385 18124
rect 28286 18034 28320 18068
rect 28354 18034 28385 18068
rect 28286 17978 28385 18034
rect 28286 17944 28320 17978
rect 28354 17944 28385 17978
rect 28286 17888 28385 17944
rect 28286 17854 28320 17888
rect 28354 17854 28385 17888
rect 28286 17798 28385 17854
rect 28286 17764 28320 17798
rect 28354 17764 28385 17798
rect 28286 17708 28385 17764
rect 28286 17674 28320 17708
rect 28354 17674 28385 17708
rect 28286 17618 28385 17674
rect 28286 17584 28320 17618
rect 28354 17584 28385 17618
rect 28286 17528 28385 17584
rect 28286 17494 28320 17528
rect 28354 17494 28385 17528
rect 28286 17438 28385 17494
rect 28449 18396 29411 18413
rect 28449 18362 28470 18396
rect 28504 18362 28560 18396
rect 28594 18394 28650 18396
rect 28684 18394 28740 18396
rect 28774 18394 28830 18396
rect 28864 18394 28920 18396
rect 28954 18394 29010 18396
rect 29044 18394 29100 18396
rect 29134 18394 29190 18396
rect 29224 18394 29280 18396
rect 29314 18394 29370 18396
rect 28614 18362 28650 18394
rect 28704 18362 28740 18394
rect 28794 18362 28830 18394
rect 28884 18362 28920 18394
rect 28974 18362 29010 18394
rect 29064 18362 29100 18394
rect 29154 18362 29190 18394
rect 29244 18362 29280 18394
rect 29334 18362 29370 18394
rect 29404 18362 29411 18396
rect 28449 18360 28580 18362
rect 28614 18360 28670 18362
rect 28704 18360 28760 18362
rect 28794 18360 28850 18362
rect 28884 18360 28940 18362
rect 28974 18360 29030 18362
rect 29064 18360 29120 18362
rect 29154 18360 29210 18362
rect 29244 18360 29300 18362
rect 29334 18360 29411 18362
rect 28449 18341 29411 18360
rect 28449 18337 28521 18341
rect 28449 18303 28468 18337
rect 28502 18303 28521 18337
rect 28449 18247 28521 18303
rect 29339 18318 29411 18341
rect 29339 18284 29358 18318
rect 29392 18284 29411 18318
rect 28449 18213 28468 18247
rect 28502 18213 28521 18247
rect 28449 18157 28521 18213
rect 28449 18123 28468 18157
rect 28502 18123 28521 18157
rect 28449 18067 28521 18123
rect 28449 18033 28468 18067
rect 28502 18033 28521 18067
rect 28449 17977 28521 18033
rect 28449 17943 28468 17977
rect 28502 17943 28521 17977
rect 28449 17887 28521 17943
rect 28449 17853 28468 17887
rect 28502 17853 28521 17887
rect 28449 17797 28521 17853
rect 28449 17763 28468 17797
rect 28502 17763 28521 17797
rect 28449 17707 28521 17763
rect 28449 17673 28468 17707
rect 28502 17673 28521 17707
rect 28449 17617 28521 17673
rect 28449 17583 28468 17617
rect 28502 17583 28521 17617
rect 28583 18220 29277 18279
rect 28583 18186 28644 18220
rect 28678 18192 28734 18220
rect 28768 18192 28824 18220
rect 28858 18192 28914 18220
rect 28690 18186 28734 18192
rect 28790 18186 28824 18192
rect 28890 18186 28914 18192
rect 28948 18192 29004 18220
rect 28948 18186 28956 18192
rect 28583 18158 28656 18186
rect 28690 18158 28756 18186
rect 28790 18158 28856 18186
rect 28890 18158 28956 18186
rect 28990 18186 29004 18192
rect 29038 18192 29094 18220
rect 29038 18186 29056 18192
rect 28990 18158 29056 18186
rect 29090 18186 29094 18192
rect 29128 18192 29184 18220
rect 29128 18186 29156 18192
rect 29218 18186 29277 18220
rect 29090 18158 29156 18186
rect 29190 18158 29277 18186
rect 28583 18130 29277 18158
rect 28583 18096 28644 18130
rect 28678 18096 28734 18130
rect 28768 18096 28824 18130
rect 28858 18096 28914 18130
rect 28948 18096 29004 18130
rect 29038 18096 29094 18130
rect 29128 18096 29184 18130
rect 29218 18096 29277 18130
rect 28583 18092 29277 18096
rect 28583 18058 28656 18092
rect 28690 18058 28756 18092
rect 28790 18058 28856 18092
rect 28890 18058 28956 18092
rect 28990 18058 29056 18092
rect 29090 18058 29156 18092
rect 29190 18058 29277 18092
rect 28583 18040 29277 18058
rect 28583 18006 28644 18040
rect 28678 18006 28734 18040
rect 28768 18006 28824 18040
rect 28858 18006 28914 18040
rect 28948 18006 29004 18040
rect 29038 18006 29094 18040
rect 29128 18006 29184 18040
rect 29218 18006 29277 18040
rect 28583 17992 29277 18006
rect 28583 17958 28656 17992
rect 28690 17958 28756 17992
rect 28790 17958 28856 17992
rect 28890 17958 28956 17992
rect 28990 17958 29056 17992
rect 29090 17958 29156 17992
rect 29190 17958 29277 17992
rect 28583 17950 29277 17958
rect 28583 17916 28644 17950
rect 28678 17916 28734 17950
rect 28768 17916 28824 17950
rect 28858 17916 28914 17950
rect 28948 17916 29004 17950
rect 29038 17916 29094 17950
rect 29128 17916 29184 17950
rect 29218 17916 29277 17950
rect 28583 17892 29277 17916
rect 28583 17860 28656 17892
rect 28690 17860 28756 17892
rect 28790 17860 28856 17892
rect 28890 17860 28956 17892
rect 28583 17826 28644 17860
rect 28690 17858 28734 17860
rect 28790 17858 28824 17860
rect 28890 17858 28914 17860
rect 28678 17826 28734 17858
rect 28768 17826 28824 17858
rect 28858 17826 28914 17858
rect 28948 17858 28956 17860
rect 28990 17860 29056 17892
rect 28990 17858 29004 17860
rect 28948 17826 29004 17858
rect 29038 17858 29056 17860
rect 29090 17860 29156 17892
rect 29190 17860 29277 17892
rect 29090 17858 29094 17860
rect 29038 17826 29094 17858
rect 29128 17858 29156 17860
rect 29128 17826 29184 17858
rect 29218 17826 29277 17860
rect 28583 17792 29277 17826
rect 28583 17770 28656 17792
rect 28690 17770 28756 17792
rect 28790 17770 28856 17792
rect 28890 17770 28956 17792
rect 28583 17736 28644 17770
rect 28690 17758 28734 17770
rect 28790 17758 28824 17770
rect 28890 17758 28914 17770
rect 28678 17736 28734 17758
rect 28768 17736 28824 17758
rect 28858 17736 28914 17758
rect 28948 17758 28956 17770
rect 28990 17770 29056 17792
rect 28990 17758 29004 17770
rect 28948 17736 29004 17758
rect 29038 17758 29056 17770
rect 29090 17770 29156 17792
rect 29190 17770 29277 17792
rect 29090 17758 29094 17770
rect 29038 17736 29094 17758
rect 29128 17758 29156 17770
rect 29128 17736 29184 17758
rect 29218 17736 29277 17770
rect 28583 17692 29277 17736
rect 28583 17680 28656 17692
rect 28690 17680 28756 17692
rect 28790 17680 28856 17692
rect 28890 17680 28956 17692
rect 28583 17646 28644 17680
rect 28690 17658 28734 17680
rect 28790 17658 28824 17680
rect 28890 17658 28914 17680
rect 28678 17646 28734 17658
rect 28768 17646 28824 17658
rect 28858 17646 28914 17658
rect 28948 17658 28956 17680
rect 28990 17680 29056 17692
rect 28990 17658 29004 17680
rect 28948 17646 29004 17658
rect 29038 17658 29056 17680
rect 29090 17680 29156 17692
rect 29190 17680 29277 17692
rect 29090 17658 29094 17680
rect 29038 17646 29094 17658
rect 29128 17658 29156 17680
rect 29128 17646 29184 17658
rect 29218 17646 29277 17680
rect 28583 17585 29277 17646
rect 29339 18228 29411 18284
rect 29339 18194 29358 18228
rect 29392 18194 29411 18228
rect 29339 18138 29411 18194
rect 29339 18104 29358 18138
rect 29392 18104 29411 18138
rect 29339 18048 29411 18104
rect 29339 18014 29358 18048
rect 29392 18014 29411 18048
rect 29339 17958 29411 18014
rect 29339 17924 29358 17958
rect 29392 17924 29411 17958
rect 29339 17868 29411 17924
rect 29339 17834 29358 17868
rect 29392 17834 29411 17868
rect 29339 17778 29411 17834
rect 29339 17744 29358 17778
rect 29392 17744 29411 17778
rect 29339 17688 29411 17744
rect 29339 17654 29358 17688
rect 29392 17654 29411 17688
rect 29339 17598 29411 17654
rect 28449 17523 28521 17583
rect 29339 17564 29358 17598
rect 29392 17564 29411 17598
rect 29339 17523 29411 17564
rect 28449 17504 29411 17523
rect 28449 17470 28546 17504
rect 28580 17470 28636 17504
rect 28670 17470 28726 17504
rect 28760 17470 28816 17504
rect 28850 17470 28906 17504
rect 28940 17470 28996 17504
rect 29030 17470 29086 17504
rect 29120 17470 29176 17504
rect 29210 17470 29266 17504
rect 29300 17470 29411 17504
rect 28449 17451 29411 17470
rect 29475 18394 29507 18428
rect 29541 18394 29660 18428
rect 29694 18394 29725 18428
rect 30815 18428 31065 18477
rect 29475 18338 29725 18394
rect 29475 18304 29507 18338
rect 29541 18304 29660 18338
rect 29694 18304 29725 18338
rect 29475 18248 29725 18304
rect 29475 18214 29507 18248
rect 29541 18214 29660 18248
rect 29694 18214 29725 18248
rect 29475 18158 29725 18214
rect 29475 18124 29507 18158
rect 29541 18124 29660 18158
rect 29694 18124 29725 18158
rect 29475 18068 29725 18124
rect 29475 18034 29507 18068
rect 29541 18034 29660 18068
rect 29694 18034 29725 18068
rect 29475 17978 29725 18034
rect 29475 17944 29507 17978
rect 29541 17944 29660 17978
rect 29694 17944 29725 17978
rect 29475 17888 29725 17944
rect 29475 17854 29507 17888
rect 29541 17854 29660 17888
rect 29694 17854 29725 17888
rect 29475 17798 29725 17854
rect 29475 17764 29507 17798
rect 29541 17764 29660 17798
rect 29694 17764 29725 17798
rect 29475 17708 29725 17764
rect 29475 17674 29507 17708
rect 29541 17674 29660 17708
rect 29694 17674 29725 17708
rect 29475 17618 29725 17674
rect 29475 17584 29507 17618
rect 29541 17584 29660 17618
rect 29694 17584 29725 17618
rect 29475 17528 29725 17584
rect 29475 17494 29507 17528
rect 29541 17494 29660 17528
rect 29694 17494 29725 17528
rect 28286 17404 28320 17438
rect 28354 17404 28385 17438
rect 28286 17387 28385 17404
rect 29475 17438 29725 17494
rect 29789 18396 30751 18413
rect 29789 18362 29810 18396
rect 29844 18362 29900 18396
rect 29934 18394 29990 18396
rect 30024 18394 30080 18396
rect 30114 18394 30170 18396
rect 30204 18394 30260 18396
rect 30294 18394 30350 18396
rect 30384 18394 30440 18396
rect 30474 18394 30530 18396
rect 30564 18394 30620 18396
rect 30654 18394 30710 18396
rect 29954 18362 29990 18394
rect 30044 18362 30080 18394
rect 30134 18362 30170 18394
rect 30224 18362 30260 18394
rect 30314 18362 30350 18394
rect 30404 18362 30440 18394
rect 30494 18362 30530 18394
rect 30584 18362 30620 18394
rect 30674 18362 30710 18394
rect 30744 18362 30751 18396
rect 29789 18360 29920 18362
rect 29954 18360 30010 18362
rect 30044 18360 30100 18362
rect 30134 18360 30190 18362
rect 30224 18360 30280 18362
rect 30314 18360 30370 18362
rect 30404 18360 30460 18362
rect 30494 18360 30550 18362
rect 30584 18360 30640 18362
rect 30674 18360 30751 18362
rect 29789 18341 30751 18360
rect 29789 18337 29861 18341
rect 29789 18303 29808 18337
rect 29842 18303 29861 18337
rect 29789 18247 29861 18303
rect 30679 18318 30751 18341
rect 30679 18284 30698 18318
rect 30732 18284 30751 18318
rect 29789 18213 29808 18247
rect 29842 18213 29861 18247
rect 29789 18157 29861 18213
rect 29789 18123 29808 18157
rect 29842 18123 29861 18157
rect 29789 18067 29861 18123
rect 29789 18033 29808 18067
rect 29842 18033 29861 18067
rect 29789 17977 29861 18033
rect 29789 17943 29808 17977
rect 29842 17943 29861 17977
rect 29789 17887 29861 17943
rect 29789 17853 29808 17887
rect 29842 17853 29861 17887
rect 29789 17797 29861 17853
rect 29789 17763 29808 17797
rect 29842 17763 29861 17797
rect 29789 17707 29861 17763
rect 29789 17673 29808 17707
rect 29842 17673 29861 17707
rect 29789 17617 29861 17673
rect 29789 17583 29808 17617
rect 29842 17583 29861 17617
rect 29923 18220 30617 18279
rect 29923 18186 29984 18220
rect 30018 18192 30074 18220
rect 30108 18192 30164 18220
rect 30198 18192 30254 18220
rect 30030 18186 30074 18192
rect 30130 18186 30164 18192
rect 30230 18186 30254 18192
rect 30288 18192 30344 18220
rect 30288 18186 30296 18192
rect 29923 18158 29996 18186
rect 30030 18158 30096 18186
rect 30130 18158 30196 18186
rect 30230 18158 30296 18186
rect 30330 18186 30344 18192
rect 30378 18192 30434 18220
rect 30378 18186 30396 18192
rect 30330 18158 30396 18186
rect 30430 18186 30434 18192
rect 30468 18192 30524 18220
rect 30468 18186 30496 18192
rect 30558 18186 30617 18220
rect 30430 18158 30496 18186
rect 30530 18158 30617 18186
rect 29923 18130 30617 18158
rect 29923 18096 29984 18130
rect 30018 18096 30074 18130
rect 30108 18096 30164 18130
rect 30198 18096 30254 18130
rect 30288 18096 30344 18130
rect 30378 18096 30434 18130
rect 30468 18096 30524 18130
rect 30558 18096 30617 18130
rect 29923 18092 30617 18096
rect 29923 18058 29996 18092
rect 30030 18058 30096 18092
rect 30130 18058 30196 18092
rect 30230 18058 30296 18092
rect 30330 18058 30396 18092
rect 30430 18058 30496 18092
rect 30530 18058 30617 18092
rect 29923 18040 30617 18058
rect 29923 18006 29984 18040
rect 30018 18006 30074 18040
rect 30108 18006 30164 18040
rect 30198 18006 30254 18040
rect 30288 18006 30344 18040
rect 30378 18006 30434 18040
rect 30468 18006 30524 18040
rect 30558 18006 30617 18040
rect 29923 17992 30617 18006
rect 29923 17958 29996 17992
rect 30030 17958 30096 17992
rect 30130 17958 30196 17992
rect 30230 17958 30296 17992
rect 30330 17958 30396 17992
rect 30430 17958 30496 17992
rect 30530 17958 30617 17992
rect 29923 17950 30617 17958
rect 29923 17916 29984 17950
rect 30018 17916 30074 17950
rect 30108 17916 30164 17950
rect 30198 17916 30254 17950
rect 30288 17916 30344 17950
rect 30378 17916 30434 17950
rect 30468 17916 30524 17950
rect 30558 17916 30617 17950
rect 29923 17892 30617 17916
rect 29923 17860 29996 17892
rect 30030 17860 30096 17892
rect 30130 17860 30196 17892
rect 30230 17860 30296 17892
rect 29923 17826 29984 17860
rect 30030 17858 30074 17860
rect 30130 17858 30164 17860
rect 30230 17858 30254 17860
rect 30018 17826 30074 17858
rect 30108 17826 30164 17858
rect 30198 17826 30254 17858
rect 30288 17858 30296 17860
rect 30330 17860 30396 17892
rect 30330 17858 30344 17860
rect 30288 17826 30344 17858
rect 30378 17858 30396 17860
rect 30430 17860 30496 17892
rect 30530 17860 30617 17892
rect 30430 17858 30434 17860
rect 30378 17826 30434 17858
rect 30468 17858 30496 17860
rect 30468 17826 30524 17858
rect 30558 17826 30617 17860
rect 29923 17792 30617 17826
rect 29923 17770 29996 17792
rect 30030 17770 30096 17792
rect 30130 17770 30196 17792
rect 30230 17770 30296 17792
rect 29923 17736 29984 17770
rect 30030 17758 30074 17770
rect 30130 17758 30164 17770
rect 30230 17758 30254 17770
rect 30018 17736 30074 17758
rect 30108 17736 30164 17758
rect 30198 17736 30254 17758
rect 30288 17758 30296 17770
rect 30330 17770 30396 17792
rect 30330 17758 30344 17770
rect 30288 17736 30344 17758
rect 30378 17758 30396 17770
rect 30430 17770 30496 17792
rect 30530 17770 30617 17792
rect 30430 17758 30434 17770
rect 30378 17736 30434 17758
rect 30468 17758 30496 17770
rect 30468 17736 30524 17758
rect 30558 17736 30617 17770
rect 29923 17692 30617 17736
rect 29923 17680 29996 17692
rect 30030 17680 30096 17692
rect 30130 17680 30196 17692
rect 30230 17680 30296 17692
rect 29923 17646 29984 17680
rect 30030 17658 30074 17680
rect 30130 17658 30164 17680
rect 30230 17658 30254 17680
rect 30018 17646 30074 17658
rect 30108 17646 30164 17658
rect 30198 17646 30254 17658
rect 30288 17658 30296 17680
rect 30330 17680 30396 17692
rect 30330 17658 30344 17680
rect 30288 17646 30344 17658
rect 30378 17658 30396 17680
rect 30430 17680 30496 17692
rect 30530 17680 30617 17692
rect 30430 17658 30434 17680
rect 30378 17646 30434 17658
rect 30468 17658 30496 17680
rect 30468 17646 30524 17658
rect 30558 17646 30617 17680
rect 29923 17585 30617 17646
rect 30679 18228 30751 18284
rect 30679 18194 30698 18228
rect 30732 18194 30751 18228
rect 30679 18138 30751 18194
rect 30679 18104 30698 18138
rect 30732 18104 30751 18138
rect 30679 18048 30751 18104
rect 30679 18014 30698 18048
rect 30732 18014 30751 18048
rect 30679 17958 30751 18014
rect 30679 17924 30698 17958
rect 30732 17924 30751 17958
rect 30679 17868 30751 17924
rect 30679 17834 30698 17868
rect 30732 17834 30751 17868
rect 30679 17778 30751 17834
rect 30679 17744 30698 17778
rect 30732 17744 30751 17778
rect 30679 17688 30751 17744
rect 30679 17654 30698 17688
rect 30732 17654 30751 17688
rect 30679 17598 30751 17654
rect 29789 17523 29861 17583
rect 30679 17564 30698 17598
rect 30732 17564 30751 17598
rect 30679 17523 30751 17564
rect 29789 17504 30751 17523
rect 29789 17470 29886 17504
rect 29920 17470 29976 17504
rect 30010 17470 30066 17504
rect 30100 17470 30156 17504
rect 30190 17470 30246 17504
rect 30280 17470 30336 17504
rect 30370 17470 30426 17504
rect 30460 17470 30516 17504
rect 30550 17470 30606 17504
rect 30640 17470 30751 17504
rect 29789 17451 30751 17470
rect 30815 18394 30847 18428
rect 30881 18394 31000 18428
rect 31034 18394 31065 18428
rect 32155 18428 32405 18477
rect 30815 18338 31065 18394
rect 30815 18304 30847 18338
rect 30881 18304 31000 18338
rect 31034 18304 31065 18338
rect 30815 18248 31065 18304
rect 30815 18214 30847 18248
rect 30881 18214 31000 18248
rect 31034 18214 31065 18248
rect 30815 18158 31065 18214
rect 30815 18124 30847 18158
rect 30881 18124 31000 18158
rect 31034 18124 31065 18158
rect 30815 18068 31065 18124
rect 30815 18034 30847 18068
rect 30881 18034 31000 18068
rect 31034 18034 31065 18068
rect 30815 17978 31065 18034
rect 30815 17944 30847 17978
rect 30881 17944 31000 17978
rect 31034 17944 31065 17978
rect 30815 17888 31065 17944
rect 30815 17854 30847 17888
rect 30881 17854 31000 17888
rect 31034 17854 31065 17888
rect 30815 17798 31065 17854
rect 30815 17764 30847 17798
rect 30881 17764 31000 17798
rect 31034 17764 31065 17798
rect 30815 17708 31065 17764
rect 30815 17674 30847 17708
rect 30881 17674 31000 17708
rect 31034 17674 31065 17708
rect 30815 17618 31065 17674
rect 30815 17584 30847 17618
rect 30881 17584 31000 17618
rect 31034 17584 31065 17618
rect 30815 17528 31065 17584
rect 30815 17494 30847 17528
rect 30881 17494 31000 17528
rect 31034 17494 31065 17528
rect 29475 17404 29507 17438
rect 29541 17404 29660 17438
rect 29694 17404 29725 17438
rect 29475 17387 29725 17404
rect 30815 17438 31065 17494
rect 31129 18396 32091 18413
rect 31129 18362 31150 18396
rect 31184 18362 31240 18396
rect 31274 18394 31330 18396
rect 31364 18394 31420 18396
rect 31454 18394 31510 18396
rect 31544 18394 31600 18396
rect 31634 18394 31690 18396
rect 31724 18394 31780 18396
rect 31814 18394 31870 18396
rect 31904 18394 31960 18396
rect 31994 18394 32050 18396
rect 31294 18362 31330 18394
rect 31384 18362 31420 18394
rect 31474 18362 31510 18394
rect 31564 18362 31600 18394
rect 31654 18362 31690 18394
rect 31744 18362 31780 18394
rect 31834 18362 31870 18394
rect 31924 18362 31960 18394
rect 32014 18362 32050 18394
rect 32084 18362 32091 18396
rect 31129 18360 31260 18362
rect 31294 18360 31350 18362
rect 31384 18360 31440 18362
rect 31474 18360 31530 18362
rect 31564 18360 31620 18362
rect 31654 18360 31710 18362
rect 31744 18360 31800 18362
rect 31834 18360 31890 18362
rect 31924 18360 31980 18362
rect 32014 18360 32091 18362
rect 31129 18341 32091 18360
rect 31129 18337 31201 18341
rect 31129 18303 31148 18337
rect 31182 18303 31201 18337
rect 31129 18247 31201 18303
rect 32019 18318 32091 18341
rect 32019 18284 32038 18318
rect 32072 18284 32091 18318
rect 31129 18213 31148 18247
rect 31182 18213 31201 18247
rect 31129 18157 31201 18213
rect 31129 18123 31148 18157
rect 31182 18123 31201 18157
rect 31129 18067 31201 18123
rect 31129 18033 31148 18067
rect 31182 18033 31201 18067
rect 31129 17977 31201 18033
rect 31129 17943 31148 17977
rect 31182 17943 31201 17977
rect 31129 17887 31201 17943
rect 31129 17853 31148 17887
rect 31182 17853 31201 17887
rect 31129 17797 31201 17853
rect 31129 17763 31148 17797
rect 31182 17763 31201 17797
rect 31129 17707 31201 17763
rect 31129 17673 31148 17707
rect 31182 17673 31201 17707
rect 31129 17617 31201 17673
rect 31129 17583 31148 17617
rect 31182 17583 31201 17617
rect 31263 18220 31957 18279
rect 31263 18186 31324 18220
rect 31358 18192 31414 18220
rect 31448 18192 31504 18220
rect 31538 18192 31594 18220
rect 31370 18186 31414 18192
rect 31470 18186 31504 18192
rect 31570 18186 31594 18192
rect 31628 18192 31684 18220
rect 31628 18186 31636 18192
rect 31263 18158 31336 18186
rect 31370 18158 31436 18186
rect 31470 18158 31536 18186
rect 31570 18158 31636 18186
rect 31670 18186 31684 18192
rect 31718 18192 31774 18220
rect 31718 18186 31736 18192
rect 31670 18158 31736 18186
rect 31770 18186 31774 18192
rect 31808 18192 31864 18220
rect 31808 18186 31836 18192
rect 31898 18186 31957 18220
rect 31770 18158 31836 18186
rect 31870 18158 31957 18186
rect 31263 18130 31957 18158
rect 31263 18096 31324 18130
rect 31358 18096 31414 18130
rect 31448 18096 31504 18130
rect 31538 18096 31594 18130
rect 31628 18096 31684 18130
rect 31718 18096 31774 18130
rect 31808 18096 31864 18130
rect 31898 18096 31957 18130
rect 31263 18092 31957 18096
rect 31263 18058 31336 18092
rect 31370 18058 31436 18092
rect 31470 18058 31536 18092
rect 31570 18058 31636 18092
rect 31670 18058 31736 18092
rect 31770 18058 31836 18092
rect 31870 18058 31957 18092
rect 31263 18040 31957 18058
rect 31263 18006 31324 18040
rect 31358 18006 31414 18040
rect 31448 18006 31504 18040
rect 31538 18006 31594 18040
rect 31628 18006 31684 18040
rect 31718 18006 31774 18040
rect 31808 18006 31864 18040
rect 31898 18006 31957 18040
rect 31263 17992 31957 18006
rect 31263 17958 31336 17992
rect 31370 17958 31436 17992
rect 31470 17958 31536 17992
rect 31570 17958 31636 17992
rect 31670 17958 31736 17992
rect 31770 17958 31836 17992
rect 31870 17958 31957 17992
rect 31263 17950 31957 17958
rect 31263 17916 31324 17950
rect 31358 17916 31414 17950
rect 31448 17916 31504 17950
rect 31538 17916 31594 17950
rect 31628 17916 31684 17950
rect 31718 17916 31774 17950
rect 31808 17916 31864 17950
rect 31898 17916 31957 17950
rect 31263 17892 31957 17916
rect 31263 17860 31336 17892
rect 31370 17860 31436 17892
rect 31470 17860 31536 17892
rect 31570 17860 31636 17892
rect 31263 17826 31324 17860
rect 31370 17858 31414 17860
rect 31470 17858 31504 17860
rect 31570 17858 31594 17860
rect 31358 17826 31414 17858
rect 31448 17826 31504 17858
rect 31538 17826 31594 17858
rect 31628 17858 31636 17860
rect 31670 17860 31736 17892
rect 31670 17858 31684 17860
rect 31628 17826 31684 17858
rect 31718 17858 31736 17860
rect 31770 17860 31836 17892
rect 31870 17860 31957 17892
rect 31770 17858 31774 17860
rect 31718 17826 31774 17858
rect 31808 17858 31836 17860
rect 31808 17826 31864 17858
rect 31898 17826 31957 17860
rect 31263 17792 31957 17826
rect 31263 17770 31336 17792
rect 31370 17770 31436 17792
rect 31470 17770 31536 17792
rect 31570 17770 31636 17792
rect 31263 17736 31324 17770
rect 31370 17758 31414 17770
rect 31470 17758 31504 17770
rect 31570 17758 31594 17770
rect 31358 17736 31414 17758
rect 31448 17736 31504 17758
rect 31538 17736 31594 17758
rect 31628 17758 31636 17770
rect 31670 17770 31736 17792
rect 31670 17758 31684 17770
rect 31628 17736 31684 17758
rect 31718 17758 31736 17770
rect 31770 17770 31836 17792
rect 31870 17770 31957 17792
rect 31770 17758 31774 17770
rect 31718 17736 31774 17758
rect 31808 17758 31836 17770
rect 31808 17736 31864 17758
rect 31898 17736 31957 17770
rect 31263 17692 31957 17736
rect 31263 17680 31336 17692
rect 31370 17680 31436 17692
rect 31470 17680 31536 17692
rect 31570 17680 31636 17692
rect 31263 17646 31324 17680
rect 31370 17658 31414 17680
rect 31470 17658 31504 17680
rect 31570 17658 31594 17680
rect 31358 17646 31414 17658
rect 31448 17646 31504 17658
rect 31538 17646 31594 17658
rect 31628 17658 31636 17680
rect 31670 17680 31736 17692
rect 31670 17658 31684 17680
rect 31628 17646 31684 17658
rect 31718 17658 31736 17680
rect 31770 17680 31836 17692
rect 31870 17680 31957 17692
rect 31770 17658 31774 17680
rect 31718 17646 31774 17658
rect 31808 17658 31836 17680
rect 31808 17646 31864 17658
rect 31898 17646 31957 17680
rect 31263 17585 31957 17646
rect 32019 18228 32091 18284
rect 32019 18194 32038 18228
rect 32072 18194 32091 18228
rect 32019 18138 32091 18194
rect 32019 18104 32038 18138
rect 32072 18104 32091 18138
rect 32019 18048 32091 18104
rect 32019 18014 32038 18048
rect 32072 18014 32091 18048
rect 32019 17958 32091 18014
rect 32019 17924 32038 17958
rect 32072 17924 32091 17958
rect 32019 17868 32091 17924
rect 32019 17834 32038 17868
rect 32072 17834 32091 17868
rect 32019 17778 32091 17834
rect 32019 17744 32038 17778
rect 32072 17744 32091 17778
rect 32019 17688 32091 17744
rect 32019 17654 32038 17688
rect 32072 17654 32091 17688
rect 32019 17598 32091 17654
rect 31129 17523 31201 17583
rect 32019 17564 32038 17598
rect 32072 17564 32091 17598
rect 32019 17523 32091 17564
rect 31129 17504 32091 17523
rect 31129 17470 31226 17504
rect 31260 17470 31316 17504
rect 31350 17470 31406 17504
rect 31440 17470 31496 17504
rect 31530 17470 31586 17504
rect 31620 17470 31676 17504
rect 31710 17470 31766 17504
rect 31800 17470 31856 17504
rect 31890 17470 31946 17504
rect 31980 17470 32091 17504
rect 31129 17451 32091 17470
rect 32155 18394 32187 18428
rect 32221 18394 32340 18428
rect 32374 18394 32405 18428
rect 33495 18428 33745 18477
rect 32155 18338 32405 18394
rect 32155 18304 32187 18338
rect 32221 18304 32340 18338
rect 32374 18304 32405 18338
rect 32155 18248 32405 18304
rect 32155 18214 32187 18248
rect 32221 18214 32340 18248
rect 32374 18214 32405 18248
rect 32155 18158 32405 18214
rect 32155 18124 32187 18158
rect 32221 18124 32340 18158
rect 32374 18124 32405 18158
rect 32155 18068 32405 18124
rect 32155 18034 32187 18068
rect 32221 18034 32340 18068
rect 32374 18034 32405 18068
rect 32155 17978 32405 18034
rect 32155 17944 32187 17978
rect 32221 17944 32340 17978
rect 32374 17944 32405 17978
rect 32155 17888 32405 17944
rect 32155 17854 32187 17888
rect 32221 17854 32340 17888
rect 32374 17854 32405 17888
rect 32155 17798 32405 17854
rect 32155 17764 32187 17798
rect 32221 17764 32340 17798
rect 32374 17764 32405 17798
rect 32155 17708 32405 17764
rect 32155 17674 32187 17708
rect 32221 17674 32340 17708
rect 32374 17674 32405 17708
rect 32155 17618 32405 17674
rect 32155 17584 32187 17618
rect 32221 17584 32340 17618
rect 32374 17584 32405 17618
rect 32155 17528 32405 17584
rect 32155 17494 32187 17528
rect 32221 17494 32340 17528
rect 32374 17494 32405 17528
rect 30815 17404 30847 17438
rect 30881 17404 31000 17438
rect 31034 17404 31065 17438
rect 30815 17387 31065 17404
rect 32155 17438 32405 17494
rect 32469 18396 33431 18413
rect 32469 18362 32490 18396
rect 32524 18362 32580 18396
rect 32614 18394 32670 18396
rect 32704 18394 32760 18396
rect 32794 18394 32850 18396
rect 32884 18394 32940 18396
rect 32974 18394 33030 18396
rect 33064 18394 33120 18396
rect 33154 18394 33210 18396
rect 33244 18394 33300 18396
rect 33334 18394 33390 18396
rect 32634 18362 32670 18394
rect 32724 18362 32760 18394
rect 32814 18362 32850 18394
rect 32904 18362 32940 18394
rect 32994 18362 33030 18394
rect 33084 18362 33120 18394
rect 33174 18362 33210 18394
rect 33264 18362 33300 18394
rect 33354 18362 33390 18394
rect 33424 18362 33431 18396
rect 32469 18360 32600 18362
rect 32634 18360 32690 18362
rect 32724 18360 32780 18362
rect 32814 18360 32870 18362
rect 32904 18360 32960 18362
rect 32994 18360 33050 18362
rect 33084 18360 33140 18362
rect 33174 18360 33230 18362
rect 33264 18360 33320 18362
rect 33354 18360 33431 18362
rect 32469 18341 33431 18360
rect 32469 18337 32541 18341
rect 32469 18303 32488 18337
rect 32522 18303 32541 18337
rect 32469 18247 32541 18303
rect 33359 18318 33431 18341
rect 33359 18284 33378 18318
rect 33412 18284 33431 18318
rect 32469 18213 32488 18247
rect 32522 18213 32541 18247
rect 32469 18157 32541 18213
rect 32469 18123 32488 18157
rect 32522 18123 32541 18157
rect 32469 18067 32541 18123
rect 32469 18033 32488 18067
rect 32522 18033 32541 18067
rect 32469 17977 32541 18033
rect 32469 17943 32488 17977
rect 32522 17943 32541 17977
rect 32469 17887 32541 17943
rect 32469 17853 32488 17887
rect 32522 17853 32541 17887
rect 32469 17797 32541 17853
rect 32469 17763 32488 17797
rect 32522 17763 32541 17797
rect 32469 17707 32541 17763
rect 32469 17673 32488 17707
rect 32522 17673 32541 17707
rect 32469 17617 32541 17673
rect 32469 17583 32488 17617
rect 32522 17583 32541 17617
rect 32603 18220 33297 18279
rect 32603 18186 32664 18220
rect 32698 18192 32754 18220
rect 32788 18192 32844 18220
rect 32878 18192 32934 18220
rect 32710 18186 32754 18192
rect 32810 18186 32844 18192
rect 32910 18186 32934 18192
rect 32968 18192 33024 18220
rect 32968 18186 32976 18192
rect 32603 18158 32676 18186
rect 32710 18158 32776 18186
rect 32810 18158 32876 18186
rect 32910 18158 32976 18186
rect 33010 18186 33024 18192
rect 33058 18192 33114 18220
rect 33058 18186 33076 18192
rect 33010 18158 33076 18186
rect 33110 18186 33114 18192
rect 33148 18192 33204 18220
rect 33148 18186 33176 18192
rect 33238 18186 33297 18220
rect 33110 18158 33176 18186
rect 33210 18158 33297 18186
rect 32603 18130 33297 18158
rect 32603 18096 32664 18130
rect 32698 18096 32754 18130
rect 32788 18096 32844 18130
rect 32878 18096 32934 18130
rect 32968 18096 33024 18130
rect 33058 18096 33114 18130
rect 33148 18096 33204 18130
rect 33238 18096 33297 18130
rect 32603 18092 33297 18096
rect 32603 18058 32676 18092
rect 32710 18058 32776 18092
rect 32810 18058 32876 18092
rect 32910 18058 32976 18092
rect 33010 18058 33076 18092
rect 33110 18058 33176 18092
rect 33210 18058 33297 18092
rect 32603 18040 33297 18058
rect 32603 18006 32664 18040
rect 32698 18006 32754 18040
rect 32788 18006 32844 18040
rect 32878 18006 32934 18040
rect 32968 18006 33024 18040
rect 33058 18006 33114 18040
rect 33148 18006 33204 18040
rect 33238 18006 33297 18040
rect 32603 17992 33297 18006
rect 32603 17958 32676 17992
rect 32710 17958 32776 17992
rect 32810 17958 32876 17992
rect 32910 17958 32976 17992
rect 33010 17958 33076 17992
rect 33110 17958 33176 17992
rect 33210 17958 33297 17992
rect 32603 17950 33297 17958
rect 32603 17916 32664 17950
rect 32698 17916 32754 17950
rect 32788 17916 32844 17950
rect 32878 17916 32934 17950
rect 32968 17916 33024 17950
rect 33058 17916 33114 17950
rect 33148 17916 33204 17950
rect 33238 17916 33297 17950
rect 32603 17892 33297 17916
rect 32603 17860 32676 17892
rect 32710 17860 32776 17892
rect 32810 17860 32876 17892
rect 32910 17860 32976 17892
rect 32603 17826 32664 17860
rect 32710 17858 32754 17860
rect 32810 17858 32844 17860
rect 32910 17858 32934 17860
rect 32698 17826 32754 17858
rect 32788 17826 32844 17858
rect 32878 17826 32934 17858
rect 32968 17858 32976 17860
rect 33010 17860 33076 17892
rect 33010 17858 33024 17860
rect 32968 17826 33024 17858
rect 33058 17858 33076 17860
rect 33110 17860 33176 17892
rect 33210 17860 33297 17892
rect 33110 17858 33114 17860
rect 33058 17826 33114 17858
rect 33148 17858 33176 17860
rect 33148 17826 33204 17858
rect 33238 17826 33297 17860
rect 32603 17792 33297 17826
rect 32603 17770 32676 17792
rect 32710 17770 32776 17792
rect 32810 17770 32876 17792
rect 32910 17770 32976 17792
rect 32603 17736 32664 17770
rect 32710 17758 32754 17770
rect 32810 17758 32844 17770
rect 32910 17758 32934 17770
rect 32698 17736 32754 17758
rect 32788 17736 32844 17758
rect 32878 17736 32934 17758
rect 32968 17758 32976 17770
rect 33010 17770 33076 17792
rect 33010 17758 33024 17770
rect 32968 17736 33024 17758
rect 33058 17758 33076 17770
rect 33110 17770 33176 17792
rect 33210 17770 33297 17792
rect 33110 17758 33114 17770
rect 33058 17736 33114 17758
rect 33148 17758 33176 17770
rect 33148 17736 33204 17758
rect 33238 17736 33297 17770
rect 32603 17692 33297 17736
rect 32603 17680 32676 17692
rect 32710 17680 32776 17692
rect 32810 17680 32876 17692
rect 32910 17680 32976 17692
rect 32603 17646 32664 17680
rect 32710 17658 32754 17680
rect 32810 17658 32844 17680
rect 32910 17658 32934 17680
rect 32698 17646 32754 17658
rect 32788 17646 32844 17658
rect 32878 17646 32934 17658
rect 32968 17658 32976 17680
rect 33010 17680 33076 17692
rect 33010 17658 33024 17680
rect 32968 17646 33024 17658
rect 33058 17658 33076 17680
rect 33110 17680 33176 17692
rect 33210 17680 33297 17692
rect 33110 17658 33114 17680
rect 33058 17646 33114 17658
rect 33148 17658 33176 17680
rect 33148 17646 33204 17658
rect 33238 17646 33297 17680
rect 32603 17585 33297 17646
rect 33359 18228 33431 18284
rect 33359 18194 33378 18228
rect 33412 18194 33431 18228
rect 33359 18138 33431 18194
rect 33359 18104 33378 18138
rect 33412 18104 33431 18138
rect 33359 18048 33431 18104
rect 33359 18014 33378 18048
rect 33412 18014 33431 18048
rect 33359 17958 33431 18014
rect 33359 17924 33378 17958
rect 33412 17924 33431 17958
rect 33359 17868 33431 17924
rect 33359 17834 33378 17868
rect 33412 17834 33431 17868
rect 33359 17778 33431 17834
rect 33359 17744 33378 17778
rect 33412 17744 33431 17778
rect 33359 17688 33431 17744
rect 33359 17654 33378 17688
rect 33412 17654 33431 17688
rect 33359 17598 33431 17654
rect 32469 17523 32541 17583
rect 33359 17564 33378 17598
rect 33412 17564 33431 17598
rect 33359 17523 33431 17564
rect 32469 17504 33431 17523
rect 32469 17470 32566 17504
rect 32600 17470 32656 17504
rect 32690 17470 32746 17504
rect 32780 17470 32836 17504
rect 32870 17470 32926 17504
rect 32960 17470 33016 17504
rect 33050 17470 33106 17504
rect 33140 17470 33196 17504
rect 33230 17470 33286 17504
rect 33320 17470 33431 17504
rect 32469 17451 33431 17470
rect 33495 18394 33527 18428
rect 33561 18394 33680 18428
rect 33714 18394 33745 18428
rect 34835 18428 35085 18477
rect 33495 18338 33745 18394
rect 33495 18304 33527 18338
rect 33561 18304 33680 18338
rect 33714 18304 33745 18338
rect 33495 18248 33745 18304
rect 33495 18214 33527 18248
rect 33561 18214 33680 18248
rect 33714 18214 33745 18248
rect 33495 18158 33745 18214
rect 33495 18124 33527 18158
rect 33561 18124 33680 18158
rect 33714 18124 33745 18158
rect 33495 18068 33745 18124
rect 33495 18034 33527 18068
rect 33561 18034 33680 18068
rect 33714 18034 33745 18068
rect 33495 17978 33745 18034
rect 33495 17944 33527 17978
rect 33561 17944 33680 17978
rect 33714 17944 33745 17978
rect 33495 17888 33745 17944
rect 33495 17854 33527 17888
rect 33561 17854 33680 17888
rect 33714 17854 33745 17888
rect 33495 17798 33745 17854
rect 33495 17764 33527 17798
rect 33561 17764 33680 17798
rect 33714 17764 33745 17798
rect 33495 17708 33745 17764
rect 33495 17674 33527 17708
rect 33561 17674 33680 17708
rect 33714 17674 33745 17708
rect 33495 17618 33745 17674
rect 33495 17584 33527 17618
rect 33561 17584 33680 17618
rect 33714 17584 33745 17618
rect 33495 17528 33745 17584
rect 33495 17494 33527 17528
rect 33561 17494 33680 17528
rect 33714 17494 33745 17528
rect 32155 17404 32187 17438
rect 32221 17404 32340 17438
rect 32374 17404 32405 17438
rect 32155 17387 32405 17404
rect 33495 17438 33745 17494
rect 33809 18396 34771 18413
rect 33809 18362 33830 18396
rect 33864 18362 33920 18396
rect 33954 18394 34010 18396
rect 34044 18394 34100 18396
rect 34134 18394 34190 18396
rect 34224 18394 34280 18396
rect 34314 18394 34370 18396
rect 34404 18394 34460 18396
rect 34494 18394 34550 18396
rect 34584 18394 34640 18396
rect 34674 18394 34730 18396
rect 33974 18362 34010 18394
rect 34064 18362 34100 18394
rect 34154 18362 34190 18394
rect 34244 18362 34280 18394
rect 34334 18362 34370 18394
rect 34424 18362 34460 18394
rect 34514 18362 34550 18394
rect 34604 18362 34640 18394
rect 34694 18362 34730 18394
rect 34764 18362 34771 18396
rect 33809 18360 33940 18362
rect 33974 18360 34030 18362
rect 34064 18360 34120 18362
rect 34154 18360 34210 18362
rect 34244 18360 34300 18362
rect 34334 18360 34390 18362
rect 34424 18360 34480 18362
rect 34514 18360 34570 18362
rect 34604 18360 34660 18362
rect 34694 18360 34771 18362
rect 33809 18341 34771 18360
rect 33809 18337 33881 18341
rect 33809 18303 33828 18337
rect 33862 18303 33881 18337
rect 33809 18247 33881 18303
rect 34699 18318 34771 18341
rect 34699 18284 34718 18318
rect 34752 18284 34771 18318
rect 33809 18213 33828 18247
rect 33862 18213 33881 18247
rect 33809 18157 33881 18213
rect 33809 18123 33828 18157
rect 33862 18123 33881 18157
rect 33809 18067 33881 18123
rect 33809 18033 33828 18067
rect 33862 18033 33881 18067
rect 33809 17977 33881 18033
rect 33809 17943 33828 17977
rect 33862 17943 33881 17977
rect 33809 17887 33881 17943
rect 33809 17853 33828 17887
rect 33862 17853 33881 17887
rect 33809 17797 33881 17853
rect 33809 17763 33828 17797
rect 33862 17763 33881 17797
rect 33809 17707 33881 17763
rect 33809 17673 33828 17707
rect 33862 17673 33881 17707
rect 33809 17617 33881 17673
rect 33809 17583 33828 17617
rect 33862 17583 33881 17617
rect 33943 18220 34637 18279
rect 33943 18186 34004 18220
rect 34038 18192 34094 18220
rect 34128 18192 34184 18220
rect 34218 18192 34274 18220
rect 34050 18186 34094 18192
rect 34150 18186 34184 18192
rect 34250 18186 34274 18192
rect 34308 18192 34364 18220
rect 34308 18186 34316 18192
rect 33943 18158 34016 18186
rect 34050 18158 34116 18186
rect 34150 18158 34216 18186
rect 34250 18158 34316 18186
rect 34350 18186 34364 18192
rect 34398 18192 34454 18220
rect 34398 18186 34416 18192
rect 34350 18158 34416 18186
rect 34450 18186 34454 18192
rect 34488 18192 34544 18220
rect 34488 18186 34516 18192
rect 34578 18186 34637 18220
rect 34450 18158 34516 18186
rect 34550 18158 34637 18186
rect 33943 18130 34637 18158
rect 33943 18096 34004 18130
rect 34038 18096 34094 18130
rect 34128 18096 34184 18130
rect 34218 18096 34274 18130
rect 34308 18096 34364 18130
rect 34398 18096 34454 18130
rect 34488 18096 34544 18130
rect 34578 18096 34637 18130
rect 33943 18092 34637 18096
rect 33943 18058 34016 18092
rect 34050 18058 34116 18092
rect 34150 18058 34216 18092
rect 34250 18058 34316 18092
rect 34350 18058 34416 18092
rect 34450 18058 34516 18092
rect 34550 18058 34637 18092
rect 33943 18040 34637 18058
rect 33943 18006 34004 18040
rect 34038 18006 34094 18040
rect 34128 18006 34184 18040
rect 34218 18006 34274 18040
rect 34308 18006 34364 18040
rect 34398 18006 34454 18040
rect 34488 18006 34544 18040
rect 34578 18006 34637 18040
rect 33943 17992 34637 18006
rect 33943 17958 34016 17992
rect 34050 17958 34116 17992
rect 34150 17958 34216 17992
rect 34250 17958 34316 17992
rect 34350 17958 34416 17992
rect 34450 17958 34516 17992
rect 34550 17958 34637 17992
rect 33943 17950 34637 17958
rect 33943 17916 34004 17950
rect 34038 17916 34094 17950
rect 34128 17916 34184 17950
rect 34218 17916 34274 17950
rect 34308 17916 34364 17950
rect 34398 17916 34454 17950
rect 34488 17916 34544 17950
rect 34578 17916 34637 17950
rect 33943 17892 34637 17916
rect 33943 17860 34016 17892
rect 34050 17860 34116 17892
rect 34150 17860 34216 17892
rect 34250 17860 34316 17892
rect 33943 17826 34004 17860
rect 34050 17858 34094 17860
rect 34150 17858 34184 17860
rect 34250 17858 34274 17860
rect 34038 17826 34094 17858
rect 34128 17826 34184 17858
rect 34218 17826 34274 17858
rect 34308 17858 34316 17860
rect 34350 17860 34416 17892
rect 34350 17858 34364 17860
rect 34308 17826 34364 17858
rect 34398 17858 34416 17860
rect 34450 17860 34516 17892
rect 34550 17860 34637 17892
rect 34450 17858 34454 17860
rect 34398 17826 34454 17858
rect 34488 17858 34516 17860
rect 34488 17826 34544 17858
rect 34578 17826 34637 17860
rect 33943 17792 34637 17826
rect 33943 17770 34016 17792
rect 34050 17770 34116 17792
rect 34150 17770 34216 17792
rect 34250 17770 34316 17792
rect 33943 17736 34004 17770
rect 34050 17758 34094 17770
rect 34150 17758 34184 17770
rect 34250 17758 34274 17770
rect 34038 17736 34094 17758
rect 34128 17736 34184 17758
rect 34218 17736 34274 17758
rect 34308 17758 34316 17770
rect 34350 17770 34416 17792
rect 34350 17758 34364 17770
rect 34308 17736 34364 17758
rect 34398 17758 34416 17770
rect 34450 17770 34516 17792
rect 34550 17770 34637 17792
rect 34450 17758 34454 17770
rect 34398 17736 34454 17758
rect 34488 17758 34516 17770
rect 34488 17736 34544 17758
rect 34578 17736 34637 17770
rect 33943 17692 34637 17736
rect 33943 17680 34016 17692
rect 34050 17680 34116 17692
rect 34150 17680 34216 17692
rect 34250 17680 34316 17692
rect 33943 17646 34004 17680
rect 34050 17658 34094 17680
rect 34150 17658 34184 17680
rect 34250 17658 34274 17680
rect 34038 17646 34094 17658
rect 34128 17646 34184 17658
rect 34218 17646 34274 17658
rect 34308 17658 34316 17680
rect 34350 17680 34416 17692
rect 34350 17658 34364 17680
rect 34308 17646 34364 17658
rect 34398 17658 34416 17680
rect 34450 17680 34516 17692
rect 34550 17680 34637 17692
rect 34450 17658 34454 17680
rect 34398 17646 34454 17658
rect 34488 17658 34516 17680
rect 34488 17646 34544 17658
rect 34578 17646 34637 17680
rect 33943 17585 34637 17646
rect 34699 18228 34771 18284
rect 34699 18194 34718 18228
rect 34752 18194 34771 18228
rect 34699 18138 34771 18194
rect 34699 18104 34718 18138
rect 34752 18104 34771 18138
rect 34699 18048 34771 18104
rect 34699 18014 34718 18048
rect 34752 18014 34771 18048
rect 34699 17958 34771 18014
rect 34699 17924 34718 17958
rect 34752 17924 34771 17958
rect 34699 17868 34771 17924
rect 34699 17834 34718 17868
rect 34752 17834 34771 17868
rect 34699 17778 34771 17834
rect 34699 17744 34718 17778
rect 34752 17744 34771 17778
rect 34699 17688 34771 17744
rect 34699 17654 34718 17688
rect 34752 17654 34771 17688
rect 34699 17598 34771 17654
rect 33809 17523 33881 17583
rect 34699 17564 34718 17598
rect 34752 17564 34771 17598
rect 34699 17523 34771 17564
rect 33809 17504 34771 17523
rect 33809 17470 33906 17504
rect 33940 17470 33996 17504
rect 34030 17470 34086 17504
rect 34120 17470 34176 17504
rect 34210 17470 34266 17504
rect 34300 17470 34356 17504
rect 34390 17470 34446 17504
rect 34480 17470 34536 17504
rect 34570 17470 34626 17504
rect 34660 17470 34771 17504
rect 33809 17451 34771 17470
rect 34835 18394 34867 18428
rect 34901 18394 35020 18428
rect 35054 18394 35085 18428
rect 36175 18428 36425 18477
rect 34835 18338 35085 18394
rect 34835 18304 34867 18338
rect 34901 18304 35020 18338
rect 35054 18304 35085 18338
rect 34835 18248 35085 18304
rect 34835 18214 34867 18248
rect 34901 18214 35020 18248
rect 35054 18214 35085 18248
rect 34835 18158 35085 18214
rect 34835 18124 34867 18158
rect 34901 18124 35020 18158
rect 35054 18124 35085 18158
rect 34835 18068 35085 18124
rect 34835 18034 34867 18068
rect 34901 18034 35020 18068
rect 35054 18034 35085 18068
rect 34835 17978 35085 18034
rect 34835 17944 34867 17978
rect 34901 17944 35020 17978
rect 35054 17944 35085 17978
rect 34835 17888 35085 17944
rect 34835 17854 34867 17888
rect 34901 17854 35020 17888
rect 35054 17854 35085 17888
rect 34835 17798 35085 17854
rect 34835 17764 34867 17798
rect 34901 17764 35020 17798
rect 35054 17764 35085 17798
rect 34835 17708 35085 17764
rect 34835 17674 34867 17708
rect 34901 17674 35020 17708
rect 35054 17674 35085 17708
rect 34835 17618 35085 17674
rect 34835 17584 34867 17618
rect 34901 17584 35020 17618
rect 35054 17584 35085 17618
rect 34835 17528 35085 17584
rect 34835 17494 34867 17528
rect 34901 17494 35020 17528
rect 35054 17494 35085 17528
rect 33495 17404 33527 17438
rect 33561 17404 33680 17438
rect 33714 17404 33745 17438
rect 33495 17387 33745 17404
rect 34835 17438 35085 17494
rect 35149 18396 36111 18413
rect 35149 18362 35170 18396
rect 35204 18362 35260 18396
rect 35294 18394 35350 18396
rect 35384 18394 35440 18396
rect 35474 18394 35530 18396
rect 35564 18394 35620 18396
rect 35654 18394 35710 18396
rect 35744 18394 35800 18396
rect 35834 18394 35890 18396
rect 35924 18394 35980 18396
rect 36014 18394 36070 18396
rect 35314 18362 35350 18394
rect 35404 18362 35440 18394
rect 35494 18362 35530 18394
rect 35584 18362 35620 18394
rect 35674 18362 35710 18394
rect 35764 18362 35800 18394
rect 35854 18362 35890 18394
rect 35944 18362 35980 18394
rect 36034 18362 36070 18394
rect 36104 18362 36111 18396
rect 35149 18360 35280 18362
rect 35314 18360 35370 18362
rect 35404 18360 35460 18362
rect 35494 18360 35550 18362
rect 35584 18360 35640 18362
rect 35674 18360 35730 18362
rect 35764 18360 35820 18362
rect 35854 18360 35910 18362
rect 35944 18360 36000 18362
rect 36034 18360 36111 18362
rect 35149 18341 36111 18360
rect 35149 18337 35221 18341
rect 35149 18303 35168 18337
rect 35202 18303 35221 18337
rect 35149 18247 35221 18303
rect 36039 18318 36111 18341
rect 36039 18284 36058 18318
rect 36092 18284 36111 18318
rect 35149 18213 35168 18247
rect 35202 18213 35221 18247
rect 35149 18157 35221 18213
rect 35149 18123 35168 18157
rect 35202 18123 35221 18157
rect 35149 18067 35221 18123
rect 35149 18033 35168 18067
rect 35202 18033 35221 18067
rect 35149 17977 35221 18033
rect 35149 17943 35168 17977
rect 35202 17943 35221 17977
rect 35149 17887 35221 17943
rect 35149 17853 35168 17887
rect 35202 17853 35221 17887
rect 35149 17797 35221 17853
rect 35149 17763 35168 17797
rect 35202 17763 35221 17797
rect 35149 17707 35221 17763
rect 35149 17673 35168 17707
rect 35202 17673 35221 17707
rect 35149 17617 35221 17673
rect 35149 17583 35168 17617
rect 35202 17583 35221 17617
rect 35283 18220 35977 18279
rect 35283 18186 35344 18220
rect 35378 18192 35434 18220
rect 35468 18192 35524 18220
rect 35558 18192 35614 18220
rect 35390 18186 35434 18192
rect 35490 18186 35524 18192
rect 35590 18186 35614 18192
rect 35648 18192 35704 18220
rect 35648 18186 35656 18192
rect 35283 18158 35356 18186
rect 35390 18158 35456 18186
rect 35490 18158 35556 18186
rect 35590 18158 35656 18186
rect 35690 18186 35704 18192
rect 35738 18192 35794 18220
rect 35738 18186 35756 18192
rect 35690 18158 35756 18186
rect 35790 18186 35794 18192
rect 35828 18192 35884 18220
rect 35828 18186 35856 18192
rect 35918 18186 35977 18220
rect 35790 18158 35856 18186
rect 35890 18158 35977 18186
rect 35283 18130 35977 18158
rect 35283 18096 35344 18130
rect 35378 18096 35434 18130
rect 35468 18096 35524 18130
rect 35558 18096 35614 18130
rect 35648 18096 35704 18130
rect 35738 18096 35794 18130
rect 35828 18096 35884 18130
rect 35918 18096 35977 18130
rect 35283 18092 35977 18096
rect 35283 18058 35356 18092
rect 35390 18058 35456 18092
rect 35490 18058 35556 18092
rect 35590 18058 35656 18092
rect 35690 18058 35756 18092
rect 35790 18058 35856 18092
rect 35890 18058 35977 18092
rect 35283 18040 35977 18058
rect 35283 18006 35344 18040
rect 35378 18006 35434 18040
rect 35468 18006 35524 18040
rect 35558 18006 35614 18040
rect 35648 18006 35704 18040
rect 35738 18006 35794 18040
rect 35828 18006 35884 18040
rect 35918 18006 35977 18040
rect 35283 17992 35977 18006
rect 35283 17958 35356 17992
rect 35390 17958 35456 17992
rect 35490 17958 35556 17992
rect 35590 17958 35656 17992
rect 35690 17958 35756 17992
rect 35790 17958 35856 17992
rect 35890 17958 35977 17992
rect 35283 17950 35977 17958
rect 35283 17916 35344 17950
rect 35378 17916 35434 17950
rect 35468 17916 35524 17950
rect 35558 17916 35614 17950
rect 35648 17916 35704 17950
rect 35738 17916 35794 17950
rect 35828 17916 35884 17950
rect 35918 17916 35977 17950
rect 35283 17892 35977 17916
rect 35283 17860 35356 17892
rect 35390 17860 35456 17892
rect 35490 17860 35556 17892
rect 35590 17860 35656 17892
rect 35283 17826 35344 17860
rect 35390 17858 35434 17860
rect 35490 17858 35524 17860
rect 35590 17858 35614 17860
rect 35378 17826 35434 17858
rect 35468 17826 35524 17858
rect 35558 17826 35614 17858
rect 35648 17858 35656 17860
rect 35690 17860 35756 17892
rect 35690 17858 35704 17860
rect 35648 17826 35704 17858
rect 35738 17858 35756 17860
rect 35790 17860 35856 17892
rect 35890 17860 35977 17892
rect 35790 17858 35794 17860
rect 35738 17826 35794 17858
rect 35828 17858 35856 17860
rect 35828 17826 35884 17858
rect 35918 17826 35977 17860
rect 35283 17792 35977 17826
rect 35283 17770 35356 17792
rect 35390 17770 35456 17792
rect 35490 17770 35556 17792
rect 35590 17770 35656 17792
rect 35283 17736 35344 17770
rect 35390 17758 35434 17770
rect 35490 17758 35524 17770
rect 35590 17758 35614 17770
rect 35378 17736 35434 17758
rect 35468 17736 35524 17758
rect 35558 17736 35614 17758
rect 35648 17758 35656 17770
rect 35690 17770 35756 17792
rect 35690 17758 35704 17770
rect 35648 17736 35704 17758
rect 35738 17758 35756 17770
rect 35790 17770 35856 17792
rect 35890 17770 35977 17792
rect 35790 17758 35794 17770
rect 35738 17736 35794 17758
rect 35828 17758 35856 17770
rect 35828 17736 35884 17758
rect 35918 17736 35977 17770
rect 35283 17692 35977 17736
rect 35283 17680 35356 17692
rect 35390 17680 35456 17692
rect 35490 17680 35556 17692
rect 35590 17680 35656 17692
rect 35283 17646 35344 17680
rect 35390 17658 35434 17680
rect 35490 17658 35524 17680
rect 35590 17658 35614 17680
rect 35378 17646 35434 17658
rect 35468 17646 35524 17658
rect 35558 17646 35614 17658
rect 35648 17658 35656 17680
rect 35690 17680 35756 17692
rect 35690 17658 35704 17680
rect 35648 17646 35704 17658
rect 35738 17658 35756 17680
rect 35790 17680 35856 17692
rect 35890 17680 35977 17692
rect 35790 17658 35794 17680
rect 35738 17646 35794 17658
rect 35828 17658 35856 17680
rect 35828 17646 35884 17658
rect 35918 17646 35977 17680
rect 35283 17585 35977 17646
rect 36039 18228 36111 18284
rect 36039 18194 36058 18228
rect 36092 18194 36111 18228
rect 36039 18138 36111 18194
rect 36039 18104 36058 18138
rect 36092 18104 36111 18138
rect 36039 18048 36111 18104
rect 36039 18014 36058 18048
rect 36092 18014 36111 18048
rect 36039 17958 36111 18014
rect 36039 17924 36058 17958
rect 36092 17924 36111 17958
rect 36039 17868 36111 17924
rect 36039 17834 36058 17868
rect 36092 17834 36111 17868
rect 36039 17778 36111 17834
rect 36039 17744 36058 17778
rect 36092 17744 36111 17778
rect 36039 17688 36111 17744
rect 36039 17654 36058 17688
rect 36092 17654 36111 17688
rect 36039 17598 36111 17654
rect 35149 17523 35221 17583
rect 36039 17564 36058 17598
rect 36092 17564 36111 17598
rect 36039 17523 36111 17564
rect 35149 17504 36111 17523
rect 35149 17470 35246 17504
rect 35280 17470 35336 17504
rect 35370 17470 35426 17504
rect 35460 17470 35516 17504
rect 35550 17470 35606 17504
rect 35640 17470 35696 17504
rect 35730 17470 35786 17504
rect 35820 17470 35876 17504
rect 35910 17470 35966 17504
rect 36000 17470 36111 17504
rect 35149 17451 36111 17470
rect 36175 18394 36207 18428
rect 36241 18394 36360 18428
rect 36394 18394 36425 18428
rect 37515 18428 37765 18477
rect 36175 18338 36425 18394
rect 36175 18304 36207 18338
rect 36241 18304 36360 18338
rect 36394 18304 36425 18338
rect 36175 18248 36425 18304
rect 36175 18214 36207 18248
rect 36241 18214 36360 18248
rect 36394 18214 36425 18248
rect 36175 18158 36425 18214
rect 36175 18124 36207 18158
rect 36241 18124 36360 18158
rect 36394 18124 36425 18158
rect 36175 18068 36425 18124
rect 36175 18034 36207 18068
rect 36241 18034 36360 18068
rect 36394 18034 36425 18068
rect 36175 17978 36425 18034
rect 36175 17944 36207 17978
rect 36241 17944 36360 17978
rect 36394 17944 36425 17978
rect 36175 17888 36425 17944
rect 36175 17854 36207 17888
rect 36241 17854 36360 17888
rect 36394 17854 36425 17888
rect 36175 17798 36425 17854
rect 36175 17764 36207 17798
rect 36241 17764 36360 17798
rect 36394 17764 36425 17798
rect 36175 17708 36425 17764
rect 36175 17674 36207 17708
rect 36241 17674 36360 17708
rect 36394 17674 36425 17708
rect 36175 17618 36425 17674
rect 36175 17584 36207 17618
rect 36241 17584 36360 17618
rect 36394 17584 36425 17618
rect 36175 17528 36425 17584
rect 36175 17494 36207 17528
rect 36241 17494 36360 17528
rect 36394 17494 36425 17528
rect 34835 17404 34867 17438
rect 34901 17404 35020 17438
rect 35054 17404 35085 17438
rect 34835 17387 35085 17404
rect 36175 17438 36425 17494
rect 36489 18396 37451 18413
rect 36489 18362 36510 18396
rect 36544 18362 36600 18396
rect 36634 18394 36690 18396
rect 36724 18394 36780 18396
rect 36814 18394 36870 18396
rect 36904 18394 36960 18396
rect 36994 18394 37050 18396
rect 37084 18394 37140 18396
rect 37174 18394 37230 18396
rect 37264 18394 37320 18396
rect 37354 18394 37410 18396
rect 36654 18362 36690 18394
rect 36744 18362 36780 18394
rect 36834 18362 36870 18394
rect 36924 18362 36960 18394
rect 37014 18362 37050 18394
rect 37104 18362 37140 18394
rect 37194 18362 37230 18394
rect 37284 18362 37320 18394
rect 37374 18362 37410 18394
rect 37444 18362 37451 18396
rect 36489 18360 36620 18362
rect 36654 18360 36710 18362
rect 36744 18360 36800 18362
rect 36834 18360 36890 18362
rect 36924 18360 36980 18362
rect 37014 18360 37070 18362
rect 37104 18360 37160 18362
rect 37194 18360 37250 18362
rect 37284 18360 37340 18362
rect 37374 18360 37451 18362
rect 36489 18341 37451 18360
rect 36489 18337 36561 18341
rect 36489 18303 36508 18337
rect 36542 18303 36561 18337
rect 36489 18247 36561 18303
rect 37379 18318 37451 18341
rect 37379 18284 37398 18318
rect 37432 18284 37451 18318
rect 36489 18213 36508 18247
rect 36542 18213 36561 18247
rect 36489 18157 36561 18213
rect 36489 18123 36508 18157
rect 36542 18123 36561 18157
rect 36489 18067 36561 18123
rect 36489 18033 36508 18067
rect 36542 18033 36561 18067
rect 36489 17977 36561 18033
rect 36489 17943 36508 17977
rect 36542 17943 36561 17977
rect 36489 17887 36561 17943
rect 36489 17853 36508 17887
rect 36542 17853 36561 17887
rect 36489 17797 36561 17853
rect 36489 17763 36508 17797
rect 36542 17763 36561 17797
rect 36489 17707 36561 17763
rect 36489 17673 36508 17707
rect 36542 17673 36561 17707
rect 36489 17617 36561 17673
rect 36489 17583 36508 17617
rect 36542 17583 36561 17617
rect 36623 18220 37317 18279
rect 36623 18186 36684 18220
rect 36718 18192 36774 18220
rect 36808 18192 36864 18220
rect 36898 18192 36954 18220
rect 36730 18186 36774 18192
rect 36830 18186 36864 18192
rect 36930 18186 36954 18192
rect 36988 18192 37044 18220
rect 36988 18186 36996 18192
rect 36623 18158 36696 18186
rect 36730 18158 36796 18186
rect 36830 18158 36896 18186
rect 36930 18158 36996 18186
rect 37030 18186 37044 18192
rect 37078 18192 37134 18220
rect 37078 18186 37096 18192
rect 37030 18158 37096 18186
rect 37130 18186 37134 18192
rect 37168 18192 37224 18220
rect 37168 18186 37196 18192
rect 37258 18186 37317 18220
rect 37130 18158 37196 18186
rect 37230 18158 37317 18186
rect 36623 18130 37317 18158
rect 36623 18096 36684 18130
rect 36718 18096 36774 18130
rect 36808 18096 36864 18130
rect 36898 18096 36954 18130
rect 36988 18096 37044 18130
rect 37078 18096 37134 18130
rect 37168 18096 37224 18130
rect 37258 18096 37317 18130
rect 36623 18092 37317 18096
rect 36623 18058 36696 18092
rect 36730 18058 36796 18092
rect 36830 18058 36896 18092
rect 36930 18058 36996 18092
rect 37030 18058 37096 18092
rect 37130 18058 37196 18092
rect 37230 18058 37317 18092
rect 36623 18040 37317 18058
rect 36623 18006 36684 18040
rect 36718 18006 36774 18040
rect 36808 18006 36864 18040
rect 36898 18006 36954 18040
rect 36988 18006 37044 18040
rect 37078 18006 37134 18040
rect 37168 18006 37224 18040
rect 37258 18006 37317 18040
rect 36623 17992 37317 18006
rect 36623 17958 36696 17992
rect 36730 17958 36796 17992
rect 36830 17958 36896 17992
rect 36930 17958 36996 17992
rect 37030 17958 37096 17992
rect 37130 17958 37196 17992
rect 37230 17958 37317 17992
rect 36623 17950 37317 17958
rect 36623 17916 36684 17950
rect 36718 17916 36774 17950
rect 36808 17916 36864 17950
rect 36898 17916 36954 17950
rect 36988 17916 37044 17950
rect 37078 17916 37134 17950
rect 37168 17916 37224 17950
rect 37258 17916 37317 17950
rect 36623 17892 37317 17916
rect 36623 17860 36696 17892
rect 36730 17860 36796 17892
rect 36830 17860 36896 17892
rect 36930 17860 36996 17892
rect 36623 17826 36684 17860
rect 36730 17858 36774 17860
rect 36830 17858 36864 17860
rect 36930 17858 36954 17860
rect 36718 17826 36774 17858
rect 36808 17826 36864 17858
rect 36898 17826 36954 17858
rect 36988 17858 36996 17860
rect 37030 17860 37096 17892
rect 37030 17858 37044 17860
rect 36988 17826 37044 17858
rect 37078 17858 37096 17860
rect 37130 17860 37196 17892
rect 37230 17860 37317 17892
rect 37130 17858 37134 17860
rect 37078 17826 37134 17858
rect 37168 17858 37196 17860
rect 37168 17826 37224 17858
rect 37258 17826 37317 17860
rect 36623 17792 37317 17826
rect 36623 17770 36696 17792
rect 36730 17770 36796 17792
rect 36830 17770 36896 17792
rect 36930 17770 36996 17792
rect 36623 17736 36684 17770
rect 36730 17758 36774 17770
rect 36830 17758 36864 17770
rect 36930 17758 36954 17770
rect 36718 17736 36774 17758
rect 36808 17736 36864 17758
rect 36898 17736 36954 17758
rect 36988 17758 36996 17770
rect 37030 17770 37096 17792
rect 37030 17758 37044 17770
rect 36988 17736 37044 17758
rect 37078 17758 37096 17770
rect 37130 17770 37196 17792
rect 37230 17770 37317 17792
rect 37130 17758 37134 17770
rect 37078 17736 37134 17758
rect 37168 17758 37196 17770
rect 37168 17736 37224 17758
rect 37258 17736 37317 17770
rect 36623 17692 37317 17736
rect 36623 17680 36696 17692
rect 36730 17680 36796 17692
rect 36830 17680 36896 17692
rect 36930 17680 36996 17692
rect 36623 17646 36684 17680
rect 36730 17658 36774 17680
rect 36830 17658 36864 17680
rect 36930 17658 36954 17680
rect 36718 17646 36774 17658
rect 36808 17646 36864 17658
rect 36898 17646 36954 17658
rect 36988 17658 36996 17680
rect 37030 17680 37096 17692
rect 37030 17658 37044 17680
rect 36988 17646 37044 17658
rect 37078 17658 37096 17680
rect 37130 17680 37196 17692
rect 37230 17680 37317 17692
rect 37130 17658 37134 17680
rect 37078 17646 37134 17658
rect 37168 17658 37196 17680
rect 37168 17646 37224 17658
rect 37258 17646 37317 17680
rect 36623 17585 37317 17646
rect 37379 18228 37451 18284
rect 37379 18194 37398 18228
rect 37432 18194 37451 18228
rect 37379 18138 37451 18194
rect 37379 18104 37398 18138
rect 37432 18104 37451 18138
rect 37379 18048 37451 18104
rect 37379 18014 37398 18048
rect 37432 18014 37451 18048
rect 37379 17958 37451 18014
rect 37379 17924 37398 17958
rect 37432 17924 37451 17958
rect 37379 17868 37451 17924
rect 37379 17834 37398 17868
rect 37432 17834 37451 17868
rect 37379 17778 37451 17834
rect 37379 17744 37398 17778
rect 37432 17744 37451 17778
rect 37379 17688 37451 17744
rect 37379 17654 37398 17688
rect 37432 17654 37451 17688
rect 37379 17598 37451 17654
rect 36489 17523 36561 17583
rect 37379 17564 37398 17598
rect 37432 17564 37451 17598
rect 37379 17523 37451 17564
rect 36489 17504 37451 17523
rect 36489 17470 36586 17504
rect 36620 17470 36676 17504
rect 36710 17470 36766 17504
rect 36800 17470 36856 17504
rect 36890 17470 36946 17504
rect 36980 17470 37036 17504
rect 37070 17470 37126 17504
rect 37160 17470 37216 17504
rect 37250 17470 37306 17504
rect 37340 17470 37451 17504
rect 36489 17451 37451 17470
rect 37515 18394 37547 18428
rect 37581 18394 37700 18428
rect 37734 18394 37765 18428
rect 38855 18428 38954 18477
rect 37515 18338 37765 18394
rect 37515 18304 37547 18338
rect 37581 18304 37700 18338
rect 37734 18304 37765 18338
rect 37515 18248 37765 18304
rect 37515 18214 37547 18248
rect 37581 18214 37700 18248
rect 37734 18214 37765 18248
rect 37515 18158 37765 18214
rect 37515 18124 37547 18158
rect 37581 18124 37700 18158
rect 37734 18124 37765 18158
rect 37515 18068 37765 18124
rect 37515 18034 37547 18068
rect 37581 18034 37700 18068
rect 37734 18034 37765 18068
rect 37515 17978 37765 18034
rect 37515 17944 37547 17978
rect 37581 17944 37700 17978
rect 37734 17944 37765 17978
rect 37515 17888 37765 17944
rect 37515 17854 37547 17888
rect 37581 17854 37700 17888
rect 37734 17854 37765 17888
rect 37515 17798 37765 17854
rect 37515 17764 37547 17798
rect 37581 17764 37700 17798
rect 37734 17764 37765 17798
rect 37515 17708 37765 17764
rect 37515 17674 37547 17708
rect 37581 17674 37700 17708
rect 37734 17674 37765 17708
rect 37515 17618 37765 17674
rect 37515 17584 37547 17618
rect 37581 17584 37700 17618
rect 37734 17584 37765 17618
rect 37515 17528 37765 17584
rect 37515 17494 37547 17528
rect 37581 17494 37700 17528
rect 37734 17494 37765 17528
rect 36175 17404 36207 17438
rect 36241 17404 36360 17438
rect 36394 17404 36425 17438
rect 36175 17387 36425 17404
rect 37515 17438 37765 17494
rect 37829 18396 38791 18413
rect 37829 18362 37850 18396
rect 37884 18362 37940 18396
rect 37974 18394 38030 18396
rect 38064 18394 38120 18396
rect 38154 18394 38210 18396
rect 38244 18394 38300 18396
rect 38334 18394 38390 18396
rect 38424 18394 38480 18396
rect 38514 18394 38570 18396
rect 38604 18394 38660 18396
rect 38694 18394 38750 18396
rect 37994 18362 38030 18394
rect 38084 18362 38120 18394
rect 38174 18362 38210 18394
rect 38264 18362 38300 18394
rect 38354 18362 38390 18394
rect 38444 18362 38480 18394
rect 38534 18362 38570 18394
rect 38624 18362 38660 18394
rect 38714 18362 38750 18394
rect 38784 18362 38791 18396
rect 37829 18360 37960 18362
rect 37994 18360 38050 18362
rect 38084 18360 38140 18362
rect 38174 18360 38230 18362
rect 38264 18360 38320 18362
rect 38354 18360 38410 18362
rect 38444 18360 38500 18362
rect 38534 18360 38590 18362
rect 38624 18360 38680 18362
rect 38714 18360 38791 18362
rect 37829 18341 38791 18360
rect 37829 18337 37901 18341
rect 37829 18303 37848 18337
rect 37882 18303 37901 18337
rect 37829 18247 37901 18303
rect 38719 18318 38791 18341
rect 38719 18284 38738 18318
rect 38772 18284 38791 18318
rect 37829 18213 37848 18247
rect 37882 18213 37901 18247
rect 37829 18157 37901 18213
rect 37829 18123 37848 18157
rect 37882 18123 37901 18157
rect 37829 18067 37901 18123
rect 37829 18033 37848 18067
rect 37882 18033 37901 18067
rect 37829 17977 37901 18033
rect 37829 17943 37848 17977
rect 37882 17943 37901 17977
rect 37829 17887 37901 17943
rect 37829 17853 37848 17887
rect 37882 17853 37901 17887
rect 37829 17797 37901 17853
rect 37829 17763 37848 17797
rect 37882 17763 37901 17797
rect 37829 17707 37901 17763
rect 37829 17673 37848 17707
rect 37882 17673 37901 17707
rect 37829 17617 37901 17673
rect 37829 17583 37848 17617
rect 37882 17583 37901 17617
rect 37963 18220 38657 18279
rect 37963 18186 38024 18220
rect 38058 18192 38114 18220
rect 38148 18192 38204 18220
rect 38238 18192 38294 18220
rect 38070 18186 38114 18192
rect 38170 18186 38204 18192
rect 38270 18186 38294 18192
rect 38328 18192 38384 18220
rect 38328 18186 38336 18192
rect 37963 18158 38036 18186
rect 38070 18158 38136 18186
rect 38170 18158 38236 18186
rect 38270 18158 38336 18186
rect 38370 18186 38384 18192
rect 38418 18192 38474 18220
rect 38418 18186 38436 18192
rect 38370 18158 38436 18186
rect 38470 18186 38474 18192
rect 38508 18192 38564 18220
rect 38508 18186 38536 18192
rect 38598 18186 38657 18220
rect 38470 18158 38536 18186
rect 38570 18158 38657 18186
rect 37963 18130 38657 18158
rect 37963 18096 38024 18130
rect 38058 18096 38114 18130
rect 38148 18096 38204 18130
rect 38238 18096 38294 18130
rect 38328 18096 38384 18130
rect 38418 18096 38474 18130
rect 38508 18096 38564 18130
rect 38598 18096 38657 18130
rect 37963 18092 38657 18096
rect 37963 18058 38036 18092
rect 38070 18058 38136 18092
rect 38170 18058 38236 18092
rect 38270 18058 38336 18092
rect 38370 18058 38436 18092
rect 38470 18058 38536 18092
rect 38570 18058 38657 18092
rect 37963 18040 38657 18058
rect 37963 18006 38024 18040
rect 38058 18006 38114 18040
rect 38148 18006 38204 18040
rect 38238 18006 38294 18040
rect 38328 18006 38384 18040
rect 38418 18006 38474 18040
rect 38508 18006 38564 18040
rect 38598 18006 38657 18040
rect 37963 17992 38657 18006
rect 37963 17958 38036 17992
rect 38070 17958 38136 17992
rect 38170 17958 38236 17992
rect 38270 17958 38336 17992
rect 38370 17958 38436 17992
rect 38470 17958 38536 17992
rect 38570 17958 38657 17992
rect 37963 17950 38657 17958
rect 37963 17916 38024 17950
rect 38058 17916 38114 17950
rect 38148 17916 38204 17950
rect 38238 17916 38294 17950
rect 38328 17916 38384 17950
rect 38418 17916 38474 17950
rect 38508 17916 38564 17950
rect 38598 17916 38657 17950
rect 37963 17892 38657 17916
rect 37963 17860 38036 17892
rect 38070 17860 38136 17892
rect 38170 17860 38236 17892
rect 38270 17860 38336 17892
rect 37963 17826 38024 17860
rect 38070 17858 38114 17860
rect 38170 17858 38204 17860
rect 38270 17858 38294 17860
rect 38058 17826 38114 17858
rect 38148 17826 38204 17858
rect 38238 17826 38294 17858
rect 38328 17858 38336 17860
rect 38370 17860 38436 17892
rect 38370 17858 38384 17860
rect 38328 17826 38384 17858
rect 38418 17858 38436 17860
rect 38470 17860 38536 17892
rect 38570 17860 38657 17892
rect 38470 17858 38474 17860
rect 38418 17826 38474 17858
rect 38508 17858 38536 17860
rect 38508 17826 38564 17858
rect 38598 17826 38657 17860
rect 37963 17792 38657 17826
rect 37963 17770 38036 17792
rect 38070 17770 38136 17792
rect 38170 17770 38236 17792
rect 38270 17770 38336 17792
rect 37963 17736 38024 17770
rect 38070 17758 38114 17770
rect 38170 17758 38204 17770
rect 38270 17758 38294 17770
rect 38058 17736 38114 17758
rect 38148 17736 38204 17758
rect 38238 17736 38294 17758
rect 38328 17758 38336 17770
rect 38370 17770 38436 17792
rect 38370 17758 38384 17770
rect 38328 17736 38384 17758
rect 38418 17758 38436 17770
rect 38470 17770 38536 17792
rect 38570 17770 38657 17792
rect 38470 17758 38474 17770
rect 38418 17736 38474 17758
rect 38508 17758 38536 17770
rect 38508 17736 38564 17758
rect 38598 17736 38657 17770
rect 37963 17692 38657 17736
rect 37963 17680 38036 17692
rect 38070 17680 38136 17692
rect 38170 17680 38236 17692
rect 38270 17680 38336 17692
rect 37963 17646 38024 17680
rect 38070 17658 38114 17680
rect 38170 17658 38204 17680
rect 38270 17658 38294 17680
rect 38058 17646 38114 17658
rect 38148 17646 38204 17658
rect 38238 17646 38294 17658
rect 38328 17658 38336 17680
rect 38370 17680 38436 17692
rect 38370 17658 38384 17680
rect 38328 17646 38384 17658
rect 38418 17658 38436 17680
rect 38470 17680 38536 17692
rect 38570 17680 38657 17692
rect 38470 17658 38474 17680
rect 38418 17646 38474 17658
rect 38508 17658 38536 17680
rect 38508 17646 38564 17658
rect 38598 17646 38657 17680
rect 37963 17585 38657 17646
rect 38719 18228 38791 18284
rect 38719 18194 38738 18228
rect 38772 18194 38791 18228
rect 38719 18138 38791 18194
rect 38719 18104 38738 18138
rect 38772 18104 38791 18138
rect 38719 18048 38791 18104
rect 38719 18014 38738 18048
rect 38772 18014 38791 18048
rect 38719 17958 38791 18014
rect 38719 17924 38738 17958
rect 38772 17924 38791 17958
rect 38719 17868 38791 17924
rect 38719 17834 38738 17868
rect 38772 17834 38791 17868
rect 38719 17778 38791 17834
rect 38719 17744 38738 17778
rect 38772 17744 38791 17778
rect 38719 17688 38791 17744
rect 38719 17654 38738 17688
rect 38772 17654 38791 17688
rect 38719 17598 38791 17654
rect 37829 17523 37901 17583
rect 38719 17564 38738 17598
rect 38772 17564 38791 17598
rect 38719 17523 38791 17564
rect 37829 17504 38791 17523
rect 37829 17470 37926 17504
rect 37960 17470 38016 17504
rect 38050 17470 38106 17504
rect 38140 17470 38196 17504
rect 38230 17470 38286 17504
rect 38320 17470 38376 17504
rect 38410 17470 38466 17504
rect 38500 17470 38556 17504
rect 38590 17470 38646 17504
rect 38680 17470 38791 17504
rect 37829 17451 38791 17470
rect 38855 18394 38887 18428
rect 38921 18394 38954 18428
rect 38855 18338 38954 18394
rect 38855 18304 38887 18338
rect 38921 18304 38954 18338
rect 38855 18248 38954 18304
rect 38855 18214 38887 18248
rect 38921 18214 38954 18248
rect 38855 18158 38954 18214
rect 38855 18124 38887 18158
rect 38921 18124 38954 18158
rect 38855 18068 38954 18124
rect 38855 18034 38887 18068
rect 38921 18034 38954 18068
rect 38855 17978 38954 18034
rect 38855 17944 38887 17978
rect 38921 17944 38954 17978
rect 38855 17888 38954 17944
rect 38855 17854 38887 17888
rect 38921 17854 38954 17888
rect 38855 17798 38954 17854
rect 38855 17764 38887 17798
rect 38921 17764 38954 17798
rect 38855 17708 38954 17764
rect 38855 17674 38887 17708
rect 38921 17674 38954 17708
rect 40168 17923 40784 17962
rect 40168 17821 40255 17923
rect 40697 17821 40784 17923
rect 38855 17618 38954 17674
rect 38855 17584 38887 17618
rect 38921 17584 38954 17618
rect 38855 17528 38954 17584
rect 38855 17494 38887 17528
rect 38921 17494 38954 17528
rect 37515 17404 37547 17438
rect 37581 17404 37700 17438
rect 37734 17404 37765 17438
rect 37515 17387 37765 17404
rect 38855 17438 38954 17494
rect 38855 17404 38887 17438
rect 38921 17404 38954 17438
rect 38855 17387 38954 17404
rect 28286 17354 38954 17387
rect 28286 17320 28416 17354
rect 28450 17320 28506 17354
rect 28540 17320 28596 17354
rect 28630 17320 28686 17354
rect 28720 17320 28776 17354
rect 28810 17320 28866 17354
rect 28900 17320 28956 17354
rect 28990 17320 29046 17354
rect 29080 17320 29136 17354
rect 29170 17320 29226 17354
rect 29260 17320 29316 17354
rect 29350 17320 29406 17354
rect 29440 17320 29756 17354
rect 29790 17320 29846 17354
rect 29880 17320 29936 17354
rect 29970 17320 30026 17354
rect 30060 17320 30116 17354
rect 30150 17320 30206 17354
rect 30240 17320 30296 17354
rect 30330 17320 30386 17354
rect 30420 17320 30476 17354
rect 30510 17320 30566 17354
rect 30600 17320 30656 17354
rect 30690 17320 30746 17354
rect 30780 17320 31096 17354
rect 31130 17320 31186 17354
rect 31220 17320 31276 17354
rect 31310 17320 31366 17354
rect 31400 17320 31456 17354
rect 31490 17320 31546 17354
rect 31580 17320 31636 17354
rect 31670 17320 31726 17354
rect 31760 17320 31816 17354
rect 31850 17320 31906 17354
rect 31940 17320 31996 17354
rect 32030 17320 32086 17354
rect 32120 17320 32436 17354
rect 32470 17320 32526 17354
rect 32560 17320 32616 17354
rect 32650 17320 32706 17354
rect 32740 17320 32796 17354
rect 32830 17320 32886 17354
rect 32920 17320 32976 17354
rect 33010 17320 33066 17354
rect 33100 17320 33156 17354
rect 33190 17320 33246 17354
rect 33280 17320 33336 17354
rect 33370 17320 33426 17354
rect 33460 17320 33776 17354
rect 33810 17320 33866 17354
rect 33900 17320 33956 17354
rect 33990 17320 34046 17354
rect 34080 17320 34136 17354
rect 34170 17320 34226 17354
rect 34260 17320 34316 17354
rect 34350 17320 34406 17354
rect 34440 17320 34496 17354
rect 34530 17320 34586 17354
rect 34620 17320 34676 17354
rect 34710 17320 34766 17354
rect 34800 17320 35116 17354
rect 35150 17320 35206 17354
rect 35240 17320 35296 17354
rect 35330 17320 35386 17354
rect 35420 17320 35476 17354
rect 35510 17320 35566 17354
rect 35600 17320 35656 17354
rect 35690 17320 35746 17354
rect 35780 17320 35836 17354
rect 35870 17320 35926 17354
rect 35960 17320 36016 17354
rect 36050 17320 36106 17354
rect 36140 17320 36456 17354
rect 36490 17320 36546 17354
rect 36580 17320 36636 17354
rect 36670 17320 36726 17354
rect 36760 17320 36816 17354
rect 36850 17320 36906 17354
rect 36940 17320 36996 17354
rect 37030 17320 37086 17354
rect 37120 17320 37176 17354
rect 37210 17320 37266 17354
rect 37300 17320 37356 17354
rect 37390 17320 37446 17354
rect 37480 17320 37796 17354
rect 37830 17320 37886 17354
rect 37920 17320 37976 17354
rect 38010 17320 38066 17354
rect 38100 17320 38156 17354
rect 38190 17320 38246 17354
rect 38280 17320 38336 17354
rect 38370 17320 38426 17354
rect 38460 17320 38516 17354
rect 38550 17320 38606 17354
rect 38640 17320 38696 17354
rect 38730 17320 38786 17354
rect 38820 17320 38954 17354
rect 28286 17288 38954 17320
rect 23948 17255 26824 17262
rect 23948 17221 23949 17255
rect 23983 17221 26824 17255
rect 23948 17202 26824 17221
rect 23948 17153 26824 17156
rect 23948 17143 26525 17153
rect 26559 17143 26824 17153
rect 23948 17109 24131 17143
rect 24165 17109 24531 17143
rect 24565 17109 24931 17143
rect 24965 17109 25331 17143
rect 25365 17109 25731 17143
rect 25765 17109 26131 17143
rect 26165 17119 26525 17143
rect 26165 17109 26531 17119
rect 26565 17109 26824 17143
rect 23948 17096 26824 17109
rect 40168 17022 40784 17821
rect 41264 17677 41696 18067
rect 5916 17009 10194 17022
rect 5916 16975 6197 17009
rect 6231 16975 6597 17009
rect 6631 16975 6997 17009
rect 7031 16975 7397 17009
rect 7431 16975 7797 17009
rect 7831 16975 8197 17009
rect 8231 16975 8597 17009
rect 8631 16975 8997 17009
rect 9031 16975 9397 17009
rect 9431 16975 9797 17009
rect 9831 16975 10194 17009
rect 5916 16962 10194 16975
rect 10640 17009 13080 17022
rect 10640 16975 10823 17009
rect 10857 16975 11023 17009
rect 11057 16975 11223 17009
rect 11257 16975 11423 17009
rect 11457 16975 11623 17009
rect 11657 16975 11823 17009
rect 11857 16975 12023 17009
rect 12057 16975 12223 17009
rect 12257 16975 12423 17009
rect 12457 16975 12623 17009
rect 12657 16975 12823 17009
rect 12857 16975 13080 17009
rect 10640 16962 13080 16975
rect 13384 17009 15824 17022
rect 13384 16975 13567 17009
rect 13601 16975 13767 17009
rect 13801 16975 13967 17009
rect 14001 16975 14167 17009
rect 14201 16975 14367 17009
rect 14401 16975 14567 17009
rect 14601 16975 14767 17009
rect 14801 16975 14967 17009
rect 15001 16975 15167 17009
rect 15201 16975 15367 17009
rect 15401 16975 15567 17009
rect 15601 16975 15824 17009
rect 13384 16962 15824 16975
rect 16110 17009 23278 17022
rect 16110 16975 16293 17009
rect 16327 16975 16693 17009
rect 16727 16975 17093 17009
rect 17127 16975 17493 17009
rect 17527 16975 17893 17009
rect 17927 16975 18293 17009
rect 18327 16975 18693 17009
rect 18727 16975 19093 17009
rect 19127 16975 19493 17009
rect 19527 16975 19893 17009
rect 19927 16975 20293 17009
rect 20327 16975 20693 17009
rect 20727 16975 21093 17009
rect 21127 16975 21493 17009
rect 21527 16975 21893 17009
rect 21927 16975 22293 17009
rect 22327 16975 22693 17009
rect 22727 16975 23093 17009
rect 23127 16975 23278 17009
rect 16110 16962 23278 16975
rect 23850 17009 26824 17022
rect 23850 16975 24131 17009
rect 24165 16975 24531 17009
rect 24565 16975 24931 17009
rect 24965 16975 25331 17009
rect 25365 16975 25731 17009
rect 25765 16975 26131 17009
rect 26165 16975 26531 17009
rect 26565 16975 26824 17009
rect 23850 16962 26824 16975
rect 28260 17009 38980 17022
rect 28260 16975 28443 17009
rect 28477 16975 28643 17009
rect 28677 16975 28843 17009
rect 28877 16975 29043 17009
rect 29077 16975 29243 17009
rect 29277 16975 29443 17009
rect 29477 16975 29643 17009
rect 29677 16975 29843 17009
rect 29877 16975 30043 17009
rect 30077 16975 30243 17009
rect 30277 16975 30443 17009
rect 30477 16975 30643 17009
rect 30677 16975 30843 17009
rect 30877 16975 31043 17009
rect 31077 16975 31243 17009
rect 31277 16975 31443 17009
rect 31477 16975 31643 17009
rect 31677 16975 31843 17009
rect 31877 16975 32043 17009
rect 32077 16975 32243 17009
rect 32277 16975 32443 17009
rect 32477 16975 32643 17009
rect 32677 16975 32843 17009
rect 32877 16975 33043 17009
rect 33077 16975 33243 17009
rect 33277 16975 33443 17009
rect 33477 16975 33643 17009
rect 33677 16975 33843 17009
rect 33877 16975 34043 17009
rect 34077 16975 34243 17009
rect 34277 16975 34443 17009
rect 34477 16975 34643 17009
rect 34677 16975 34843 17009
rect 34877 16975 35043 17009
rect 35077 16975 35243 17009
rect 35277 16975 35443 17009
rect 35477 16975 35643 17009
rect 35677 16975 35843 17009
rect 35877 16975 36043 17009
rect 36077 16975 36243 17009
rect 36277 16975 36443 17009
rect 36477 16975 36643 17009
rect 36677 16975 36843 17009
rect 36877 16975 37043 17009
rect 37077 16975 37243 17009
rect 37277 16975 37443 17009
rect 37477 16975 37643 17009
rect 37677 16975 37843 17009
rect 37877 16975 38043 17009
rect 38077 16975 38243 17009
rect 38277 16975 38443 17009
rect 38477 16975 38643 17009
rect 38677 16975 38843 17009
rect 38877 16975 38980 17009
rect 28260 16962 38980 16975
rect 39256 17009 41696 17022
rect 39256 16975 39439 17009
rect 39473 16975 39639 17009
rect 39673 16975 39839 17009
rect 39873 16975 40039 17009
rect 40073 16975 40239 17009
rect 40273 16975 40439 17009
rect 40473 16975 40639 17009
rect 40673 16975 40839 17009
rect 40873 16975 41039 17009
rect 41073 16975 41239 17009
rect 41273 16975 41439 17009
rect 41473 16975 41696 17009
rect 39256 16962 41696 16975
rect 7896 15129 10336 15142
rect 7896 15095 8079 15129
rect 8113 15095 8279 15129
rect 8313 15095 8479 15129
rect 8513 15095 8679 15129
rect 8713 15095 8879 15129
rect 8913 15095 9079 15129
rect 9113 15095 9279 15129
rect 9313 15095 9479 15129
rect 9513 15095 9679 15129
rect 9713 15095 9879 15129
rect 9913 15095 10079 15129
rect 10113 15095 10336 15129
rect 7896 15082 10336 15095
rect 10640 15129 13080 15142
rect 10640 15095 10823 15129
rect 10857 15095 11023 15129
rect 11057 15095 11223 15129
rect 11257 15095 11423 15129
rect 11457 15095 11623 15129
rect 11657 15095 11823 15129
rect 11857 15095 12023 15129
rect 12057 15095 12223 15129
rect 12257 15095 12423 15129
rect 12457 15095 12623 15129
rect 12657 15095 12823 15129
rect 12857 15095 13080 15129
rect 10640 15082 13080 15095
rect 13384 15129 15824 15142
rect 13384 15095 13567 15129
rect 13601 15095 13767 15129
rect 13801 15095 13967 15129
rect 14001 15095 14167 15129
rect 14201 15095 14367 15129
rect 14401 15095 14567 15129
rect 14601 15095 14767 15129
rect 14801 15095 14967 15129
rect 15001 15095 15167 15129
rect 15201 15095 15367 15129
rect 15401 15095 15567 15129
rect 15601 15095 15824 15129
rect 13384 15082 15824 15095
rect 16110 15129 23278 15142
rect 16110 15095 16293 15129
rect 16327 15095 16693 15129
rect 16727 15095 17093 15129
rect 17127 15095 17493 15129
rect 17527 15095 17893 15129
rect 17927 15095 18293 15129
rect 18327 15095 18693 15129
rect 18727 15095 19093 15129
rect 19127 15095 19493 15129
rect 19527 15095 19893 15129
rect 19927 15095 20293 15129
rect 20327 15095 20693 15129
rect 20727 15095 21093 15129
rect 21127 15095 21493 15129
rect 21527 15095 21893 15129
rect 21927 15095 22293 15129
rect 22327 15095 22693 15129
rect 22727 15095 23093 15129
rect 23127 15095 23278 15129
rect 16110 15082 23278 15095
rect 23576 15129 26016 15142
rect 23576 15095 23759 15129
rect 23793 15095 23959 15129
rect 23993 15095 24159 15129
rect 24193 15095 24359 15129
rect 24393 15095 24559 15129
rect 24593 15095 24759 15129
rect 24793 15095 24959 15129
rect 24993 15095 25159 15129
rect 25193 15095 25359 15129
rect 25393 15095 25559 15129
rect 25593 15095 25759 15129
rect 25793 15095 26016 15129
rect 23576 15082 26016 15095
rect 28260 15129 38980 15142
rect 28260 15095 28443 15129
rect 28477 15095 28643 15129
rect 28677 15095 28843 15129
rect 28877 15095 29043 15129
rect 29077 15095 29243 15129
rect 29277 15095 29443 15129
rect 29477 15095 29643 15129
rect 29677 15095 29843 15129
rect 29877 15095 30043 15129
rect 30077 15095 30243 15129
rect 30277 15095 30443 15129
rect 30477 15095 30643 15129
rect 30677 15095 30843 15129
rect 30877 15095 31043 15129
rect 31077 15095 31243 15129
rect 31277 15095 31443 15129
rect 31477 15095 31643 15129
rect 31677 15095 31843 15129
rect 31877 15095 32043 15129
rect 32077 15095 32243 15129
rect 32277 15095 32443 15129
rect 32477 15095 32643 15129
rect 32677 15095 32843 15129
rect 32877 15095 33043 15129
rect 33077 15095 33243 15129
rect 33277 15095 33443 15129
rect 33477 15095 33643 15129
rect 33677 15095 33843 15129
rect 33877 15095 34043 15129
rect 34077 15095 34243 15129
rect 34277 15095 34443 15129
rect 34477 15095 34643 15129
rect 34677 15095 34843 15129
rect 34877 15095 35043 15129
rect 35077 15095 35243 15129
rect 35277 15095 35443 15129
rect 35477 15095 35643 15129
rect 35677 15095 35843 15129
rect 35877 15095 36043 15129
rect 36077 15095 36243 15129
rect 36277 15095 36443 15129
rect 36477 15095 36643 15129
rect 36677 15095 36843 15129
rect 36877 15095 37043 15129
rect 37077 15095 37243 15129
rect 37277 15095 37443 15129
rect 37477 15095 37643 15129
rect 37677 15095 37843 15129
rect 37877 15095 38043 15129
rect 38077 15095 38243 15129
rect 38277 15095 38443 15129
rect 38477 15095 38643 15129
rect 38677 15095 38843 15129
rect 38877 15095 38980 15129
rect 28260 15082 38980 15095
rect 39256 15129 41696 15142
rect 39256 15095 39439 15129
rect 39473 15095 39639 15129
rect 39673 15095 39839 15129
rect 39873 15095 40039 15129
rect 40073 15095 40239 15129
rect 40273 15095 40439 15129
rect 40473 15095 40639 15129
rect 40673 15095 40839 15129
rect 40873 15095 41039 15129
rect 41073 15095 41239 15129
rect 41273 15095 41439 15129
rect 41473 15095 41696 15129
rect 39256 15082 41696 15095
rect 8808 14163 9424 14202
rect 8808 14061 8895 14163
rect 9337 14061 9424 14163
rect 8808 13262 9424 14061
rect 9904 13917 10336 14307
rect 11552 14163 12168 14202
rect 11552 14061 11639 14163
rect 12081 14061 12168 14163
rect 11552 13262 12168 14061
rect 12648 13917 13080 14307
rect 14296 14163 14912 14202
rect 14296 14061 14383 14163
rect 14825 14061 14912 14163
rect 14296 13262 14912 14061
rect 15392 13917 15824 14307
rect 24488 14163 25104 14202
rect 24488 14061 24575 14163
rect 25017 14061 25104 14163
rect 24488 13262 25104 14061
rect 25584 13917 26016 14307
rect 28286 14796 38954 14816
rect 28286 14762 28306 14796
rect 28340 14762 28396 14796
rect 28430 14781 28486 14796
rect 28520 14781 28576 14796
rect 28610 14781 28666 14796
rect 28700 14781 28756 14796
rect 28790 14781 28846 14796
rect 28880 14781 28936 14796
rect 28970 14781 29026 14796
rect 29060 14781 29116 14796
rect 29150 14781 29206 14796
rect 29240 14781 29296 14796
rect 29330 14781 29386 14796
rect 29420 14781 29476 14796
rect 28450 14762 28486 14781
rect 28540 14762 28576 14781
rect 28630 14762 28666 14781
rect 28720 14762 28756 14781
rect 28810 14762 28846 14781
rect 28900 14762 28936 14781
rect 28990 14762 29026 14781
rect 29080 14762 29116 14781
rect 29170 14762 29206 14781
rect 29260 14762 29296 14781
rect 29350 14762 29386 14781
rect 29440 14762 29476 14781
rect 29510 14762 29646 14796
rect 29680 14762 29736 14796
rect 29770 14781 29826 14796
rect 29860 14781 29916 14796
rect 29950 14781 30006 14796
rect 30040 14781 30096 14796
rect 30130 14781 30186 14796
rect 30220 14781 30276 14796
rect 30310 14781 30366 14796
rect 30400 14781 30456 14796
rect 30490 14781 30546 14796
rect 30580 14781 30636 14796
rect 30670 14781 30726 14796
rect 30760 14781 30816 14796
rect 29790 14762 29826 14781
rect 29880 14762 29916 14781
rect 29970 14762 30006 14781
rect 30060 14762 30096 14781
rect 30150 14762 30186 14781
rect 30240 14762 30276 14781
rect 30330 14762 30366 14781
rect 30420 14762 30456 14781
rect 30510 14762 30546 14781
rect 30600 14762 30636 14781
rect 30690 14762 30726 14781
rect 30780 14762 30816 14781
rect 30850 14762 30986 14796
rect 31020 14762 31076 14796
rect 31110 14781 31166 14796
rect 31200 14781 31256 14796
rect 31290 14781 31346 14796
rect 31380 14781 31436 14796
rect 31470 14781 31526 14796
rect 31560 14781 31616 14796
rect 31650 14781 31706 14796
rect 31740 14781 31796 14796
rect 31830 14781 31886 14796
rect 31920 14781 31976 14796
rect 32010 14781 32066 14796
rect 32100 14781 32156 14796
rect 31130 14762 31166 14781
rect 31220 14762 31256 14781
rect 31310 14762 31346 14781
rect 31400 14762 31436 14781
rect 31490 14762 31526 14781
rect 31580 14762 31616 14781
rect 31670 14762 31706 14781
rect 31760 14762 31796 14781
rect 31850 14762 31886 14781
rect 31940 14762 31976 14781
rect 32030 14762 32066 14781
rect 32120 14762 32156 14781
rect 32190 14762 32326 14796
rect 32360 14762 32416 14796
rect 32450 14781 32506 14796
rect 32540 14781 32596 14796
rect 32630 14781 32686 14796
rect 32720 14781 32776 14796
rect 32810 14781 32866 14796
rect 32900 14781 32956 14796
rect 32990 14781 33046 14796
rect 33080 14781 33136 14796
rect 33170 14781 33226 14796
rect 33260 14781 33316 14796
rect 33350 14781 33406 14796
rect 33440 14781 33496 14796
rect 32470 14762 32506 14781
rect 32560 14762 32596 14781
rect 32650 14762 32686 14781
rect 32740 14762 32776 14781
rect 32830 14762 32866 14781
rect 32920 14762 32956 14781
rect 33010 14762 33046 14781
rect 33100 14762 33136 14781
rect 33190 14762 33226 14781
rect 33280 14762 33316 14781
rect 33370 14762 33406 14781
rect 33460 14762 33496 14781
rect 33530 14762 33666 14796
rect 33700 14762 33756 14796
rect 33790 14781 33846 14796
rect 33880 14781 33936 14796
rect 33970 14781 34026 14796
rect 34060 14781 34116 14796
rect 34150 14781 34206 14796
rect 34240 14781 34296 14796
rect 34330 14781 34386 14796
rect 34420 14781 34476 14796
rect 34510 14781 34566 14796
rect 34600 14781 34656 14796
rect 34690 14781 34746 14796
rect 34780 14781 34836 14796
rect 33810 14762 33846 14781
rect 33900 14762 33936 14781
rect 33990 14762 34026 14781
rect 34080 14762 34116 14781
rect 34170 14762 34206 14781
rect 34260 14762 34296 14781
rect 34350 14762 34386 14781
rect 34440 14762 34476 14781
rect 34530 14762 34566 14781
rect 34620 14762 34656 14781
rect 34710 14762 34746 14781
rect 34800 14762 34836 14781
rect 34870 14762 35006 14796
rect 35040 14762 35096 14796
rect 35130 14781 35186 14796
rect 35220 14781 35276 14796
rect 35310 14781 35366 14796
rect 35400 14781 35456 14796
rect 35490 14781 35546 14796
rect 35580 14781 35636 14796
rect 35670 14781 35726 14796
rect 35760 14781 35816 14796
rect 35850 14781 35906 14796
rect 35940 14781 35996 14796
rect 36030 14781 36086 14796
rect 36120 14781 36176 14796
rect 35150 14762 35186 14781
rect 35240 14762 35276 14781
rect 35330 14762 35366 14781
rect 35420 14762 35456 14781
rect 35510 14762 35546 14781
rect 35600 14762 35636 14781
rect 35690 14762 35726 14781
rect 35780 14762 35816 14781
rect 35870 14762 35906 14781
rect 35960 14762 35996 14781
rect 36050 14762 36086 14781
rect 36140 14762 36176 14781
rect 36210 14762 36346 14796
rect 36380 14762 36436 14796
rect 36470 14781 36526 14796
rect 36560 14781 36616 14796
rect 36650 14781 36706 14796
rect 36740 14781 36796 14796
rect 36830 14781 36886 14796
rect 36920 14781 36976 14796
rect 37010 14781 37066 14796
rect 37100 14781 37156 14796
rect 37190 14781 37246 14796
rect 37280 14781 37336 14796
rect 37370 14781 37426 14796
rect 37460 14781 37516 14796
rect 36490 14762 36526 14781
rect 36580 14762 36616 14781
rect 36670 14762 36706 14781
rect 36760 14762 36796 14781
rect 36850 14762 36886 14781
rect 36940 14762 36976 14781
rect 37030 14762 37066 14781
rect 37120 14762 37156 14781
rect 37210 14762 37246 14781
rect 37300 14762 37336 14781
rect 37390 14762 37426 14781
rect 37480 14762 37516 14781
rect 37550 14762 37686 14796
rect 37720 14762 37776 14796
rect 37810 14781 37866 14796
rect 37900 14781 37956 14796
rect 37990 14781 38046 14796
rect 38080 14781 38136 14796
rect 38170 14781 38226 14796
rect 38260 14781 38316 14796
rect 38350 14781 38406 14796
rect 38440 14781 38496 14796
rect 38530 14781 38586 14796
rect 38620 14781 38676 14796
rect 38710 14781 38766 14796
rect 38800 14781 38856 14796
rect 37830 14762 37866 14781
rect 37920 14762 37956 14781
rect 38010 14762 38046 14781
rect 38100 14762 38136 14781
rect 38190 14762 38226 14781
rect 38280 14762 38316 14781
rect 38370 14762 38406 14781
rect 38460 14762 38496 14781
rect 38550 14762 38586 14781
rect 38640 14762 38676 14781
rect 38730 14762 38766 14781
rect 38820 14762 38856 14781
rect 38890 14762 38954 14796
rect 28286 14758 28416 14762
rect 28286 14724 28320 14758
rect 28354 14747 28416 14758
rect 28450 14747 28506 14762
rect 28540 14747 28596 14762
rect 28630 14747 28686 14762
rect 28720 14747 28776 14762
rect 28810 14747 28866 14762
rect 28900 14747 28956 14762
rect 28990 14747 29046 14762
rect 29080 14747 29136 14762
rect 29170 14747 29226 14762
rect 29260 14747 29316 14762
rect 29350 14747 29406 14762
rect 29440 14758 29756 14762
rect 29440 14747 29507 14758
rect 28354 14724 29507 14747
rect 29541 14724 29660 14758
rect 29694 14747 29756 14758
rect 29790 14747 29846 14762
rect 29880 14747 29936 14762
rect 29970 14747 30026 14762
rect 30060 14747 30116 14762
rect 30150 14747 30206 14762
rect 30240 14747 30296 14762
rect 30330 14747 30386 14762
rect 30420 14747 30476 14762
rect 30510 14747 30566 14762
rect 30600 14747 30656 14762
rect 30690 14747 30746 14762
rect 30780 14758 31096 14762
rect 30780 14747 30847 14758
rect 29694 14724 30847 14747
rect 30881 14724 31000 14758
rect 31034 14747 31096 14758
rect 31130 14747 31186 14762
rect 31220 14747 31276 14762
rect 31310 14747 31366 14762
rect 31400 14747 31456 14762
rect 31490 14747 31546 14762
rect 31580 14747 31636 14762
rect 31670 14747 31726 14762
rect 31760 14747 31816 14762
rect 31850 14747 31906 14762
rect 31940 14747 31996 14762
rect 32030 14747 32086 14762
rect 32120 14758 32436 14762
rect 32120 14747 32187 14758
rect 31034 14724 32187 14747
rect 32221 14724 32340 14758
rect 32374 14747 32436 14758
rect 32470 14747 32526 14762
rect 32560 14747 32616 14762
rect 32650 14747 32706 14762
rect 32740 14747 32796 14762
rect 32830 14747 32886 14762
rect 32920 14747 32976 14762
rect 33010 14747 33066 14762
rect 33100 14747 33156 14762
rect 33190 14747 33246 14762
rect 33280 14747 33336 14762
rect 33370 14747 33426 14762
rect 33460 14758 33776 14762
rect 33460 14747 33527 14758
rect 32374 14724 33527 14747
rect 33561 14724 33680 14758
rect 33714 14747 33776 14758
rect 33810 14747 33866 14762
rect 33900 14747 33956 14762
rect 33990 14747 34046 14762
rect 34080 14747 34136 14762
rect 34170 14747 34226 14762
rect 34260 14747 34316 14762
rect 34350 14747 34406 14762
rect 34440 14747 34496 14762
rect 34530 14747 34586 14762
rect 34620 14747 34676 14762
rect 34710 14747 34766 14762
rect 34800 14758 35116 14762
rect 34800 14747 34867 14758
rect 33714 14724 34867 14747
rect 34901 14724 35020 14758
rect 35054 14747 35116 14758
rect 35150 14747 35206 14762
rect 35240 14747 35296 14762
rect 35330 14747 35386 14762
rect 35420 14747 35476 14762
rect 35510 14747 35566 14762
rect 35600 14747 35656 14762
rect 35690 14747 35746 14762
rect 35780 14747 35836 14762
rect 35870 14747 35926 14762
rect 35960 14747 36016 14762
rect 36050 14747 36106 14762
rect 36140 14758 36456 14762
rect 36140 14747 36207 14758
rect 35054 14724 36207 14747
rect 36241 14724 36360 14758
rect 36394 14747 36456 14758
rect 36490 14747 36546 14762
rect 36580 14747 36636 14762
rect 36670 14747 36726 14762
rect 36760 14747 36816 14762
rect 36850 14747 36906 14762
rect 36940 14747 36996 14762
rect 37030 14747 37086 14762
rect 37120 14747 37176 14762
rect 37210 14747 37266 14762
rect 37300 14747 37356 14762
rect 37390 14747 37446 14762
rect 37480 14758 37796 14762
rect 37480 14747 37547 14758
rect 36394 14724 37547 14747
rect 37581 14724 37700 14758
rect 37734 14747 37796 14758
rect 37830 14747 37886 14762
rect 37920 14747 37976 14762
rect 38010 14747 38066 14762
rect 38100 14747 38156 14762
rect 38190 14747 38246 14762
rect 38280 14747 38336 14762
rect 38370 14747 38426 14762
rect 38460 14747 38516 14762
rect 38550 14747 38606 14762
rect 38640 14747 38696 14762
rect 38730 14747 38786 14762
rect 38820 14758 38954 14762
rect 38820 14747 38887 14758
rect 37734 14724 38887 14747
rect 38921 14724 38954 14758
rect 28286 14717 38954 14724
rect 28286 14668 28385 14717
rect 28286 14634 28320 14668
rect 28354 14634 28385 14668
rect 29475 14668 29725 14717
rect 28286 14578 28385 14634
rect 28286 14544 28320 14578
rect 28354 14544 28385 14578
rect 28286 14488 28385 14544
rect 28286 14454 28320 14488
rect 28354 14454 28385 14488
rect 28286 14398 28385 14454
rect 28286 14364 28320 14398
rect 28354 14364 28385 14398
rect 28286 14308 28385 14364
rect 28286 14274 28320 14308
rect 28354 14274 28385 14308
rect 28286 14218 28385 14274
rect 28286 14184 28320 14218
rect 28354 14184 28385 14218
rect 28286 14128 28385 14184
rect 28286 14094 28320 14128
rect 28354 14094 28385 14128
rect 28286 14038 28385 14094
rect 28286 14004 28320 14038
rect 28354 14004 28385 14038
rect 28286 13948 28385 14004
rect 28286 13914 28320 13948
rect 28354 13914 28385 13948
rect 28286 13858 28385 13914
rect 28286 13824 28320 13858
rect 28354 13824 28385 13858
rect 28286 13768 28385 13824
rect 28286 13734 28320 13768
rect 28354 13734 28385 13768
rect 28286 13678 28385 13734
rect 28449 14636 29411 14653
rect 28449 14602 28470 14636
rect 28504 14602 28560 14636
rect 28594 14634 28650 14636
rect 28684 14634 28740 14636
rect 28774 14634 28830 14636
rect 28864 14634 28920 14636
rect 28954 14634 29010 14636
rect 29044 14634 29100 14636
rect 29134 14634 29190 14636
rect 29224 14634 29280 14636
rect 29314 14634 29370 14636
rect 28614 14602 28650 14634
rect 28704 14602 28740 14634
rect 28794 14602 28830 14634
rect 28884 14602 28920 14634
rect 28974 14602 29010 14634
rect 29064 14602 29100 14634
rect 29154 14602 29190 14634
rect 29244 14602 29280 14634
rect 29334 14602 29370 14634
rect 29404 14602 29411 14636
rect 28449 14600 28580 14602
rect 28614 14600 28670 14602
rect 28704 14600 28760 14602
rect 28794 14600 28850 14602
rect 28884 14600 28940 14602
rect 28974 14600 29030 14602
rect 29064 14600 29120 14602
rect 29154 14600 29210 14602
rect 29244 14600 29300 14602
rect 29334 14600 29411 14602
rect 28449 14581 29411 14600
rect 28449 14577 28521 14581
rect 28449 14543 28468 14577
rect 28502 14543 28521 14577
rect 28449 14487 28521 14543
rect 29339 14558 29411 14581
rect 29339 14524 29358 14558
rect 29392 14524 29411 14558
rect 28449 14453 28468 14487
rect 28502 14453 28521 14487
rect 28449 14397 28521 14453
rect 28449 14363 28468 14397
rect 28502 14363 28521 14397
rect 28449 14307 28521 14363
rect 28449 14273 28468 14307
rect 28502 14273 28521 14307
rect 28449 14217 28521 14273
rect 28449 14183 28468 14217
rect 28502 14183 28521 14217
rect 28449 14127 28521 14183
rect 28449 14093 28468 14127
rect 28502 14093 28521 14127
rect 28449 14037 28521 14093
rect 28449 14003 28468 14037
rect 28502 14003 28521 14037
rect 28449 13947 28521 14003
rect 28449 13913 28468 13947
rect 28502 13913 28521 13947
rect 28449 13857 28521 13913
rect 28449 13823 28468 13857
rect 28502 13823 28521 13857
rect 28583 14460 29277 14519
rect 28583 14426 28644 14460
rect 28678 14432 28734 14460
rect 28768 14432 28824 14460
rect 28858 14432 28914 14460
rect 28690 14426 28734 14432
rect 28790 14426 28824 14432
rect 28890 14426 28914 14432
rect 28948 14432 29004 14460
rect 28948 14426 28956 14432
rect 28583 14398 28656 14426
rect 28690 14398 28756 14426
rect 28790 14398 28856 14426
rect 28890 14398 28956 14426
rect 28990 14426 29004 14432
rect 29038 14432 29094 14460
rect 29038 14426 29056 14432
rect 28990 14398 29056 14426
rect 29090 14426 29094 14432
rect 29128 14432 29184 14460
rect 29128 14426 29156 14432
rect 29218 14426 29277 14460
rect 29090 14398 29156 14426
rect 29190 14398 29277 14426
rect 28583 14370 29277 14398
rect 28583 14336 28644 14370
rect 28678 14336 28734 14370
rect 28768 14336 28824 14370
rect 28858 14336 28914 14370
rect 28948 14336 29004 14370
rect 29038 14336 29094 14370
rect 29128 14336 29184 14370
rect 29218 14336 29277 14370
rect 28583 14332 29277 14336
rect 28583 14298 28656 14332
rect 28690 14298 28756 14332
rect 28790 14298 28856 14332
rect 28890 14298 28956 14332
rect 28990 14298 29056 14332
rect 29090 14298 29156 14332
rect 29190 14298 29277 14332
rect 28583 14280 29277 14298
rect 28583 14246 28644 14280
rect 28678 14246 28734 14280
rect 28768 14246 28824 14280
rect 28858 14246 28914 14280
rect 28948 14246 29004 14280
rect 29038 14246 29094 14280
rect 29128 14246 29184 14280
rect 29218 14246 29277 14280
rect 28583 14232 29277 14246
rect 28583 14198 28656 14232
rect 28690 14198 28756 14232
rect 28790 14198 28856 14232
rect 28890 14198 28956 14232
rect 28990 14198 29056 14232
rect 29090 14198 29156 14232
rect 29190 14198 29277 14232
rect 28583 14190 29277 14198
rect 28583 14156 28644 14190
rect 28678 14156 28734 14190
rect 28768 14156 28824 14190
rect 28858 14156 28914 14190
rect 28948 14156 29004 14190
rect 29038 14156 29094 14190
rect 29128 14156 29184 14190
rect 29218 14156 29277 14190
rect 28583 14132 29277 14156
rect 28583 14100 28656 14132
rect 28690 14100 28756 14132
rect 28790 14100 28856 14132
rect 28890 14100 28956 14132
rect 28583 14066 28644 14100
rect 28690 14098 28734 14100
rect 28790 14098 28824 14100
rect 28890 14098 28914 14100
rect 28678 14066 28734 14098
rect 28768 14066 28824 14098
rect 28858 14066 28914 14098
rect 28948 14098 28956 14100
rect 28990 14100 29056 14132
rect 28990 14098 29004 14100
rect 28948 14066 29004 14098
rect 29038 14098 29056 14100
rect 29090 14100 29156 14132
rect 29190 14100 29277 14132
rect 29090 14098 29094 14100
rect 29038 14066 29094 14098
rect 29128 14098 29156 14100
rect 29128 14066 29184 14098
rect 29218 14066 29277 14100
rect 28583 14032 29277 14066
rect 28583 14010 28656 14032
rect 28690 14010 28756 14032
rect 28790 14010 28856 14032
rect 28890 14010 28956 14032
rect 28583 13976 28644 14010
rect 28690 13998 28734 14010
rect 28790 13998 28824 14010
rect 28890 13998 28914 14010
rect 28678 13976 28734 13998
rect 28768 13976 28824 13998
rect 28858 13976 28914 13998
rect 28948 13998 28956 14010
rect 28990 14010 29056 14032
rect 28990 13998 29004 14010
rect 28948 13976 29004 13998
rect 29038 13998 29056 14010
rect 29090 14010 29156 14032
rect 29190 14010 29277 14032
rect 29090 13998 29094 14010
rect 29038 13976 29094 13998
rect 29128 13998 29156 14010
rect 29128 13976 29184 13998
rect 29218 13976 29277 14010
rect 28583 13932 29277 13976
rect 28583 13920 28656 13932
rect 28690 13920 28756 13932
rect 28790 13920 28856 13932
rect 28890 13920 28956 13932
rect 28583 13886 28644 13920
rect 28690 13898 28734 13920
rect 28790 13898 28824 13920
rect 28890 13898 28914 13920
rect 28678 13886 28734 13898
rect 28768 13886 28824 13898
rect 28858 13886 28914 13898
rect 28948 13898 28956 13920
rect 28990 13920 29056 13932
rect 28990 13898 29004 13920
rect 28948 13886 29004 13898
rect 29038 13898 29056 13920
rect 29090 13920 29156 13932
rect 29190 13920 29277 13932
rect 29090 13898 29094 13920
rect 29038 13886 29094 13898
rect 29128 13898 29156 13920
rect 29128 13886 29184 13898
rect 29218 13886 29277 13920
rect 28583 13825 29277 13886
rect 29339 14468 29411 14524
rect 29339 14434 29358 14468
rect 29392 14434 29411 14468
rect 29339 14378 29411 14434
rect 29339 14344 29358 14378
rect 29392 14344 29411 14378
rect 29339 14288 29411 14344
rect 29339 14254 29358 14288
rect 29392 14254 29411 14288
rect 29339 14198 29411 14254
rect 29339 14164 29358 14198
rect 29392 14164 29411 14198
rect 29339 14108 29411 14164
rect 29339 14074 29358 14108
rect 29392 14074 29411 14108
rect 29339 14018 29411 14074
rect 29339 13984 29358 14018
rect 29392 13984 29411 14018
rect 29339 13928 29411 13984
rect 29339 13894 29358 13928
rect 29392 13894 29411 13928
rect 29339 13838 29411 13894
rect 28449 13763 28521 13823
rect 29339 13804 29358 13838
rect 29392 13804 29411 13838
rect 29339 13763 29411 13804
rect 28449 13744 29411 13763
rect 28449 13710 28546 13744
rect 28580 13710 28636 13744
rect 28670 13710 28726 13744
rect 28760 13710 28816 13744
rect 28850 13710 28906 13744
rect 28940 13710 28996 13744
rect 29030 13710 29086 13744
rect 29120 13710 29176 13744
rect 29210 13710 29266 13744
rect 29300 13710 29411 13744
rect 28449 13691 29411 13710
rect 29475 14634 29507 14668
rect 29541 14634 29660 14668
rect 29694 14634 29725 14668
rect 30815 14668 31065 14717
rect 29475 14578 29725 14634
rect 29475 14544 29507 14578
rect 29541 14544 29660 14578
rect 29694 14544 29725 14578
rect 29475 14488 29725 14544
rect 29475 14454 29507 14488
rect 29541 14454 29660 14488
rect 29694 14454 29725 14488
rect 29475 14398 29725 14454
rect 29475 14364 29507 14398
rect 29541 14364 29660 14398
rect 29694 14364 29725 14398
rect 29475 14308 29725 14364
rect 29475 14274 29507 14308
rect 29541 14274 29660 14308
rect 29694 14274 29725 14308
rect 29475 14218 29725 14274
rect 29475 14184 29507 14218
rect 29541 14184 29660 14218
rect 29694 14184 29725 14218
rect 29475 14128 29725 14184
rect 29475 14094 29507 14128
rect 29541 14094 29660 14128
rect 29694 14094 29725 14128
rect 29475 14038 29725 14094
rect 29475 14004 29507 14038
rect 29541 14004 29660 14038
rect 29694 14004 29725 14038
rect 29475 13948 29725 14004
rect 29475 13914 29507 13948
rect 29541 13914 29660 13948
rect 29694 13914 29725 13948
rect 29475 13858 29725 13914
rect 29475 13824 29507 13858
rect 29541 13824 29660 13858
rect 29694 13824 29725 13858
rect 29475 13768 29725 13824
rect 29475 13734 29507 13768
rect 29541 13734 29660 13768
rect 29694 13734 29725 13768
rect 28286 13644 28320 13678
rect 28354 13644 28385 13678
rect 28286 13627 28385 13644
rect 29475 13678 29725 13734
rect 29789 14636 30751 14653
rect 29789 14602 29810 14636
rect 29844 14602 29900 14636
rect 29934 14634 29990 14636
rect 30024 14634 30080 14636
rect 30114 14634 30170 14636
rect 30204 14634 30260 14636
rect 30294 14634 30350 14636
rect 30384 14634 30440 14636
rect 30474 14634 30530 14636
rect 30564 14634 30620 14636
rect 30654 14634 30710 14636
rect 29954 14602 29990 14634
rect 30044 14602 30080 14634
rect 30134 14602 30170 14634
rect 30224 14602 30260 14634
rect 30314 14602 30350 14634
rect 30404 14602 30440 14634
rect 30494 14602 30530 14634
rect 30584 14602 30620 14634
rect 30674 14602 30710 14634
rect 30744 14602 30751 14636
rect 29789 14600 29920 14602
rect 29954 14600 30010 14602
rect 30044 14600 30100 14602
rect 30134 14600 30190 14602
rect 30224 14600 30280 14602
rect 30314 14600 30370 14602
rect 30404 14600 30460 14602
rect 30494 14600 30550 14602
rect 30584 14600 30640 14602
rect 30674 14600 30751 14602
rect 29789 14581 30751 14600
rect 29789 14577 29861 14581
rect 29789 14543 29808 14577
rect 29842 14543 29861 14577
rect 29789 14487 29861 14543
rect 30679 14558 30751 14581
rect 30679 14524 30698 14558
rect 30732 14524 30751 14558
rect 29789 14453 29808 14487
rect 29842 14453 29861 14487
rect 29789 14397 29861 14453
rect 29789 14363 29808 14397
rect 29842 14363 29861 14397
rect 29789 14307 29861 14363
rect 29789 14273 29808 14307
rect 29842 14273 29861 14307
rect 29789 14217 29861 14273
rect 29789 14183 29808 14217
rect 29842 14183 29861 14217
rect 29789 14127 29861 14183
rect 29789 14093 29808 14127
rect 29842 14093 29861 14127
rect 29789 14037 29861 14093
rect 29789 14003 29808 14037
rect 29842 14003 29861 14037
rect 29789 13947 29861 14003
rect 29789 13913 29808 13947
rect 29842 13913 29861 13947
rect 29789 13857 29861 13913
rect 29789 13823 29808 13857
rect 29842 13823 29861 13857
rect 29923 14460 30617 14519
rect 29923 14426 29984 14460
rect 30018 14432 30074 14460
rect 30108 14432 30164 14460
rect 30198 14432 30254 14460
rect 30030 14426 30074 14432
rect 30130 14426 30164 14432
rect 30230 14426 30254 14432
rect 30288 14432 30344 14460
rect 30288 14426 30296 14432
rect 29923 14398 29996 14426
rect 30030 14398 30096 14426
rect 30130 14398 30196 14426
rect 30230 14398 30296 14426
rect 30330 14426 30344 14432
rect 30378 14432 30434 14460
rect 30378 14426 30396 14432
rect 30330 14398 30396 14426
rect 30430 14426 30434 14432
rect 30468 14432 30524 14460
rect 30468 14426 30496 14432
rect 30558 14426 30617 14460
rect 30430 14398 30496 14426
rect 30530 14398 30617 14426
rect 29923 14370 30617 14398
rect 29923 14336 29984 14370
rect 30018 14336 30074 14370
rect 30108 14336 30164 14370
rect 30198 14336 30254 14370
rect 30288 14336 30344 14370
rect 30378 14336 30434 14370
rect 30468 14336 30524 14370
rect 30558 14336 30617 14370
rect 29923 14332 30617 14336
rect 29923 14298 29996 14332
rect 30030 14298 30096 14332
rect 30130 14298 30196 14332
rect 30230 14298 30296 14332
rect 30330 14298 30396 14332
rect 30430 14298 30496 14332
rect 30530 14298 30617 14332
rect 29923 14280 30617 14298
rect 29923 14246 29984 14280
rect 30018 14246 30074 14280
rect 30108 14246 30164 14280
rect 30198 14246 30254 14280
rect 30288 14246 30344 14280
rect 30378 14246 30434 14280
rect 30468 14246 30524 14280
rect 30558 14246 30617 14280
rect 29923 14232 30617 14246
rect 29923 14198 29996 14232
rect 30030 14198 30096 14232
rect 30130 14198 30196 14232
rect 30230 14198 30296 14232
rect 30330 14198 30396 14232
rect 30430 14198 30496 14232
rect 30530 14198 30617 14232
rect 29923 14190 30617 14198
rect 29923 14156 29984 14190
rect 30018 14156 30074 14190
rect 30108 14156 30164 14190
rect 30198 14156 30254 14190
rect 30288 14156 30344 14190
rect 30378 14156 30434 14190
rect 30468 14156 30524 14190
rect 30558 14156 30617 14190
rect 29923 14132 30617 14156
rect 29923 14100 29996 14132
rect 30030 14100 30096 14132
rect 30130 14100 30196 14132
rect 30230 14100 30296 14132
rect 29923 14066 29984 14100
rect 30030 14098 30074 14100
rect 30130 14098 30164 14100
rect 30230 14098 30254 14100
rect 30018 14066 30074 14098
rect 30108 14066 30164 14098
rect 30198 14066 30254 14098
rect 30288 14098 30296 14100
rect 30330 14100 30396 14132
rect 30330 14098 30344 14100
rect 30288 14066 30344 14098
rect 30378 14098 30396 14100
rect 30430 14100 30496 14132
rect 30530 14100 30617 14132
rect 30430 14098 30434 14100
rect 30378 14066 30434 14098
rect 30468 14098 30496 14100
rect 30468 14066 30524 14098
rect 30558 14066 30617 14100
rect 29923 14032 30617 14066
rect 29923 14010 29996 14032
rect 30030 14010 30096 14032
rect 30130 14010 30196 14032
rect 30230 14010 30296 14032
rect 29923 13976 29984 14010
rect 30030 13998 30074 14010
rect 30130 13998 30164 14010
rect 30230 13998 30254 14010
rect 30018 13976 30074 13998
rect 30108 13976 30164 13998
rect 30198 13976 30254 13998
rect 30288 13998 30296 14010
rect 30330 14010 30396 14032
rect 30330 13998 30344 14010
rect 30288 13976 30344 13998
rect 30378 13998 30396 14010
rect 30430 14010 30496 14032
rect 30530 14010 30617 14032
rect 30430 13998 30434 14010
rect 30378 13976 30434 13998
rect 30468 13998 30496 14010
rect 30468 13976 30524 13998
rect 30558 13976 30617 14010
rect 29923 13932 30617 13976
rect 29923 13920 29996 13932
rect 30030 13920 30096 13932
rect 30130 13920 30196 13932
rect 30230 13920 30296 13932
rect 29923 13886 29984 13920
rect 30030 13898 30074 13920
rect 30130 13898 30164 13920
rect 30230 13898 30254 13920
rect 30018 13886 30074 13898
rect 30108 13886 30164 13898
rect 30198 13886 30254 13898
rect 30288 13898 30296 13920
rect 30330 13920 30396 13932
rect 30330 13898 30344 13920
rect 30288 13886 30344 13898
rect 30378 13898 30396 13920
rect 30430 13920 30496 13932
rect 30530 13920 30617 13932
rect 30430 13898 30434 13920
rect 30378 13886 30434 13898
rect 30468 13898 30496 13920
rect 30468 13886 30524 13898
rect 30558 13886 30617 13920
rect 29923 13825 30617 13886
rect 30679 14468 30751 14524
rect 30679 14434 30698 14468
rect 30732 14434 30751 14468
rect 30679 14378 30751 14434
rect 30679 14344 30698 14378
rect 30732 14344 30751 14378
rect 30679 14288 30751 14344
rect 30679 14254 30698 14288
rect 30732 14254 30751 14288
rect 30679 14198 30751 14254
rect 30679 14164 30698 14198
rect 30732 14164 30751 14198
rect 30679 14108 30751 14164
rect 30679 14074 30698 14108
rect 30732 14074 30751 14108
rect 30679 14018 30751 14074
rect 30679 13984 30698 14018
rect 30732 13984 30751 14018
rect 30679 13928 30751 13984
rect 30679 13894 30698 13928
rect 30732 13894 30751 13928
rect 30679 13838 30751 13894
rect 29789 13763 29861 13823
rect 30679 13804 30698 13838
rect 30732 13804 30751 13838
rect 30679 13763 30751 13804
rect 29789 13744 30751 13763
rect 29789 13710 29886 13744
rect 29920 13710 29976 13744
rect 30010 13710 30066 13744
rect 30100 13710 30156 13744
rect 30190 13710 30246 13744
rect 30280 13710 30336 13744
rect 30370 13710 30426 13744
rect 30460 13710 30516 13744
rect 30550 13710 30606 13744
rect 30640 13710 30751 13744
rect 29789 13691 30751 13710
rect 30815 14634 30847 14668
rect 30881 14634 31000 14668
rect 31034 14634 31065 14668
rect 32155 14668 32405 14717
rect 30815 14578 31065 14634
rect 30815 14544 30847 14578
rect 30881 14544 31000 14578
rect 31034 14544 31065 14578
rect 30815 14488 31065 14544
rect 30815 14454 30847 14488
rect 30881 14454 31000 14488
rect 31034 14454 31065 14488
rect 30815 14398 31065 14454
rect 30815 14364 30847 14398
rect 30881 14364 31000 14398
rect 31034 14364 31065 14398
rect 30815 14308 31065 14364
rect 30815 14274 30847 14308
rect 30881 14274 31000 14308
rect 31034 14274 31065 14308
rect 30815 14218 31065 14274
rect 30815 14184 30847 14218
rect 30881 14184 31000 14218
rect 31034 14184 31065 14218
rect 30815 14128 31065 14184
rect 30815 14094 30847 14128
rect 30881 14094 31000 14128
rect 31034 14094 31065 14128
rect 30815 14038 31065 14094
rect 30815 14004 30847 14038
rect 30881 14004 31000 14038
rect 31034 14004 31065 14038
rect 30815 13948 31065 14004
rect 30815 13914 30847 13948
rect 30881 13914 31000 13948
rect 31034 13914 31065 13948
rect 30815 13858 31065 13914
rect 30815 13824 30847 13858
rect 30881 13824 31000 13858
rect 31034 13824 31065 13858
rect 30815 13768 31065 13824
rect 30815 13734 30847 13768
rect 30881 13734 31000 13768
rect 31034 13734 31065 13768
rect 29475 13644 29507 13678
rect 29541 13644 29660 13678
rect 29694 13644 29725 13678
rect 29475 13627 29725 13644
rect 30815 13678 31065 13734
rect 31129 14636 32091 14653
rect 31129 14602 31150 14636
rect 31184 14602 31240 14636
rect 31274 14634 31330 14636
rect 31364 14634 31420 14636
rect 31454 14634 31510 14636
rect 31544 14634 31600 14636
rect 31634 14634 31690 14636
rect 31724 14634 31780 14636
rect 31814 14634 31870 14636
rect 31904 14634 31960 14636
rect 31994 14634 32050 14636
rect 31294 14602 31330 14634
rect 31384 14602 31420 14634
rect 31474 14602 31510 14634
rect 31564 14602 31600 14634
rect 31654 14602 31690 14634
rect 31744 14602 31780 14634
rect 31834 14602 31870 14634
rect 31924 14602 31960 14634
rect 32014 14602 32050 14634
rect 32084 14602 32091 14636
rect 31129 14600 31260 14602
rect 31294 14600 31350 14602
rect 31384 14600 31440 14602
rect 31474 14600 31530 14602
rect 31564 14600 31620 14602
rect 31654 14600 31710 14602
rect 31744 14600 31800 14602
rect 31834 14600 31890 14602
rect 31924 14600 31980 14602
rect 32014 14600 32091 14602
rect 31129 14581 32091 14600
rect 31129 14577 31201 14581
rect 31129 14543 31148 14577
rect 31182 14543 31201 14577
rect 31129 14487 31201 14543
rect 32019 14558 32091 14581
rect 32019 14524 32038 14558
rect 32072 14524 32091 14558
rect 31129 14453 31148 14487
rect 31182 14453 31201 14487
rect 31129 14397 31201 14453
rect 31129 14363 31148 14397
rect 31182 14363 31201 14397
rect 31129 14307 31201 14363
rect 31129 14273 31148 14307
rect 31182 14273 31201 14307
rect 31129 14217 31201 14273
rect 31129 14183 31148 14217
rect 31182 14183 31201 14217
rect 31129 14127 31201 14183
rect 31129 14093 31148 14127
rect 31182 14093 31201 14127
rect 31129 14037 31201 14093
rect 31129 14003 31148 14037
rect 31182 14003 31201 14037
rect 31129 13947 31201 14003
rect 31129 13913 31148 13947
rect 31182 13913 31201 13947
rect 31129 13857 31201 13913
rect 31129 13823 31148 13857
rect 31182 13823 31201 13857
rect 31263 14460 31957 14519
rect 31263 14426 31324 14460
rect 31358 14432 31414 14460
rect 31448 14432 31504 14460
rect 31538 14432 31594 14460
rect 31370 14426 31414 14432
rect 31470 14426 31504 14432
rect 31570 14426 31594 14432
rect 31628 14432 31684 14460
rect 31628 14426 31636 14432
rect 31263 14398 31336 14426
rect 31370 14398 31436 14426
rect 31470 14398 31536 14426
rect 31570 14398 31636 14426
rect 31670 14426 31684 14432
rect 31718 14432 31774 14460
rect 31718 14426 31736 14432
rect 31670 14398 31736 14426
rect 31770 14426 31774 14432
rect 31808 14432 31864 14460
rect 31808 14426 31836 14432
rect 31898 14426 31957 14460
rect 31770 14398 31836 14426
rect 31870 14398 31957 14426
rect 31263 14370 31957 14398
rect 31263 14336 31324 14370
rect 31358 14336 31414 14370
rect 31448 14336 31504 14370
rect 31538 14336 31594 14370
rect 31628 14336 31684 14370
rect 31718 14336 31774 14370
rect 31808 14336 31864 14370
rect 31898 14336 31957 14370
rect 31263 14332 31957 14336
rect 31263 14298 31336 14332
rect 31370 14298 31436 14332
rect 31470 14298 31536 14332
rect 31570 14298 31636 14332
rect 31670 14298 31736 14332
rect 31770 14298 31836 14332
rect 31870 14298 31957 14332
rect 31263 14280 31957 14298
rect 31263 14246 31324 14280
rect 31358 14246 31414 14280
rect 31448 14246 31504 14280
rect 31538 14246 31594 14280
rect 31628 14246 31684 14280
rect 31718 14246 31774 14280
rect 31808 14246 31864 14280
rect 31898 14246 31957 14280
rect 31263 14232 31957 14246
rect 31263 14198 31336 14232
rect 31370 14198 31436 14232
rect 31470 14198 31536 14232
rect 31570 14198 31636 14232
rect 31670 14198 31736 14232
rect 31770 14198 31836 14232
rect 31870 14198 31957 14232
rect 31263 14190 31957 14198
rect 31263 14156 31324 14190
rect 31358 14156 31414 14190
rect 31448 14156 31504 14190
rect 31538 14156 31594 14190
rect 31628 14156 31684 14190
rect 31718 14156 31774 14190
rect 31808 14156 31864 14190
rect 31898 14156 31957 14190
rect 31263 14132 31957 14156
rect 31263 14100 31336 14132
rect 31370 14100 31436 14132
rect 31470 14100 31536 14132
rect 31570 14100 31636 14132
rect 31263 14066 31324 14100
rect 31370 14098 31414 14100
rect 31470 14098 31504 14100
rect 31570 14098 31594 14100
rect 31358 14066 31414 14098
rect 31448 14066 31504 14098
rect 31538 14066 31594 14098
rect 31628 14098 31636 14100
rect 31670 14100 31736 14132
rect 31670 14098 31684 14100
rect 31628 14066 31684 14098
rect 31718 14098 31736 14100
rect 31770 14100 31836 14132
rect 31870 14100 31957 14132
rect 31770 14098 31774 14100
rect 31718 14066 31774 14098
rect 31808 14098 31836 14100
rect 31808 14066 31864 14098
rect 31898 14066 31957 14100
rect 31263 14032 31957 14066
rect 31263 14010 31336 14032
rect 31370 14010 31436 14032
rect 31470 14010 31536 14032
rect 31570 14010 31636 14032
rect 31263 13976 31324 14010
rect 31370 13998 31414 14010
rect 31470 13998 31504 14010
rect 31570 13998 31594 14010
rect 31358 13976 31414 13998
rect 31448 13976 31504 13998
rect 31538 13976 31594 13998
rect 31628 13998 31636 14010
rect 31670 14010 31736 14032
rect 31670 13998 31684 14010
rect 31628 13976 31684 13998
rect 31718 13998 31736 14010
rect 31770 14010 31836 14032
rect 31870 14010 31957 14032
rect 31770 13998 31774 14010
rect 31718 13976 31774 13998
rect 31808 13998 31836 14010
rect 31808 13976 31864 13998
rect 31898 13976 31957 14010
rect 31263 13932 31957 13976
rect 31263 13920 31336 13932
rect 31370 13920 31436 13932
rect 31470 13920 31536 13932
rect 31570 13920 31636 13932
rect 31263 13886 31324 13920
rect 31370 13898 31414 13920
rect 31470 13898 31504 13920
rect 31570 13898 31594 13920
rect 31358 13886 31414 13898
rect 31448 13886 31504 13898
rect 31538 13886 31594 13898
rect 31628 13898 31636 13920
rect 31670 13920 31736 13932
rect 31670 13898 31684 13920
rect 31628 13886 31684 13898
rect 31718 13898 31736 13920
rect 31770 13920 31836 13932
rect 31870 13920 31957 13932
rect 31770 13898 31774 13920
rect 31718 13886 31774 13898
rect 31808 13898 31836 13920
rect 31808 13886 31864 13898
rect 31898 13886 31957 13920
rect 31263 13825 31957 13886
rect 32019 14468 32091 14524
rect 32019 14434 32038 14468
rect 32072 14434 32091 14468
rect 32019 14378 32091 14434
rect 32019 14344 32038 14378
rect 32072 14344 32091 14378
rect 32019 14288 32091 14344
rect 32019 14254 32038 14288
rect 32072 14254 32091 14288
rect 32019 14198 32091 14254
rect 32019 14164 32038 14198
rect 32072 14164 32091 14198
rect 32019 14108 32091 14164
rect 32019 14074 32038 14108
rect 32072 14074 32091 14108
rect 32019 14018 32091 14074
rect 32019 13984 32038 14018
rect 32072 13984 32091 14018
rect 32019 13928 32091 13984
rect 32019 13894 32038 13928
rect 32072 13894 32091 13928
rect 32019 13838 32091 13894
rect 31129 13763 31201 13823
rect 32019 13804 32038 13838
rect 32072 13804 32091 13838
rect 32019 13763 32091 13804
rect 31129 13744 32091 13763
rect 31129 13710 31226 13744
rect 31260 13710 31316 13744
rect 31350 13710 31406 13744
rect 31440 13710 31496 13744
rect 31530 13710 31586 13744
rect 31620 13710 31676 13744
rect 31710 13710 31766 13744
rect 31800 13710 31856 13744
rect 31890 13710 31946 13744
rect 31980 13710 32091 13744
rect 31129 13691 32091 13710
rect 32155 14634 32187 14668
rect 32221 14634 32340 14668
rect 32374 14634 32405 14668
rect 33495 14668 33745 14717
rect 32155 14578 32405 14634
rect 32155 14544 32187 14578
rect 32221 14544 32340 14578
rect 32374 14544 32405 14578
rect 32155 14488 32405 14544
rect 32155 14454 32187 14488
rect 32221 14454 32340 14488
rect 32374 14454 32405 14488
rect 32155 14398 32405 14454
rect 32155 14364 32187 14398
rect 32221 14364 32340 14398
rect 32374 14364 32405 14398
rect 32155 14308 32405 14364
rect 32155 14274 32187 14308
rect 32221 14274 32340 14308
rect 32374 14274 32405 14308
rect 32155 14218 32405 14274
rect 32155 14184 32187 14218
rect 32221 14184 32340 14218
rect 32374 14184 32405 14218
rect 32155 14128 32405 14184
rect 32155 14094 32187 14128
rect 32221 14094 32340 14128
rect 32374 14094 32405 14128
rect 32155 14038 32405 14094
rect 32155 14004 32187 14038
rect 32221 14004 32340 14038
rect 32374 14004 32405 14038
rect 32155 13948 32405 14004
rect 32155 13914 32187 13948
rect 32221 13914 32340 13948
rect 32374 13914 32405 13948
rect 32155 13858 32405 13914
rect 32155 13824 32187 13858
rect 32221 13824 32340 13858
rect 32374 13824 32405 13858
rect 32155 13768 32405 13824
rect 32155 13734 32187 13768
rect 32221 13734 32340 13768
rect 32374 13734 32405 13768
rect 30815 13644 30847 13678
rect 30881 13644 31000 13678
rect 31034 13644 31065 13678
rect 30815 13627 31065 13644
rect 32155 13678 32405 13734
rect 32469 14636 33431 14653
rect 32469 14602 32490 14636
rect 32524 14602 32580 14636
rect 32614 14634 32670 14636
rect 32704 14634 32760 14636
rect 32794 14634 32850 14636
rect 32884 14634 32940 14636
rect 32974 14634 33030 14636
rect 33064 14634 33120 14636
rect 33154 14634 33210 14636
rect 33244 14634 33300 14636
rect 33334 14634 33390 14636
rect 32634 14602 32670 14634
rect 32724 14602 32760 14634
rect 32814 14602 32850 14634
rect 32904 14602 32940 14634
rect 32994 14602 33030 14634
rect 33084 14602 33120 14634
rect 33174 14602 33210 14634
rect 33264 14602 33300 14634
rect 33354 14602 33390 14634
rect 33424 14602 33431 14636
rect 32469 14600 32600 14602
rect 32634 14600 32690 14602
rect 32724 14600 32780 14602
rect 32814 14600 32870 14602
rect 32904 14600 32960 14602
rect 32994 14600 33050 14602
rect 33084 14600 33140 14602
rect 33174 14600 33230 14602
rect 33264 14600 33320 14602
rect 33354 14600 33431 14602
rect 32469 14581 33431 14600
rect 32469 14577 32541 14581
rect 32469 14543 32488 14577
rect 32522 14543 32541 14577
rect 32469 14487 32541 14543
rect 33359 14558 33431 14581
rect 33359 14524 33378 14558
rect 33412 14524 33431 14558
rect 32469 14453 32488 14487
rect 32522 14453 32541 14487
rect 32469 14397 32541 14453
rect 32469 14363 32488 14397
rect 32522 14363 32541 14397
rect 32469 14307 32541 14363
rect 32469 14273 32488 14307
rect 32522 14273 32541 14307
rect 32469 14217 32541 14273
rect 32469 14183 32488 14217
rect 32522 14183 32541 14217
rect 32469 14127 32541 14183
rect 32469 14093 32488 14127
rect 32522 14093 32541 14127
rect 32469 14037 32541 14093
rect 32469 14003 32488 14037
rect 32522 14003 32541 14037
rect 32469 13947 32541 14003
rect 32469 13913 32488 13947
rect 32522 13913 32541 13947
rect 32469 13857 32541 13913
rect 32469 13823 32488 13857
rect 32522 13823 32541 13857
rect 32603 14460 33297 14519
rect 32603 14426 32664 14460
rect 32698 14432 32754 14460
rect 32788 14432 32844 14460
rect 32878 14432 32934 14460
rect 32710 14426 32754 14432
rect 32810 14426 32844 14432
rect 32910 14426 32934 14432
rect 32968 14432 33024 14460
rect 32968 14426 32976 14432
rect 32603 14398 32676 14426
rect 32710 14398 32776 14426
rect 32810 14398 32876 14426
rect 32910 14398 32976 14426
rect 33010 14426 33024 14432
rect 33058 14432 33114 14460
rect 33058 14426 33076 14432
rect 33010 14398 33076 14426
rect 33110 14426 33114 14432
rect 33148 14432 33204 14460
rect 33148 14426 33176 14432
rect 33238 14426 33297 14460
rect 33110 14398 33176 14426
rect 33210 14398 33297 14426
rect 32603 14370 33297 14398
rect 32603 14336 32664 14370
rect 32698 14336 32754 14370
rect 32788 14336 32844 14370
rect 32878 14336 32934 14370
rect 32968 14336 33024 14370
rect 33058 14336 33114 14370
rect 33148 14336 33204 14370
rect 33238 14336 33297 14370
rect 32603 14332 33297 14336
rect 32603 14298 32676 14332
rect 32710 14298 32776 14332
rect 32810 14298 32876 14332
rect 32910 14298 32976 14332
rect 33010 14298 33076 14332
rect 33110 14298 33176 14332
rect 33210 14298 33297 14332
rect 32603 14280 33297 14298
rect 32603 14246 32664 14280
rect 32698 14246 32754 14280
rect 32788 14246 32844 14280
rect 32878 14246 32934 14280
rect 32968 14246 33024 14280
rect 33058 14246 33114 14280
rect 33148 14246 33204 14280
rect 33238 14246 33297 14280
rect 32603 14232 33297 14246
rect 32603 14198 32676 14232
rect 32710 14198 32776 14232
rect 32810 14198 32876 14232
rect 32910 14198 32976 14232
rect 33010 14198 33076 14232
rect 33110 14198 33176 14232
rect 33210 14198 33297 14232
rect 32603 14190 33297 14198
rect 32603 14156 32664 14190
rect 32698 14156 32754 14190
rect 32788 14156 32844 14190
rect 32878 14156 32934 14190
rect 32968 14156 33024 14190
rect 33058 14156 33114 14190
rect 33148 14156 33204 14190
rect 33238 14156 33297 14190
rect 32603 14132 33297 14156
rect 32603 14100 32676 14132
rect 32710 14100 32776 14132
rect 32810 14100 32876 14132
rect 32910 14100 32976 14132
rect 32603 14066 32664 14100
rect 32710 14098 32754 14100
rect 32810 14098 32844 14100
rect 32910 14098 32934 14100
rect 32698 14066 32754 14098
rect 32788 14066 32844 14098
rect 32878 14066 32934 14098
rect 32968 14098 32976 14100
rect 33010 14100 33076 14132
rect 33010 14098 33024 14100
rect 32968 14066 33024 14098
rect 33058 14098 33076 14100
rect 33110 14100 33176 14132
rect 33210 14100 33297 14132
rect 33110 14098 33114 14100
rect 33058 14066 33114 14098
rect 33148 14098 33176 14100
rect 33148 14066 33204 14098
rect 33238 14066 33297 14100
rect 32603 14032 33297 14066
rect 32603 14010 32676 14032
rect 32710 14010 32776 14032
rect 32810 14010 32876 14032
rect 32910 14010 32976 14032
rect 32603 13976 32664 14010
rect 32710 13998 32754 14010
rect 32810 13998 32844 14010
rect 32910 13998 32934 14010
rect 32698 13976 32754 13998
rect 32788 13976 32844 13998
rect 32878 13976 32934 13998
rect 32968 13998 32976 14010
rect 33010 14010 33076 14032
rect 33010 13998 33024 14010
rect 32968 13976 33024 13998
rect 33058 13998 33076 14010
rect 33110 14010 33176 14032
rect 33210 14010 33297 14032
rect 33110 13998 33114 14010
rect 33058 13976 33114 13998
rect 33148 13998 33176 14010
rect 33148 13976 33204 13998
rect 33238 13976 33297 14010
rect 32603 13932 33297 13976
rect 32603 13920 32676 13932
rect 32710 13920 32776 13932
rect 32810 13920 32876 13932
rect 32910 13920 32976 13932
rect 32603 13886 32664 13920
rect 32710 13898 32754 13920
rect 32810 13898 32844 13920
rect 32910 13898 32934 13920
rect 32698 13886 32754 13898
rect 32788 13886 32844 13898
rect 32878 13886 32934 13898
rect 32968 13898 32976 13920
rect 33010 13920 33076 13932
rect 33010 13898 33024 13920
rect 32968 13886 33024 13898
rect 33058 13898 33076 13920
rect 33110 13920 33176 13932
rect 33210 13920 33297 13932
rect 33110 13898 33114 13920
rect 33058 13886 33114 13898
rect 33148 13898 33176 13920
rect 33148 13886 33204 13898
rect 33238 13886 33297 13920
rect 32603 13825 33297 13886
rect 33359 14468 33431 14524
rect 33359 14434 33378 14468
rect 33412 14434 33431 14468
rect 33359 14378 33431 14434
rect 33359 14344 33378 14378
rect 33412 14344 33431 14378
rect 33359 14288 33431 14344
rect 33359 14254 33378 14288
rect 33412 14254 33431 14288
rect 33359 14198 33431 14254
rect 33359 14164 33378 14198
rect 33412 14164 33431 14198
rect 33359 14108 33431 14164
rect 33359 14074 33378 14108
rect 33412 14074 33431 14108
rect 33359 14018 33431 14074
rect 33359 13984 33378 14018
rect 33412 13984 33431 14018
rect 33359 13928 33431 13984
rect 33359 13894 33378 13928
rect 33412 13894 33431 13928
rect 33359 13838 33431 13894
rect 32469 13763 32541 13823
rect 33359 13804 33378 13838
rect 33412 13804 33431 13838
rect 33359 13763 33431 13804
rect 32469 13744 33431 13763
rect 32469 13710 32566 13744
rect 32600 13710 32656 13744
rect 32690 13710 32746 13744
rect 32780 13710 32836 13744
rect 32870 13710 32926 13744
rect 32960 13710 33016 13744
rect 33050 13710 33106 13744
rect 33140 13710 33196 13744
rect 33230 13710 33286 13744
rect 33320 13710 33431 13744
rect 32469 13691 33431 13710
rect 33495 14634 33527 14668
rect 33561 14634 33680 14668
rect 33714 14634 33745 14668
rect 34835 14668 35085 14717
rect 33495 14578 33745 14634
rect 33495 14544 33527 14578
rect 33561 14544 33680 14578
rect 33714 14544 33745 14578
rect 33495 14488 33745 14544
rect 33495 14454 33527 14488
rect 33561 14454 33680 14488
rect 33714 14454 33745 14488
rect 33495 14398 33745 14454
rect 33495 14364 33527 14398
rect 33561 14364 33680 14398
rect 33714 14364 33745 14398
rect 33495 14308 33745 14364
rect 33495 14274 33527 14308
rect 33561 14274 33680 14308
rect 33714 14274 33745 14308
rect 33495 14218 33745 14274
rect 33495 14184 33527 14218
rect 33561 14184 33680 14218
rect 33714 14184 33745 14218
rect 33495 14128 33745 14184
rect 33495 14094 33527 14128
rect 33561 14094 33680 14128
rect 33714 14094 33745 14128
rect 33495 14038 33745 14094
rect 33495 14004 33527 14038
rect 33561 14004 33680 14038
rect 33714 14004 33745 14038
rect 33495 13948 33745 14004
rect 33495 13914 33527 13948
rect 33561 13914 33680 13948
rect 33714 13914 33745 13948
rect 33495 13858 33745 13914
rect 33495 13824 33527 13858
rect 33561 13824 33680 13858
rect 33714 13824 33745 13858
rect 33495 13768 33745 13824
rect 33495 13734 33527 13768
rect 33561 13734 33680 13768
rect 33714 13734 33745 13768
rect 32155 13644 32187 13678
rect 32221 13644 32340 13678
rect 32374 13644 32405 13678
rect 32155 13627 32405 13644
rect 33495 13678 33745 13734
rect 33809 14636 34771 14653
rect 33809 14602 33830 14636
rect 33864 14602 33920 14636
rect 33954 14634 34010 14636
rect 34044 14634 34100 14636
rect 34134 14634 34190 14636
rect 34224 14634 34280 14636
rect 34314 14634 34370 14636
rect 34404 14634 34460 14636
rect 34494 14634 34550 14636
rect 34584 14634 34640 14636
rect 34674 14634 34730 14636
rect 33974 14602 34010 14634
rect 34064 14602 34100 14634
rect 34154 14602 34190 14634
rect 34244 14602 34280 14634
rect 34334 14602 34370 14634
rect 34424 14602 34460 14634
rect 34514 14602 34550 14634
rect 34604 14602 34640 14634
rect 34694 14602 34730 14634
rect 34764 14602 34771 14636
rect 33809 14600 33940 14602
rect 33974 14600 34030 14602
rect 34064 14600 34120 14602
rect 34154 14600 34210 14602
rect 34244 14600 34300 14602
rect 34334 14600 34390 14602
rect 34424 14600 34480 14602
rect 34514 14600 34570 14602
rect 34604 14600 34660 14602
rect 34694 14600 34771 14602
rect 33809 14581 34771 14600
rect 33809 14577 33881 14581
rect 33809 14543 33828 14577
rect 33862 14543 33881 14577
rect 33809 14487 33881 14543
rect 34699 14558 34771 14581
rect 34699 14524 34718 14558
rect 34752 14524 34771 14558
rect 33809 14453 33828 14487
rect 33862 14453 33881 14487
rect 33809 14397 33881 14453
rect 33809 14363 33828 14397
rect 33862 14363 33881 14397
rect 33809 14307 33881 14363
rect 33809 14273 33828 14307
rect 33862 14273 33881 14307
rect 33809 14217 33881 14273
rect 33809 14183 33828 14217
rect 33862 14183 33881 14217
rect 33809 14127 33881 14183
rect 33809 14093 33828 14127
rect 33862 14093 33881 14127
rect 33809 14037 33881 14093
rect 33809 14003 33828 14037
rect 33862 14003 33881 14037
rect 33809 13947 33881 14003
rect 33809 13913 33828 13947
rect 33862 13913 33881 13947
rect 33809 13857 33881 13913
rect 33809 13823 33828 13857
rect 33862 13823 33881 13857
rect 33943 14460 34637 14519
rect 33943 14426 34004 14460
rect 34038 14432 34094 14460
rect 34128 14432 34184 14460
rect 34218 14432 34274 14460
rect 34050 14426 34094 14432
rect 34150 14426 34184 14432
rect 34250 14426 34274 14432
rect 34308 14432 34364 14460
rect 34308 14426 34316 14432
rect 33943 14398 34016 14426
rect 34050 14398 34116 14426
rect 34150 14398 34216 14426
rect 34250 14398 34316 14426
rect 34350 14426 34364 14432
rect 34398 14432 34454 14460
rect 34398 14426 34416 14432
rect 34350 14398 34416 14426
rect 34450 14426 34454 14432
rect 34488 14432 34544 14460
rect 34488 14426 34516 14432
rect 34578 14426 34637 14460
rect 34450 14398 34516 14426
rect 34550 14398 34637 14426
rect 33943 14370 34637 14398
rect 33943 14336 34004 14370
rect 34038 14336 34094 14370
rect 34128 14336 34184 14370
rect 34218 14336 34274 14370
rect 34308 14336 34364 14370
rect 34398 14336 34454 14370
rect 34488 14336 34544 14370
rect 34578 14336 34637 14370
rect 33943 14332 34637 14336
rect 33943 14298 34016 14332
rect 34050 14298 34116 14332
rect 34150 14298 34216 14332
rect 34250 14298 34316 14332
rect 34350 14298 34416 14332
rect 34450 14298 34516 14332
rect 34550 14298 34637 14332
rect 33943 14280 34637 14298
rect 33943 14246 34004 14280
rect 34038 14246 34094 14280
rect 34128 14246 34184 14280
rect 34218 14246 34274 14280
rect 34308 14246 34364 14280
rect 34398 14246 34454 14280
rect 34488 14246 34544 14280
rect 34578 14246 34637 14280
rect 33943 14232 34637 14246
rect 33943 14198 34016 14232
rect 34050 14198 34116 14232
rect 34150 14198 34216 14232
rect 34250 14198 34316 14232
rect 34350 14198 34416 14232
rect 34450 14198 34516 14232
rect 34550 14198 34637 14232
rect 33943 14190 34637 14198
rect 33943 14156 34004 14190
rect 34038 14156 34094 14190
rect 34128 14156 34184 14190
rect 34218 14156 34274 14190
rect 34308 14156 34364 14190
rect 34398 14156 34454 14190
rect 34488 14156 34544 14190
rect 34578 14156 34637 14190
rect 33943 14132 34637 14156
rect 33943 14100 34016 14132
rect 34050 14100 34116 14132
rect 34150 14100 34216 14132
rect 34250 14100 34316 14132
rect 33943 14066 34004 14100
rect 34050 14098 34094 14100
rect 34150 14098 34184 14100
rect 34250 14098 34274 14100
rect 34038 14066 34094 14098
rect 34128 14066 34184 14098
rect 34218 14066 34274 14098
rect 34308 14098 34316 14100
rect 34350 14100 34416 14132
rect 34350 14098 34364 14100
rect 34308 14066 34364 14098
rect 34398 14098 34416 14100
rect 34450 14100 34516 14132
rect 34550 14100 34637 14132
rect 34450 14098 34454 14100
rect 34398 14066 34454 14098
rect 34488 14098 34516 14100
rect 34488 14066 34544 14098
rect 34578 14066 34637 14100
rect 33943 14032 34637 14066
rect 33943 14010 34016 14032
rect 34050 14010 34116 14032
rect 34150 14010 34216 14032
rect 34250 14010 34316 14032
rect 33943 13976 34004 14010
rect 34050 13998 34094 14010
rect 34150 13998 34184 14010
rect 34250 13998 34274 14010
rect 34038 13976 34094 13998
rect 34128 13976 34184 13998
rect 34218 13976 34274 13998
rect 34308 13998 34316 14010
rect 34350 14010 34416 14032
rect 34350 13998 34364 14010
rect 34308 13976 34364 13998
rect 34398 13998 34416 14010
rect 34450 14010 34516 14032
rect 34550 14010 34637 14032
rect 34450 13998 34454 14010
rect 34398 13976 34454 13998
rect 34488 13998 34516 14010
rect 34488 13976 34544 13998
rect 34578 13976 34637 14010
rect 33943 13932 34637 13976
rect 33943 13920 34016 13932
rect 34050 13920 34116 13932
rect 34150 13920 34216 13932
rect 34250 13920 34316 13932
rect 33943 13886 34004 13920
rect 34050 13898 34094 13920
rect 34150 13898 34184 13920
rect 34250 13898 34274 13920
rect 34038 13886 34094 13898
rect 34128 13886 34184 13898
rect 34218 13886 34274 13898
rect 34308 13898 34316 13920
rect 34350 13920 34416 13932
rect 34350 13898 34364 13920
rect 34308 13886 34364 13898
rect 34398 13898 34416 13920
rect 34450 13920 34516 13932
rect 34550 13920 34637 13932
rect 34450 13898 34454 13920
rect 34398 13886 34454 13898
rect 34488 13898 34516 13920
rect 34488 13886 34544 13898
rect 34578 13886 34637 13920
rect 33943 13825 34637 13886
rect 34699 14468 34771 14524
rect 34699 14434 34718 14468
rect 34752 14434 34771 14468
rect 34699 14378 34771 14434
rect 34699 14344 34718 14378
rect 34752 14344 34771 14378
rect 34699 14288 34771 14344
rect 34699 14254 34718 14288
rect 34752 14254 34771 14288
rect 34699 14198 34771 14254
rect 34699 14164 34718 14198
rect 34752 14164 34771 14198
rect 34699 14108 34771 14164
rect 34699 14074 34718 14108
rect 34752 14074 34771 14108
rect 34699 14018 34771 14074
rect 34699 13984 34718 14018
rect 34752 13984 34771 14018
rect 34699 13928 34771 13984
rect 34699 13894 34718 13928
rect 34752 13894 34771 13928
rect 34699 13838 34771 13894
rect 33809 13763 33881 13823
rect 34699 13804 34718 13838
rect 34752 13804 34771 13838
rect 34699 13763 34771 13804
rect 33809 13744 34771 13763
rect 33809 13710 33906 13744
rect 33940 13710 33996 13744
rect 34030 13710 34086 13744
rect 34120 13710 34176 13744
rect 34210 13710 34266 13744
rect 34300 13710 34356 13744
rect 34390 13710 34446 13744
rect 34480 13710 34536 13744
rect 34570 13710 34626 13744
rect 34660 13710 34771 13744
rect 33809 13691 34771 13710
rect 34835 14634 34867 14668
rect 34901 14634 35020 14668
rect 35054 14634 35085 14668
rect 36175 14668 36425 14717
rect 34835 14578 35085 14634
rect 34835 14544 34867 14578
rect 34901 14544 35020 14578
rect 35054 14544 35085 14578
rect 34835 14488 35085 14544
rect 34835 14454 34867 14488
rect 34901 14454 35020 14488
rect 35054 14454 35085 14488
rect 34835 14398 35085 14454
rect 34835 14364 34867 14398
rect 34901 14364 35020 14398
rect 35054 14364 35085 14398
rect 34835 14308 35085 14364
rect 34835 14274 34867 14308
rect 34901 14274 35020 14308
rect 35054 14274 35085 14308
rect 34835 14218 35085 14274
rect 34835 14184 34867 14218
rect 34901 14184 35020 14218
rect 35054 14184 35085 14218
rect 34835 14128 35085 14184
rect 34835 14094 34867 14128
rect 34901 14094 35020 14128
rect 35054 14094 35085 14128
rect 34835 14038 35085 14094
rect 34835 14004 34867 14038
rect 34901 14004 35020 14038
rect 35054 14004 35085 14038
rect 34835 13948 35085 14004
rect 34835 13914 34867 13948
rect 34901 13914 35020 13948
rect 35054 13914 35085 13948
rect 34835 13858 35085 13914
rect 34835 13824 34867 13858
rect 34901 13824 35020 13858
rect 35054 13824 35085 13858
rect 34835 13768 35085 13824
rect 34835 13734 34867 13768
rect 34901 13734 35020 13768
rect 35054 13734 35085 13768
rect 33495 13644 33527 13678
rect 33561 13644 33680 13678
rect 33714 13644 33745 13678
rect 33495 13627 33745 13644
rect 34835 13678 35085 13734
rect 35149 14636 36111 14653
rect 35149 14602 35170 14636
rect 35204 14602 35260 14636
rect 35294 14634 35350 14636
rect 35384 14634 35440 14636
rect 35474 14634 35530 14636
rect 35564 14634 35620 14636
rect 35654 14634 35710 14636
rect 35744 14634 35800 14636
rect 35834 14634 35890 14636
rect 35924 14634 35980 14636
rect 36014 14634 36070 14636
rect 35314 14602 35350 14634
rect 35404 14602 35440 14634
rect 35494 14602 35530 14634
rect 35584 14602 35620 14634
rect 35674 14602 35710 14634
rect 35764 14602 35800 14634
rect 35854 14602 35890 14634
rect 35944 14602 35980 14634
rect 36034 14602 36070 14634
rect 36104 14602 36111 14636
rect 35149 14600 35280 14602
rect 35314 14600 35370 14602
rect 35404 14600 35460 14602
rect 35494 14600 35550 14602
rect 35584 14600 35640 14602
rect 35674 14600 35730 14602
rect 35764 14600 35820 14602
rect 35854 14600 35910 14602
rect 35944 14600 36000 14602
rect 36034 14600 36111 14602
rect 35149 14581 36111 14600
rect 35149 14577 35221 14581
rect 35149 14543 35168 14577
rect 35202 14543 35221 14577
rect 35149 14487 35221 14543
rect 36039 14558 36111 14581
rect 36039 14524 36058 14558
rect 36092 14524 36111 14558
rect 35149 14453 35168 14487
rect 35202 14453 35221 14487
rect 35149 14397 35221 14453
rect 35149 14363 35168 14397
rect 35202 14363 35221 14397
rect 35149 14307 35221 14363
rect 35149 14273 35168 14307
rect 35202 14273 35221 14307
rect 35149 14217 35221 14273
rect 35149 14183 35168 14217
rect 35202 14183 35221 14217
rect 35149 14127 35221 14183
rect 35149 14093 35168 14127
rect 35202 14093 35221 14127
rect 35149 14037 35221 14093
rect 35149 14003 35168 14037
rect 35202 14003 35221 14037
rect 35149 13947 35221 14003
rect 35149 13913 35168 13947
rect 35202 13913 35221 13947
rect 35149 13857 35221 13913
rect 35149 13823 35168 13857
rect 35202 13823 35221 13857
rect 35283 14460 35977 14519
rect 35283 14426 35344 14460
rect 35378 14432 35434 14460
rect 35468 14432 35524 14460
rect 35558 14432 35614 14460
rect 35390 14426 35434 14432
rect 35490 14426 35524 14432
rect 35590 14426 35614 14432
rect 35648 14432 35704 14460
rect 35648 14426 35656 14432
rect 35283 14398 35356 14426
rect 35390 14398 35456 14426
rect 35490 14398 35556 14426
rect 35590 14398 35656 14426
rect 35690 14426 35704 14432
rect 35738 14432 35794 14460
rect 35738 14426 35756 14432
rect 35690 14398 35756 14426
rect 35790 14426 35794 14432
rect 35828 14432 35884 14460
rect 35828 14426 35856 14432
rect 35918 14426 35977 14460
rect 35790 14398 35856 14426
rect 35890 14398 35977 14426
rect 35283 14370 35977 14398
rect 35283 14336 35344 14370
rect 35378 14336 35434 14370
rect 35468 14336 35524 14370
rect 35558 14336 35614 14370
rect 35648 14336 35704 14370
rect 35738 14336 35794 14370
rect 35828 14336 35884 14370
rect 35918 14336 35977 14370
rect 35283 14332 35977 14336
rect 35283 14298 35356 14332
rect 35390 14298 35456 14332
rect 35490 14298 35556 14332
rect 35590 14298 35656 14332
rect 35690 14298 35756 14332
rect 35790 14298 35856 14332
rect 35890 14298 35977 14332
rect 35283 14280 35977 14298
rect 35283 14246 35344 14280
rect 35378 14246 35434 14280
rect 35468 14246 35524 14280
rect 35558 14246 35614 14280
rect 35648 14246 35704 14280
rect 35738 14246 35794 14280
rect 35828 14246 35884 14280
rect 35918 14246 35977 14280
rect 35283 14232 35977 14246
rect 35283 14198 35356 14232
rect 35390 14198 35456 14232
rect 35490 14198 35556 14232
rect 35590 14198 35656 14232
rect 35690 14198 35756 14232
rect 35790 14198 35856 14232
rect 35890 14198 35977 14232
rect 35283 14190 35977 14198
rect 35283 14156 35344 14190
rect 35378 14156 35434 14190
rect 35468 14156 35524 14190
rect 35558 14156 35614 14190
rect 35648 14156 35704 14190
rect 35738 14156 35794 14190
rect 35828 14156 35884 14190
rect 35918 14156 35977 14190
rect 35283 14132 35977 14156
rect 35283 14100 35356 14132
rect 35390 14100 35456 14132
rect 35490 14100 35556 14132
rect 35590 14100 35656 14132
rect 35283 14066 35344 14100
rect 35390 14098 35434 14100
rect 35490 14098 35524 14100
rect 35590 14098 35614 14100
rect 35378 14066 35434 14098
rect 35468 14066 35524 14098
rect 35558 14066 35614 14098
rect 35648 14098 35656 14100
rect 35690 14100 35756 14132
rect 35690 14098 35704 14100
rect 35648 14066 35704 14098
rect 35738 14098 35756 14100
rect 35790 14100 35856 14132
rect 35890 14100 35977 14132
rect 35790 14098 35794 14100
rect 35738 14066 35794 14098
rect 35828 14098 35856 14100
rect 35828 14066 35884 14098
rect 35918 14066 35977 14100
rect 35283 14032 35977 14066
rect 35283 14010 35356 14032
rect 35390 14010 35456 14032
rect 35490 14010 35556 14032
rect 35590 14010 35656 14032
rect 35283 13976 35344 14010
rect 35390 13998 35434 14010
rect 35490 13998 35524 14010
rect 35590 13998 35614 14010
rect 35378 13976 35434 13998
rect 35468 13976 35524 13998
rect 35558 13976 35614 13998
rect 35648 13998 35656 14010
rect 35690 14010 35756 14032
rect 35690 13998 35704 14010
rect 35648 13976 35704 13998
rect 35738 13998 35756 14010
rect 35790 14010 35856 14032
rect 35890 14010 35977 14032
rect 35790 13998 35794 14010
rect 35738 13976 35794 13998
rect 35828 13998 35856 14010
rect 35828 13976 35884 13998
rect 35918 13976 35977 14010
rect 35283 13932 35977 13976
rect 35283 13920 35356 13932
rect 35390 13920 35456 13932
rect 35490 13920 35556 13932
rect 35590 13920 35656 13932
rect 35283 13886 35344 13920
rect 35390 13898 35434 13920
rect 35490 13898 35524 13920
rect 35590 13898 35614 13920
rect 35378 13886 35434 13898
rect 35468 13886 35524 13898
rect 35558 13886 35614 13898
rect 35648 13898 35656 13920
rect 35690 13920 35756 13932
rect 35690 13898 35704 13920
rect 35648 13886 35704 13898
rect 35738 13898 35756 13920
rect 35790 13920 35856 13932
rect 35890 13920 35977 13932
rect 35790 13898 35794 13920
rect 35738 13886 35794 13898
rect 35828 13898 35856 13920
rect 35828 13886 35884 13898
rect 35918 13886 35977 13920
rect 35283 13825 35977 13886
rect 36039 14468 36111 14524
rect 36039 14434 36058 14468
rect 36092 14434 36111 14468
rect 36039 14378 36111 14434
rect 36039 14344 36058 14378
rect 36092 14344 36111 14378
rect 36039 14288 36111 14344
rect 36039 14254 36058 14288
rect 36092 14254 36111 14288
rect 36039 14198 36111 14254
rect 36039 14164 36058 14198
rect 36092 14164 36111 14198
rect 36039 14108 36111 14164
rect 36039 14074 36058 14108
rect 36092 14074 36111 14108
rect 36039 14018 36111 14074
rect 36039 13984 36058 14018
rect 36092 13984 36111 14018
rect 36039 13928 36111 13984
rect 36039 13894 36058 13928
rect 36092 13894 36111 13928
rect 36039 13838 36111 13894
rect 35149 13763 35221 13823
rect 36039 13804 36058 13838
rect 36092 13804 36111 13838
rect 36039 13763 36111 13804
rect 35149 13744 36111 13763
rect 35149 13710 35246 13744
rect 35280 13710 35336 13744
rect 35370 13710 35426 13744
rect 35460 13710 35516 13744
rect 35550 13710 35606 13744
rect 35640 13710 35696 13744
rect 35730 13710 35786 13744
rect 35820 13710 35876 13744
rect 35910 13710 35966 13744
rect 36000 13710 36111 13744
rect 35149 13691 36111 13710
rect 36175 14634 36207 14668
rect 36241 14634 36360 14668
rect 36394 14634 36425 14668
rect 37515 14668 37765 14717
rect 36175 14578 36425 14634
rect 36175 14544 36207 14578
rect 36241 14544 36360 14578
rect 36394 14544 36425 14578
rect 36175 14488 36425 14544
rect 36175 14454 36207 14488
rect 36241 14454 36360 14488
rect 36394 14454 36425 14488
rect 36175 14398 36425 14454
rect 36175 14364 36207 14398
rect 36241 14364 36360 14398
rect 36394 14364 36425 14398
rect 36175 14308 36425 14364
rect 36175 14274 36207 14308
rect 36241 14274 36360 14308
rect 36394 14274 36425 14308
rect 36175 14218 36425 14274
rect 36175 14184 36207 14218
rect 36241 14184 36360 14218
rect 36394 14184 36425 14218
rect 36175 14128 36425 14184
rect 36175 14094 36207 14128
rect 36241 14094 36360 14128
rect 36394 14094 36425 14128
rect 36175 14038 36425 14094
rect 36175 14004 36207 14038
rect 36241 14004 36360 14038
rect 36394 14004 36425 14038
rect 36175 13948 36425 14004
rect 36175 13914 36207 13948
rect 36241 13914 36360 13948
rect 36394 13914 36425 13948
rect 36175 13858 36425 13914
rect 36175 13824 36207 13858
rect 36241 13824 36360 13858
rect 36394 13824 36425 13858
rect 36175 13768 36425 13824
rect 36175 13734 36207 13768
rect 36241 13734 36360 13768
rect 36394 13734 36425 13768
rect 34835 13644 34867 13678
rect 34901 13644 35020 13678
rect 35054 13644 35085 13678
rect 34835 13627 35085 13644
rect 36175 13678 36425 13734
rect 36489 14636 37451 14653
rect 36489 14602 36510 14636
rect 36544 14602 36600 14636
rect 36634 14634 36690 14636
rect 36724 14634 36780 14636
rect 36814 14634 36870 14636
rect 36904 14634 36960 14636
rect 36994 14634 37050 14636
rect 37084 14634 37140 14636
rect 37174 14634 37230 14636
rect 37264 14634 37320 14636
rect 37354 14634 37410 14636
rect 36654 14602 36690 14634
rect 36744 14602 36780 14634
rect 36834 14602 36870 14634
rect 36924 14602 36960 14634
rect 37014 14602 37050 14634
rect 37104 14602 37140 14634
rect 37194 14602 37230 14634
rect 37284 14602 37320 14634
rect 37374 14602 37410 14634
rect 37444 14602 37451 14636
rect 36489 14600 36620 14602
rect 36654 14600 36710 14602
rect 36744 14600 36800 14602
rect 36834 14600 36890 14602
rect 36924 14600 36980 14602
rect 37014 14600 37070 14602
rect 37104 14600 37160 14602
rect 37194 14600 37250 14602
rect 37284 14600 37340 14602
rect 37374 14600 37451 14602
rect 36489 14581 37451 14600
rect 36489 14577 36561 14581
rect 36489 14543 36508 14577
rect 36542 14543 36561 14577
rect 36489 14487 36561 14543
rect 37379 14558 37451 14581
rect 37379 14524 37398 14558
rect 37432 14524 37451 14558
rect 36489 14453 36508 14487
rect 36542 14453 36561 14487
rect 36489 14397 36561 14453
rect 36489 14363 36508 14397
rect 36542 14363 36561 14397
rect 36489 14307 36561 14363
rect 36489 14273 36508 14307
rect 36542 14273 36561 14307
rect 36489 14217 36561 14273
rect 36489 14183 36508 14217
rect 36542 14183 36561 14217
rect 36489 14127 36561 14183
rect 36489 14093 36508 14127
rect 36542 14093 36561 14127
rect 36489 14037 36561 14093
rect 36489 14003 36508 14037
rect 36542 14003 36561 14037
rect 36489 13947 36561 14003
rect 36489 13913 36508 13947
rect 36542 13913 36561 13947
rect 36489 13857 36561 13913
rect 36489 13823 36508 13857
rect 36542 13823 36561 13857
rect 36623 14460 37317 14519
rect 36623 14426 36684 14460
rect 36718 14432 36774 14460
rect 36808 14432 36864 14460
rect 36898 14432 36954 14460
rect 36730 14426 36774 14432
rect 36830 14426 36864 14432
rect 36930 14426 36954 14432
rect 36988 14432 37044 14460
rect 36988 14426 36996 14432
rect 36623 14398 36696 14426
rect 36730 14398 36796 14426
rect 36830 14398 36896 14426
rect 36930 14398 36996 14426
rect 37030 14426 37044 14432
rect 37078 14432 37134 14460
rect 37078 14426 37096 14432
rect 37030 14398 37096 14426
rect 37130 14426 37134 14432
rect 37168 14432 37224 14460
rect 37168 14426 37196 14432
rect 37258 14426 37317 14460
rect 37130 14398 37196 14426
rect 37230 14398 37317 14426
rect 36623 14370 37317 14398
rect 36623 14336 36684 14370
rect 36718 14336 36774 14370
rect 36808 14336 36864 14370
rect 36898 14336 36954 14370
rect 36988 14336 37044 14370
rect 37078 14336 37134 14370
rect 37168 14336 37224 14370
rect 37258 14336 37317 14370
rect 36623 14332 37317 14336
rect 36623 14298 36696 14332
rect 36730 14298 36796 14332
rect 36830 14298 36896 14332
rect 36930 14298 36996 14332
rect 37030 14298 37096 14332
rect 37130 14298 37196 14332
rect 37230 14298 37317 14332
rect 36623 14280 37317 14298
rect 36623 14246 36684 14280
rect 36718 14246 36774 14280
rect 36808 14246 36864 14280
rect 36898 14246 36954 14280
rect 36988 14246 37044 14280
rect 37078 14246 37134 14280
rect 37168 14246 37224 14280
rect 37258 14246 37317 14280
rect 36623 14232 37317 14246
rect 36623 14198 36696 14232
rect 36730 14198 36796 14232
rect 36830 14198 36896 14232
rect 36930 14198 36996 14232
rect 37030 14198 37096 14232
rect 37130 14198 37196 14232
rect 37230 14198 37317 14232
rect 36623 14190 37317 14198
rect 36623 14156 36684 14190
rect 36718 14156 36774 14190
rect 36808 14156 36864 14190
rect 36898 14156 36954 14190
rect 36988 14156 37044 14190
rect 37078 14156 37134 14190
rect 37168 14156 37224 14190
rect 37258 14156 37317 14190
rect 36623 14132 37317 14156
rect 36623 14100 36696 14132
rect 36730 14100 36796 14132
rect 36830 14100 36896 14132
rect 36930 14100 36996 14132
rect 36623 14066 36684 14100
rect 36730 14098 36774 14100
rect 36830 14098 36864 14100
rect 36930 14098 36954 14100
rect 36718 14066 36774 14098
rect 36808 14066 36864 14098
rect 36898 14066 36954 14098
rect 36988 14098 36996 14100
rect 37030 14100 37096 14132
rect 37030 14098 37044 14100
rect 36988 14066 37044 14098
rect 37078 14098 37096 14100
rect 37130 14100 37196 14132
rect 37230 14100 37317 14132
rect 37130 14098 37134 14100
rect 37078 14066 37134 14098
rect 37168 14098 37196 14100
rect 37168 14066 37224 14098
rect 37258 14066 37317 14100
rect 36623 14032 37317 14066
rect 36623 14010 36696 14032
rect 36730 14010 36796 14032
rect 36830 14010 36896 14032
rect 36930 14010 36996 14032
rect 36623 13976 36684 14010
rect 36730 13998 36774 14010
rect 36830 13998 36864 14010
rect 36930 13998 36954 14010
rect 36718 13976 36774 13998
rect 36808 13976 36864 13998
rect 36898 13976 36954 13998
rect 36988 13998 36996 14010
rect 37030 14010 37096 14032
rect 37030 13998 37044 14010
rect 36988 13976 37044 13998
rect 37078 13998 37096 14010
rect 37130 14010 37196 14032
rect 37230 14010 37317 14032
rect 37130 13998 37134 14010
rect 37078 13976 37134 13998
rect 37168 13998 37196 14010
rect 37168 13976 37224 13998
rect 37258 13976 37317 14010
rect 36623 13932 37317 13976
rect 36623 13920 36696 13932
rect 36730 13920 36796 13932
rect 36830 13920 36896 13932
rect 36930 13920 36996 13932
rect 36623 13886 36684 13920
rect 36730 13898 36774 13920
rect 36830 13898 36864 13920
rect 36930 13898 36954 13920
rect 36718 13886 36774 13898
rect 36808 13886 36864 13898
rect 36898 13886 36954 13898
rect 36988 13898 36996 13920
rect 37030 13920 37096 13932
rect 37030 13898 37044 13920
rect 36988 13886 37044 13898
rect 37078 13898 37096 13920
rect 37130 13920 37196 13932
rect 37230 13920 37317 13932
rect 37130 13898 37134 13920
rect 37078 13886 37134 13898
rect 37168 13898 37196 13920
rect 37168 13886 37224 13898
rect 37258 13886 37317 13920
rect 36623 13825 37317 13886
rect 37379 14468 37451 14524
rect 37379 14434 37398 14468
rect 37432 14434 37451 14468
rect 37379 14378 37451 14434
rect 37379 14344 37398 14378
rect 37432 14344 37451 14378
rect 37379 14288 37451 14344
rect 37379 14254 37398 14288
rect 37432 14254 37451 14288
rect 37379 14198 37451 14254
rect 37379 14164 37398 14198
rect 37432 14164 37451 14198
rect 37379 14108 37451 14164
rect 37379 14074 37398 14108
rect 37432 14074 37451 14108
rect 37379 14018 37451 14074
rect 37379 13984 37398 14018
rect 37432 13984 37451 14018
rect 37379 13928 37451 13984
rect 37379 13894 37398 13928
rect 37432 13894 37451 13928
rect 37379 13838 37451 13894
rect 36489 13763 36561 13823
rect 37379 13804 37398 13838
rect 37432 13804 37451 13838
rect 37379 13763 37451 13804
rect 36489 13744 37451 13763
rect 36489 13710 36586 13744
rect 36620 13710 36676 13744
rect 36710 13710 36766 13744
rect 36800 13710 36856 13744
rect 36890 13710 36946 13744
rect 36980 13710 37036 13744
rect 37070 13710 37126 13744
rect 37160 13710 37216 13744
rect 37250 13710 37306 13744
rect 37340 13710 37451 13744
rect 36489 13691 37451 13710
rect 37515 14634 37547 14668
rect 37581 14634 37700 14668
rect 37734 14634 37765 14668
rect 38855 14668 38954 14717
rect 37515 14578 37765 14634
rect 37515 14544 37547 14578
rect 37581 14544 37700 14578
rect 37734 14544 37765 14578
rect 37515 14488 37765 14544
rect 37515 14454 37547 14488
rect 37581 14454 37700 14488
rect 37734 14454 37765 14488
rect 37515 14398 37765 14454
rect 37515 14364 37547 14398
rect 37581 14364 37700 14398
rect 37734 14364 37765 14398
rect 37515 14308 37765 14364
rect 37515 14274 37547 14308
rect 37581 14274 37700 14308
rect 37734 14274 37765 14308
rect 37515 14218 37765 14274
rect 37515 14184 37547 14218
rect 37581 14184 37700 14218
rect 37734 14184 37765 14218
rect 37515 14128 37765 14184
rect 37515 14094 37547 14128
rect 37581 14094 37700 14128
rect 37734 14094 37765 14128
rect 37515 14038 37765 14094
rect 37515 14004 37547 14038
rect 37581 14004 37700 14038
rect 37734 14004 37765 14038
rect 37515 13948 37765 14004
rect 37515 13914 37547 13948
rect 37581 13914 37700 13948
rect 37734 13914 37765 13948
rect 37515 13858 37765 13914
rect 37515 13824 37547 13858
rect 37581 13824 37700 13858
rect 37734 13824 37765 13858
rect 37515 13768 37765 13824
rect 37515 13734 37547 13768
rect 37581 13734 37700 13768
rect 37734 13734 37765 13768
rect 36175 13644 36207 13678
rect 36241 13644 36360 13678
rect 36394 13644 36425 13678
rect 36175 13627 36425 13644
rect 37515 13678 37765 13734
rect 37829 14636 38791 14653
rect 37829 14602 37850 14636
rect 37884 14602 37940 14636
rect 37974 14634 38030 14636
rect 38064 14634 38120 14636
rect 38154 14634 38210 14636
rect 38244 14634 38300 14636
rect 38334 14634 38390 14636
rect 38424 14634 38480 14636
rect 38514 14634 38570 14636
rect 38604 14634 38660 14636
rect 38694 14634 38750 14636
rect 37994 14602 38030 14634
rect 38084 14602 38120 14634
rect 38174 14602 38210 14634
rect 38264 14602 38300 14634
rect 38354 14602 38390 14634
rect 38444 14602 38480 14634
rect 38534 14602 38570 14634
rect 38624 14602 38660 14634
rect 38714 14602 38750 14634
rect 38784 14602 38791 14636
rect 37829 14600 37960 14602
rect 37994 14600 38050 14602
rect 38084 14600 38140 14602
rect 38174 14600 38230 14602
rect 38264 14600 38320 14602
rect 38354 14600 38410 14602
rect 38444 14600 38500 14602
rect 38534 14600 38590 14602
rect 38624 14600 38680 14602
rect 38714 14600 38791 14602
rect 37829 14581 38791 14600
rect 37829 14577 37901 14581
rect 37829 14543 37848 14577
rect 37882 14543 37901 14577
rect 37829 14487 37901 14543
rect 38719 14558 38791 14581
rect 38719 14524 38738 14558
rect 38772 14524 38791 14558
rect 37829 14453 37848 14487
rect 37882 14453 37901 14487
rect 37829 14397 37901 14453
rect 37829 14363 37848 14397
rect 37882 14363 37901 14397
rect 37829 14307 37901 14363
rect 37829 14273 37848 14307
rect 37882 14273 37901 14307
rect 37829 14217 37901 14273
rect 37829 14183 37848 14217
rect 37882 14183 37901 14217
rect 37829 14127 37901 14183
rect 37829 14093 37848 14127
rect 37882 14093 37901 14127
rect 37829 14037 37901 14093
rect 37829 14003 37848 14037
rect 37882 14003 37901 14037
rect 37829 13947 37901 14003
rect 37829 13913 37848 13947
rect 37882 13913 37901 13947
rect 37829 13857 37901 13913
rect 37829 13823 37848 13857
rect 37882 13823 37901 13857
rect 37963 14460 38657 14519
rect 37963 14426 38024 14460
rect 38058 14432 38114 14460
rect 38148 14432 38204 14460
rect 38238 14432 38294 14460
rect 38070 14426 38114 14432
rect 38170 14426 38204 14432
rect 38270 14426 38294 14432
rect 38328 14432 38384 14460
rect 38328 14426 38336 14432
rect 37963 14398 38036 14426
rect 38070 14398 38136 14426
rect 38170 14398 38236 14426
rect 38270 14398 38336 14426
rect 38370 14426 38384 14432
rect 38418 14432 38474 14460
rect 38418 14426 38436 14432
rect 38370 14398 38436 14426
rect 38470 14426 38474 14432
rect 38508 14432 38564 14460
rect 38508 14426 38536 14432
rect 38598 14426 38657 14460
rect 38470 14398 38536 14426
rect 38570 14398 38657 14426
rect 37963 14370 38657 14398
rect 37963 14336 38024 14370
rect 38058 14336 38114 14370
rect 38148 14336 38204 14370
rect 38238 14336 38294 14370
rect 38328 14336 38384 14370
rect 38418 14336 38474 14370
rect 38508 14336 38564 14370
rect 38598 14336 38657 14370
rect 37963 14332 38657 14336
rect 37963 14298 38036 14332
rect 38070 14298 38136 14332
rect 38170 14298 38236 14332
rect 38270 14298 38336 14332
rect 38370 14298 38436 14332
rect 38470 14298 38536 14332
rect 38570 14298 38657 14332
rect 37963 14280 38657 14298
rect 37963 14246 38024 14280
rect 38058 14246 38114 14280
rect 38148 14246 38204 14280
rect 38238 14246 38294 14280
rect 38328 14246 38384 14280
rect 38418 14246 38474 14280
rect 38508 14246 38564 14280
rect 38598 14246 38657 14280
rect 37963 14232 38657 14246
rect 37963 14198 38036 14232
rect 38070 14198 38136 14232
rect 38170 14198 38236 14232
rect 38270 14198 38336 14232
rect 38370 14198 38436 14232
rect 38470 14198 38536 14232
rect 38570 14198 38657 14232
rect 37963 14190 38657 14198
rect 37963 14156 38024 14190
rect 38058 14156 38114 14190
rect 38148 14156 38204 14190
rect 38238 14156 38294 14190
rect 38328 14156 38384 14190
rect 38418 14156 38474 14190
rect 38508 14156 38564 14190
rect 38598 14156 38657 14190
rect 37963 14132 38657 14156
rect 37963 14100 38036 14132
rect 38070 14100 38136 14132
rect 38170 14100 38236 14132
rect 38270 14100 38336 14132
rect 37963 14066 38024 14100
rect 38070 14098 38114 14100
rect 38170 14098 38204 14100
rect 38270 14098 38294 14100
rect 38058 14066 38114 14098
rect 38148 14066 38204 14098
rect 38238 14066 38294 14098
rect 38328 14098 38336 14100
rect 38370 14100 38436 14132
rect 38370 14098 38384 14100
rect 38328 14066 38384 14098
rect 38418 14098 38436 14100
rect 38470 14100 38536 14132
rect 38570 14100 38657 14132
rect 38470 14098 38474 14100
rect 38418 14066 38474 14098
rect 38508 14098 38536 14100
rect 38508 14066 38564 14098
rect 38598 14066 38657 14100
rect 37963 14032 38657 14066
rect 37963 14010 38036 14032
rect 38070 14010 38136 14032
rect 38170 14010 38236 14032
rect 38270 14010 38336 14032
rect 37963 13976 38024 14010
rect 38070 13998 38114 14010
rect 38170 13998 38204 14010
rect 38270 13998 38294 14010
rect 38058 13976 38114 13998
rect 38148 13976 38204 13998
rect 38238 13976 38294 13998
rect 38328 13998 38336 14010
rect 38370 14010 38436 14032
rect 38370 13998 38384 14010
rect 38328 13976 38384 13998
rect 38418 13998 38436 14010
rect 38470 14010 38536 14032
rect 38570 14010 38657 14032
rect 38470 13998 38474 14010
rect 38418 13976 38474 13998
rect 38508 13998 38536 14010
rect 38508 13976 38564 13998
rect 38598 13976 38657 14010
rect 37963 13932 38657 13976
rect 37963 13920 38036 13932
rect 38070 13920 38136 13932
rect 38170 13920 38236 13932
rect 38270 13920 38336 13932
rect 37963 13886 38024 13920
rect 38070 13898 38114 13920
rect 38170 13898 38204 13920
rect 38270 13898 38294 13920
rect 38058 13886 38114 13898
rect 38148 13886 38204 13898
rect 38238 13886 38294 13898
rect 38328 13898 38336 13920
rect 38370 13920 38436 13932
rect 38370 13898 38384 13920
rect 38328 13886 38384 13898
rect 38418 13898 38436 13920
rect 38470 13920 38536 13932
rect 38570 13920 38657 13932
rect 38470 13898 38474 13920
rect 38418 13886 38474 13898
rect 38508 13898 38536 13920
rect 38508 13886 38564 13898
rect 38598 13886 38657 13920
rect 37963 13825 38657 13886
rect 38719 14468 38791 14524
rect 38719 14434 38738 14468
rect 38772 14434 38791 14468
rect 38719 14378 38791 14434
rect 38719 14344 38738 14378
rect 38772 14344 38791 14378
rect 38719 14288 38791 14344
rect 38719 14254 38738 14288
rect 38772 14254 38791 14288
rect 38719 14198 38791 14254
rect 38719 14164 38738 14198
rect 38772 14164 38791 14198
rect 38719 14108 38791 14164
rect 38719 14074 38738 14108
rect 38772 14074 38791 14108
rect 38719 14018 38791 14074
rect 38719 13984 38738 14018
rect 38772 13984 38791 14018
rect 38719 13928 38791 13984
rect 38719 13894 38738 13928
rect 38772 13894 38791 13928
rect 38719 13838 38791 13894
rect 37829 13763 37901 13823
rect 38719 13804 38738 13838
rect 38772 13804 38791 13838
rect 38719 13763 38791 13804
rect 37829 13744 38791 13763
rect 37829 13710 37926 13744
rect 37960 13710 38016 13744
rect 38050 13710 38106 13744
rect 38140 13710 38196 13744
rect 38230 13710 38286 13744
rect 38320 13710 38376 13744
rect 38410 13710 38466 13744
rect 38500 13710 38556 13744
rect 38590 13710 38646 13744
rect 38680 13710 38791 13744
rect 37829 13691 38791 13710
rect 38855 14634 38887 14668
rect 38921 14634 38954 14668
rect 38855 14578 38954 14634
rect 38855 14544 38887 14578
rect 38921 14544 38954 14578
rect 38855 14488 38954 14544
rect 38855 14454 38887 14488
rect 38921 14454 38954 14488
rect 38855 14398 38954 14454
rect 38855 14364 38887 14398
rect 38921 14364 38954 14398
rect 38855 14308 38954 14364
rect 38855 14274 38887 14308
rect 38921 14274 38954 14308
rect 38855 14218 38954 14274
rect 38855 14184 38887 14218
rect 38921 14184 38954 14218
rect 38855 14128 38954 14184
rect 38855 14094 38887 14128
rect 38921 14094 38954 14128
rect 38855 14038 38954 14094
rect 38855 14004 38887 14038
rect 38921 14004 38954 14038
rect 38855 13948 38954 14004
rect 38855 13914 38887 13948
rect 38921 13914 38954 13948
rect 40168 14163 40784 14202
rect 40168 14061 40255 14163
rect 40697 14061 40784 14163
rect 38855 13858 38954 13914
rect 38855 13824 38887 13858
rect 38921 13824 38954 13858
rect 38855 13768 38954 13824
rect 38855 13734 38887 13768
rect 38921 13734 38954 13768
rect 37515 13644 37547 13678
rect 37581 13644 37700 13678
rect 37734 13644 37765 13678
rect 37515 13627 37765 13644
rect 38855 13678 38954 13734
rect 38855 13644 38887 13678
rect 38921 13644 38954 13678
rect 38855 13627 38954 13644
rect 28286 13594 38954 13627
rect 28286 13560 28416 13594
rect 28450 13560 28506 13594
rect 28540 13560 28596 13594
rect 28630 13560 28686 13594
rect 28720 13560 28776 13594
rect 28810 13560 28866 13594
rect 28900 13560 28956 13594
rect 28990 13560 29046 13594
rect 29080 13560 29136 13594
rect 29170 13560 29226 13594
rect 29260 13560 29316 13594
rect 29350 13560 29406 13594
rect 29440 13560 29756 13594
rect 29790 13560 29846 13594
rect 29880 13560 29936 13594
rect 29970 13560 30026 13594
rect 30060 13560 30116 13594
rect 30150 13560 30206 13594
rect 30240 13560 30296 13594
rect 30330 13560 30386 13594
rect 30420 13560 30476 13594
rect 30510 13560 30566 13594
rect 30600 13560 30656 13594
rect 30690 13560 30746 13594
rect 30780 13560 31096 13594
rect 31130 13560 31186 13594
rect 31220 13560 31276 13594
rect 31310 13560 31366 13594
rect 31400 13560 31456 13594
rect 31490 13560 31546 13594
rect 31580 13560 31636 13594
rect 31670 13560 31726 13594
rect 31760 13560 31816 13594
rect 31850 13560 31906 13594
rect 31940 13560 31996 13594
rect 32030 13560 32086 13594
rect 32120 13560 32436 13594
rect 32470 13560 32526 13594
rect 32560 13560 32616 13594
rect 32650 13560 32706 13594
rect 32740 13560 32796 13594
rect 32830 13560 32886 13594
rect 32920 13560 32976 13594
rect 33010 13560 33066 13594
rect 33100 13560 33156 13594
rect 33190 13560 33246 13594
rect 33280 13560 33336 13594
rect 33370 13560 33426 13594
rect 33460 13560 33776 13594
rect 33810 13560 33866 13594
rect 33900 13560 33956 13594
rect 33990 13560 34046 13594
rect 34080 13560 34136 13594
rect 34170 13560 34226 13594
rect 34260 13560 34316 13594
rect 34350 13560 34406 13594
rect 34440 13560 34496 13594
rect 34530 13560 34586 13594
rect 34620 13560 34676 13594
rect 34710 13560 34766 13594
rect 34800 13560 35116 13594
rect 35150 13560 35206 13594
rect 35240 13560 35296 13594
rect 35330 13560 35386 13594
rect 35420 13560 35476 13594
rect 35510 13560 35566 13594
rect 35600 13560 35656 13594
rect 35690 13560 35746 13594
rect 35780 13560 35836 13594
rect 35870 13560 35926 13594
rect 35960 13560 36016 13594
rect 36050 13560 36106 13594
rect 36140 13560 36456 13594
rect 36490 13560 36546 13594
rect 36580 13560 36636 13594
rect 36670 13560 36726 13594
rect 36760 13560 36816 13594
rect 36850 13560 36906 13594
rect 36940 13560 36996 13594
rect 37030 13560 37086 13594
rect 37120 13560 37176 13594
rect 37210 13560 37266 13594
rect 37300 13560 37356 13594
rect 37390 13560 37446 13594
rect 37480 13560 37796 13594
rect 37830 13560 37886 13594
rect 37920 13560 37976 13594
rect 38010 13560 38066 13594
rect 38100 13560 38156 13594
rect 38190 13560 38246 13594
rect 38280 13560 38336 13594
rect 38370 13560 38426 13594
rect 38460 13560 38516 13594
rect 38550 13560 38606 13594
rect 38640 13560 38696 13594
rect 38730 13560 38786 13594
rect 38820 13560 38954 13594
rect 28286 13528 38954 13560
rect 40168 13262 40784 14061
rect 41264 13917 41696 14307
rect 7896 13249 10336 13262
rect 7896 13215 8079 13249
rect 8113 13215 8279 13249
rect 8313 13215 8479 13249
rect 8513 13215 8679 13249
rect 8713 13215 8879 13249
rect 8913 13215 9079 13249
rect 9113 13215 9279 13249
rect 9313 13215 9479 13249
rect 9513 13215 9679 13249
rect 9713 13215 9879 13249
rect 9913 13215 10079 13249
rect 10113 13215 10336 13249
rect 7896 13202 10336 13215
rect 10640 13249 13080 13262
rect 10640 13215 10823 13249
rect 10857 13215 11023 13249
rect 11057 13215 11223 13249
rect 11257 13215 11423 13249
rect 11457 13215 11623 13249
rect 11657 13215 11823 13249
rect 11857 13215 12023 13249
rect 12057 13215 12223 13249
rect 12257 13215 12423 13249
rect 12457 13215 12623 13249
rect 12657 13215 12823 13249
rect 12857 13215 13080 13249
rect 10640 13202 13080 13215
rect 13384 13249 15824 13262
rect 13384 13215 13567 13249
rect 13601 13215 13767 13249
rect 13801 13215 13967 13249
rect 14001 13215 14167 13249
rect 14201 13215 14367 13249
rect 14401 13215 14567 13249
rect 14601 13215 14767 13249
rect 14801 13215 14967 13249
rect 15001 13215 15167 13249
rect 15201 13215 15367 13249
rect 15401 13215 15567 13249
rect 15601 13215 15824 13249
rect 13384 13202 15824 13215
rect 16110 13249 23278 13262
rect 16110 13215 16293 13249
rect 16327 13215 16693 13249
rect 16727 13215 17093 13249
rect 17127 13215 17493 13249
rect 17527 13215 17893 13249
rect 17927 13215 18293 13249
rect 18327 13215 18693 13249
rect 18727 13215 19093 13249
rect 19127 13215 19493 13249
rect 19527 13215 19893 13249
rect 19927 13215 20293 13249
rect 20327 13215 20693 13249
rect 20727 13215 21093 13249
rect 21127 13215 21493 13249
rect 21527 13215 21893 13249
rect 21927 13215 22293 13249
rect 22327 13215 22693 13249
rect 22727 13215 23093 13249
rect 23127 13215 23278 13249
rect 16110 13202 23278 13215
rect 23576 13249 26016 13262
rect 23576 13215 23759 13249
rect 23793 13215 23959 13249
rect 23993 13215 24159 13249
rect 24193 13215 24359 13249
rect 24393 13215 24559 13249
rect 24593 13215 24759 13249
rect 24793 13215 24959 13249
rect 24993 13215 25159 13249
rect 25193 13215 25359 13249
rect 25393 13215 25559 13249
rect 25593 13215 25759 13249
rect 25793 13215 26016 13249
rect 23576 13202 26016 13215
rect 28260 13249 38980 13262
rect 28260 13215 28443 13249
rect 28477 13215 28643 13249
rect 28677 13215 28843 13249
rect 28877 13215 29043 13249
rect 29077 13215 29243 13249
rect 29277 13215 29443 13249
rect 29477 13215 29643 13249
rect 29677 13215 29843 13249
rect 29877 13215 30043 13249
rect 30077 13215 30243 13249
rect 30277 13215 30443 13249
rect 30477 13215 30643 13249
rect 30677 13215 30843 13249
rect 30877 13215 31043 13249
rect 31077 13215 31243 13249
rect 31277 13215 31443 13249
rect 31477 13215 31643 13249
rect 31677 13215 31843 13249
rect 31877 13215 32043 13249
rect 32077 13215 32243 13249
rect 32277 13215 32443 13249
rect 32477 13215 32643 13249
rect 32677 13215 32843 13249
rect 32877 13215 33043 13249
rect 33077 13215 33243 13249
rect 33277 13215 33443 13249
rect 33477 13215 33643 13249
rect 33677 13215 33843 13249
rect 33877 13215 34043 13249
rect 34077 13215 34243 13249
rect 34277 13215 34443 13249
rect 34477 13215 34643 13249
rect 34677 13215 34843 13249
rect 34877 13215 35043 13249
rect 35077 13215 35243 13249
rect 35277 13215 35443 13249
rect 35477 13215 35643 13249
rect 35677 13215 35843 13249
rect 35877 13215 36043 13249
rect 36077 13215 36243 13249
rect 36277 13215 36443 13249
rect 36477 13215 36643 13249
rect 36677 13215 36843 13249
rect 36877 13215 37043 13249
rect 37077 13215 37243 13249
rect 37277 13215 37443 13249
rect 37477 13215 37643 13249
rect 37677 13215 37843 13249
rect 37877 13215 38043 13249
rect 38077 13215 38243 13249
rect 38277 13215 38443 13249
rect 38477 13215 38643 13249
rect 38677 13215 38843 13249
rect 38877 13215 38980 13249
rect 28260 13202 38980 13215
rect 39256 13249 41696 13262
rect 39256 13215 39439 13249
rect 39473 13215 39639 13249
rect 39673 13215 39839 13249
rect 39873 13215 40039 13249
rect 40073 13215 40239 13249
rect 40273 13215 40439 13249
rect 40473 13215 40639 13249
rect 40673 13215 40839 13249
rect 40873 13215 41039 13249
rect 41073 13215 41239 13249
rect 41273 13215 41439 13249
rect 41473 13215 41696 13249
rect 39256 13202 41696 13215
rect 7896 11369 10336 11382
rect 7896 11335 8079 11369
rect 8113 11335 8279 11369
rect 8313 11335 8479 11369
rect 8513 11335 8679 11369
rect 8713 11335 8879 11369
rect 8913 11335 9079 11369
rect 9113 11335 9279 11369
rect 9313 11335 9479 11369
rect 9513 11335 9679 11369
rect 9713 11335 9879 11369
rect 9913 11335 10079 11369
rect 10113 11335 10336 11369
rect 7896 11322 10336 11335
rect 10640 11369 13080 11382
rect 10640 11335 10823 11369
rect 10857 11335 11023 11369
rect 11057 11335 11223 11369
rect 11257 11335 11423 11369
rect 11457 11335 11623 11369
rect 11657 11335 11823 11369
rect 11857 11335 12023 11369
rect 12057 11335 12223 11369
rect 12257 11335 12423 11369
rect 12457 11335 12623 11369
rect 12657 11335 12823 11369
rect 12857 11335 13080 11369
rect 10640 11322 13080 11335
rect 13384 11369 15824 11382
rect 13384 11335 13567 11369
rect 13601 11335 13767 11369
rect 13801 11335 13967 11369
rect 14001 11335 14167 11369
rect 14201 11335 14367 11369
rect 14401 11335 14567 11369
rect 14601 11335 14767 11369
rect 14801 11335 14967 11369
rect 15001 11335 15167 11369
rect 15201 11335 15367 11369
rect 15401 11335 15567 11369
rect 15601 11335 15824 11369
rect 13384 11322 15824 11335
rect 16110 11369 23278 11382
rect 16110 11335 16293 11369
rect 16327 11335 16693 11369
rect 16727 11335 17093 11369
rect 17127 11335 17493 11369
rect 17527 11335 17893 11369
rect 17927 11335 18293 11369
rect 18327 11335 18693 11369
rect 18727 11335 19093 11369
rect 19127 11335 19493 11369
rect 19527 11335 19893 11369
rect 19927 11335 20293 11369
rect 20327 11335 20693 11369
rect 20727 11335 21093 11369
rect 21127 11335 21493 11369
rect 21527 11335 21893 11369
rect 21927 11335 22293 11369
rect 22327 11335 22693 11369
rect 22727 11335 23093 11369
rect 23127 11335 23278 11369
rect 16110 11322 23278 11335
rect 23578 11369 26590 11382
rect 23578 11335 23761 11369
rect 23795 11335 23961 11369
rect 23995 11335 24161 11369
rect 24195 11335 24361 11369
rect 24395 11335 24561 11369
rect 24595 11335 24761 11369
rect 24795 11335 24961 11369
rect 24995 11335 25161 11369
rect 25195 11335 25361 11369
rect 25395 11335 25561 11369
rect 25595 11335 25761 11369
rect 25795 11335 25961 11369
rect 25995 11335 26161 11369
rect 26195 11335 26361 11369
rect 26395 11335 26590 11369
rect 23578 11322 26590 11335
rect 26908 11369 29348 11382
rect 26908 11335 27091 11369
rect 27125 11335 27291 11369
rect 27325 11335 27491 11369
rect 27525 11335 27691 11369
rect 27725 11335 27891 11369
rect 27925 11335 28091 11369
rect 28125 11335 28291 11369
rect 28325 11335 28491 11369
rect 28525 11335 28691 11369
rect 28725 11335 28891 11369
rect 28925 11335 29091 11369
rect 29125 11335 29348 11369
rect 26908 11322 29348 11335
rect 29652 11369 32092 11382
rect 29652 11335 29835 11369
rect 29869 11335 30035 11369
rect 30069 11335 30235 11369
rect 30269 11335 30435 11369
rect 30469 11335 30635 11369
rect 30669 11335 30835 11369
rect 30869 11335 31035 11369
rect 31069 11335 31235 11369
rect 31269 11335 31435 11369
rect 31469 11335 31635 11369
rect 31669 11335 31835 11369
rect 31869 11335 32092 11369
rect 29652 11322 32092 11335
rect 32396 11369 34836 11382
rect 32396 11335 32579 11369
rect 32613 11335 32779 11369
rect 32813 11335 32979 11369
rect 33013 11335 33179 11369
rect 33213 11335 33379 11369
rect 33413 11335 33579 11369
rect 33613 11335 33779 11369
rect 33813 11335 33979 11369
rect 34013 11335 34179 11369
rect 34213 11335 34379 11369
rect 34413 11335 34579 11369
rect 34613 11335 34836 11369
rect 32396 11322 34836 11335
rect 35140 11369 37580 11382
rect 35140 11335 35323 11369
rect 35357 11335 35523 11369
rect 35557 11335 35723 11369
rect 35757 11335 35923 11369
rect 35957 11335 36123 11369
rect 36157 11335 36323 11369
rect 36357 11335 36523 11369
rect 36557 11335 36723 11369
rect 36757 11335 36923 11369
rect 36957 11335 37123 11369
rect 37157 11335 37323 11369
rect 37357 11335 37580 11369
rect 35140 11322 37580 11335
rect 37884 11369 40324 11382
rect 37884 11335 38067 11369
rect 38101 11335 38267 11369
rect 38301 11335 38467 11369
rect 38501 11335 38667 11369
rect 38701 11335 38867 11369
rect 38901 11335 39067 11369
rect 39101 11335 39267 11369
rect 39301 11335 39467 11369
rect 39501 11335 39667 11369
rect 39701 11335 39867 11369
rect 39901 11335 40067 11369
rect 40101 11335 40324 11369
rect 37884 11322 40324 11335
rect 8808 10403 9424 10442
rect 8808 10301 8895 10403
rect 9337 10301 9424 10403
rect 8808 9502 9424 10301
rect 9904 10157 10336 10547
rect 11552 10403 12168 10442
rect 11552 10301 11639 10403
rect 12081 10301 12168 10403
rect 11552 9502 12168 10301
rect 12648 10157 13080 10547
rect 14296 10403 14912 10442
rect 14296 10301 14383 10403
rect 14825 10301 14912 10403
rect 14296 9502 14912 10301
rect 15392 10157 15824 10547
rect 24776 10403 25392 10442
rect 24776 10301 24863 10403
rect 25305 10301 25392 10403
rect 24776 9502 25392 10301
rect 26159 10157 26591 10547
rect 27820 10403 28436 10442
rect 27820 10301 27907 10403
rect 28349 10301 28436 10403
rect 27820 9502 28436 10301
rect 28916 10157 29348 10547
rect 30564 10403 31180 10442
rect 30564 10301 30651 10403
rect 31093 10301 31180 10403
rect 30564 9502 31180 10301
rect 31660 10157 32092 10547
rect 33308 10403 33924 10442
rect 33308 10301 33395 10403
rect 33837 10301 33924 10403
rect 33308 9502 33924 10301
rect 34404 10157 34836 10547
rect 36052 10403 36668 10442
rect 36052 10301 36139 10403
rect 36581 10301 36668 10403
rect 36052 9502 36668 10301
rect 37148 10157 37580 10547
rect 38796 10403 39412 10442
rect 38796 10301 38883 10403
rect 39325 10301 39412 10403
rect 38796 9502 39412 10301
rect 39892 10157 40324 10547
rect 7896 9489 10336 9502
rect 7896 9455 8079 9489
rect 8113 9455 8279 9489
rect 8313 9455 8479 9489
rect 8513 9455 8679 9489
rect 8713 9455 8879 9489
rect 8913 9455 9079 9489
rect 9113 9455 9279 9489
rect 9313 9455 9479 9489
rect 9513 9455 9679 9489
rect 9713 9455 9879 9489
rect 9913 9455 10079 9489
rect 10113 9455 10336 9489
rect 7896 9442 10336 9455
rect 10640 9489 13080 9502
rect 10640 9455 10823 9489
rect 10857 9455 11023 9489
rect 11057 9455 11223 9489
rect 11257 9455 11423 9489
rect 11457 9455 11623 9489
rect 11657 9455 11823 9489
rect 11857 9455 12023 9489
rect 12057 9455 12223 9489
rect 12257 9455 12423 9489
rect 12457 9455 12623 9489
rect 12657 9455 12823 9489
rect 12857 9455 13080 9489
rect 10640 9442 13080 9455
rect 13384 9489 15824 9502
rect 13384 9455 13567 9489
rect 13601 9455 13767 9489
rect 13801 9455 13967 9489
rect 14001 9455 14167 9489
rect 14201 9455 14367 9489
rect 14401 9455 14567 9489
rect 14601 9455 14767 9489
rect 14801 9455 14967 9489
rect 15001 9455 15167 9489
rect 15201 9455 15367 9489
rect 15401 9455 15567 9489
rect 15601 9455 15824 9489
rect 13384 9442 15824 9455
rect 16110 9489 23278 9502
rect 16110 9455 16293 9489
rect 16327 9455 16693 9489
rect 16727 9455 17093 9489
rect 17127 9455 17493 9489
rect 17527 9455 17893 9489
rect 17927 9455 18293 9489
rect 18327 9455 18693 9489
rect 18727 9455 19093 9489
rect 19127 9455 19493 9489
rect 19527 9455 19893 9489
rect 19927 9455 20293 9489
rect 20327 9455 20693 9489
rect 20727 9455 21093 9489
rect 21127 9455 21493 9489
rect 21527 9455 21893 9489
rect 21927 9455 22293 9489
rect 22327 9455 22693 9489
rect 22727 9455 23093 9489
rect 23127 9455 23278 9489
rect 16110 9442 23278 9455
rect 23578 9489 26590 9502
rect 23578 9455 23761 9489
rect 23795 9455 23961 9489
rect 23995 9455 24161 9489
rect 24195 9455 24361 9489
rect 24395 9455 24561 9489
rect 24595 9455 24761 9489
rect 24795 9455 24961 9489
rect 24995 9455 25161 9489
rect 25195 9455 25361 9489
rect 25395 9455 25561 9489
rect 25595 9455 25761 9489
rect 25795 9455 25961 9489
rect 25995 9455 26161 9489
rect 26195 9455 26361 9489
rect 26395 9455 26590 9489
rect 23578 9442 26590 9455
rect 26908 9489 29348 9502
rect 26908 9455 27091 9489
rect 27125 9455 27291 9489
rect 27325 9455 27491 9489
rect 27525 9455 27691 9489
rect 27725 9455 27891 9489
rect 27925 9455 28091 9489
rect 28125 9455 28291 9489
rect 28325 9455 28491 9489
rect 28525 9455 28691 9489
rect 28725 9455 28891 9489
rect 28925 9455 29091 9489
rect 29125 9455 29348 9489
rect 26908 9442 29348 9455
rect 29652 9489 32092 9502
rect 29652 9455 29835 9489
rect 29869 9455 30035 9489
rect 30069 9455 30235 9489
rect 30269 9455 30435 9489
rect 30469 9455 30635 9489
rect 30669 9455 30835 9489
rect 30869 9455 31035 9489
rect 31069 9455 31235 9489
rect 31269 9455 31435 9489
rect 31469 9455 31635 9489
rect 31669 9455 31835 9489
rect 31869 9455 32092 9489
rect 29652 9442 32092 9455
rect 32396 9489 34836 9502
rect 32396 9455 32579 9489
rect 32613 9455 32779 9489
rect 32813 9455 32979 9489
rect 33013 9455 33179 9489
rect 33213 9455 33379 9489
rect 33413 9455 33579 9489
rect 33613 9455 33779 9489
rect 33813 9455 33979 9489
rect 34013 9455 34179 9489
rect 34213 9455 34379 9489
rect 34413 9455 34579 9489
rect 34613 9455 34836 9489
rect 32396 9442 34836 9455
rect 35140 9489 37580 9502
rect 35140 9455 35323 9489
rect 35357 9455 35523 9489
rect 35557 9455 35723 9489
rect 35757 9455 35923 9489
rect 35957 9455 36123 9489
rect 36157 9455 36323 9489
rect 36357 9455 36523 9489
rect 36557 9455 36723 9489
rect 36757 9455 36923 9489
rect 36957 9455 37123 9489
rect 37157 9455 37323 9489
rect 37357 9455 37580 9489
rect 35140 9442 37580 9455
rect 37884 9489 40324 9502
rect 37884 9455 38067 9489
rect 38101 9455 38267 9489
rect 38301 9455 38467 9489
rect 38501 9455 38667 9489
rect 38701 9455 38867 9489
rect 38901 9455 39067 9489
rect 39101 9455 39267 9489
rect 39301 9455 39467 9489
rect 39501 9455 39667 9489
rect 39701 9455 39867 9489
rect 39901 9455 40067 9489
rect 40101 9455 40324 9489
rect 37884 9442 40324 9455
rect 7896 7609 10336 7622
rect 7896 7575 8079 7609
rect 8113 7575 8279 7609
rect 8313 7575 8479 7609
rect 8513 7575 8679 7609
rect 8713 7575 8879 7609
rect 8913 7575 9079 7609
rect 9113 7575 9279 7609
rect 9313 7575 9479 7609
rect 9513 7575 9679 7609
rect 9713 7575 9879 7609
rect 9913 7575 10079 7609
rect 10113 7575 10336 7609
rect 7896 7562 10336 7575
rect 14268 7609 17280 7622
rect 14268 7575 14451 7609
rect 14485 7575 14651 7609
rect 14685 7575 14851 7609
rect 14885 7575 15051 7609
rect 15085 7575 15251 7609
rect 15285 7575 15451 7609
rect 15485 7575 15651 7609
rect 15685 7575 15851 7609
rect 15885 7575 16051 7609
rect 16085 7575 16251 7609
rect 16285 7575 16451 7609
rect 16485 7575 16651 7609
rect 16685 7575 16851 7609
rect 16885 7575 17051 7609
rect 17085 7575 17280 7609
rect 14268 7562 17280 7575
rect 17598 7609 20038 7622
rect 17598 7575 17781 7609
rect 17815 7575 17981 7609
rect 18015 7575 18181 7609
rect 18215 7575 18381 7609
rect 18415 7575 18581 7609
rect 18615 7575 18781 7609
rect 18815 7575 18981 7609
rect 19015 7575 19181 7609
rect 19215 7575 19381 7609
rect 19415 7575 19581 7609
rect 19615 7575 19781 7609
rect 19815 7575 20038 7609
rect 17598 7562 20038 7575
rect 20342 7609 22782 7622
rect 20342 7575 20525 7609
rect 20559 7575 20725 7609
rect 20759 7575 20925 7609
rect 20959 7575 21125 7609
rect 21159 7575 21325 7609
rect 21359 7575 21525 7609
rect 21559 7575 21725 7609
rect 21759 7575 21925 7609
rect 21959 7575 22125 7609
rect 22159 7575 22325 7609
rect 22359 7575 22525 7609
rect 22559 7575 22782 7609
rect 20342 7562 22782 7575
rect 23086 7609 25526 7622
rect 23086 7575 23269 7609
rect 23303 7575 23469 7609
rect 23503 7575 23669 7609
rect 23703 7575 23869 7609
rect 23903 7575 24069 7609
rect 24103 7575 24269 7609
rect 24303 7575 24469 7609
rect 24503 7575 24669 7609
rect 24703 7575 24869 7609
rect 24903 7575 25069 7609
rect 25103 7575 25269 7609
rect 25303 7575 25526 7609
rect 23086 7562 25526 7575
rect 25830 7609 28270 7622
rect 25830 7575 26013 7609
rect 26047 7575 26213 7609
rect 26247 7575 26413 7609
rect 26447 7575 26613 7609
rect 26647 7575 26813 7609
rect 26847 7575 27013 7609
rect 27047 7575 27213 7609
rect 27247 7575 27413 7609
rect 27447 7575 27613 7609
rect 27647 7575 27813 7609
rect 27847 7575 28013 7609
rect 28047 7575 28270 7609
rect 25830 7562 28270 7575
rect 28574 7609 31014 7622
rect 28574 7575 28757 7609
rect 28791 7575 28957 7609
rect 28991 7575 29157 7609
rect 29191 7575 29357 7609
rect 29391 7575 29557 7609
rect 29591 7575 29757 7609
rect 29791 7575 29957 7609
rect 29991 7575 30157 7609
rect 30191 7575 30357 7609
rect 30391 7575 30557 7609
rect 30591 7575 30757 7609
rect 30791 7575 31014 7609
rect 28574 7562 31014 7575
rect 31318 7609 33758 7622
rect 31318 7575 31501 7609
rect 31535 7575 31701 7609
rect 31735 7575 31901 7609
rect 31935 7575 32101 7609
rect 32135 7575 32301 7609
rect 32335 7575 32501 7609
rect 32535 7575 32701 7609
rect 32735 7575 32901 7609
rect 32935 7575 33101 7609
rect 33135 7575 33301 7609
rect 33335 7575 33501 7609
rect 33535 7575 33758 7609
rect 31318 7562 33758 7575
rect 35140 7609 37580 7622
rect 35140 7575 35323 7609
rect 35357 7575 35523 7609
rect 35557 7575 35723 7609
rect 35757 7575 35923 7609
rect 35957 7575 36123 7609
rect 36157 7575 36323 7609
rect 36357 7575 36523 7609
rect 36557 7575 36723 7609
rect 36757 7575 36923 7609
rect 36957 7575 37123 7609
rect 37157 7575 37323 7609
rect 37357 7575 37580 7609
rect 35140 7562 37580 7575
rect 37884 7609 40324 7622
rect 37884 7575 38067 7609
rect 38101 7575 38267 7609
rect 38301 7575 38467 7609
rect 38501 7575 38667 7609
rect 38701 7575 38867 7609
rect 38901 7575 39067 7609
rect 39101 7575 39267 7609
rect 39301 7575 39467 7609
rect 39501 7575 39667 7609
rect 39701 7575 39867 7609
rect 39901 7575 40067 7609
rect 40101 7575 40324 7609
rect 37884 7562 40324 7575
rect 8808 6643 9424 6682
rect 8808 6541 8895 6643
rect 9337 6541 9424 6643
rect 8808 5742 9424 6541
rect 9904 6397 10336 6787
rect 15466 6643 16082 6682
rect 15466 6541 15553 6643
rect 15995 6541 16082 6643
rect 15466 5742 16082 6541
rect 16849 6397 17281 6787
rect 18510 6643 19126 6682
rect 18510 6541 18597 6643
rect 19039 6541 19126 6643
rect 18510 5742 19126 6541
rect 19606 6397 20038 6787
rect 21254 6643 21870 6682
rect 21254 6541 21341 6643
rect 21783 6541 21870 6643
rect 21254 5742 21870 6541
rect 22350 6397 22782 6787
rect 23998 6643 24614 6682
rect 23998 6541 24085 6643
rect 24527 6541 24614 6643
rect 23998 5742 24614 6541
rect 25094 6397 25526 6787
rect 26742 6643 27358 6682
rect 26742 6541 26829 6643
rect 27271 6541 27358 6643
rect 26742 5742 27358 6541
rect 27838 6397 28270 6787
rect 29486 6643 30102 6682
rect 29486 6541 29573 6643
rect 30015 6541 30102 6643
rect 29486 5742 30102 6541
rect 30582 6397 31014 6787
rect 32230 6643 32846 6682
rect 32230 6541 32317 6643
rect 32759 6541 32846 6643
rect 32230 5742 32846 6541
rect 33326 6397 33758 6787
rect 36052 6643 36668 6682
rect 36052 6541 36139 6643
rect 36581 6541 36668 6643
rect 36052 5742 36668 6541
rect 37148 6397 37580 6787
rect 38796 6643 39412 6682
rect 38796 6541 38883 6643
rect 39325 6541 39412 6643
rect 38796 5742 39412 6541
rect 39892 6397 40324 6787
rect 7896 5729 10336 5742
rect 7896 5695 8079 5729
rect 8113 5695 8279 5729
rect 8313 5695 8479 5729
rect 8513 5695 8679 5729
rect 8713 5695 8879 5729
rect 8913 5695 9079 5729
rect 9113 5695 9279 5729
rect 9313 5695 9479 5729
rect 9513 5695 9679 5729
rect 9713 5695 9879 5729
rect 9913 5695 10079 5729
rect 10113 5695 10336 5729
rect 7896 5682 10336 5695
rect 14268 5729 17280 5742
rect 14268 5695 14451 5729
rect 14485 5695 14651 5729
rect 14685 5695 14851 5729
rect 14885 5695 15051 5729
rect 15085 5695 15251 5729
rect 15285 5695 15451 5729
rect 15485 5695 15651 5729
rect 15685 5695 15851 5729
rect 15885 5695 16051 5729
rect 16085 5695 16251 5729
rect 16285 5695 16451 5729
rect 16485 5695 16651 5729
rect 16685 5695 16851 5729
rect 16885 5695 17051 5729
rect 17085 5695 17280 5729
rect 14268 5682 17280 5695
rect 17598 5729 20038 5742
rect 17598 5695 17781 5729
rect 17815 5695 17981 5729
rect 18015 5695 18181 5729
rect 18215 5695 18381 5729
rect 18415 5695 18581 5729
rect 18615 5695 18781 5729
rect 18815 5695 18981 5729
rect 19015 5695 19181 5729
rect 19215 5695 19381 5729
rect 19415 5695 19581 5729
rect 19615 5695 19781 5729
rect 19815 5695 20038 5729
rect 17598 5682 20038 5695
rect 20342 5729 22782 5742
rect 20342 5695 20525 5729
rect 20559 5695 20725 5729
rect 20759 5695 20925 5729
rect 20959 5695 21125 5729
rect 21159 5695 21325 5729
rect 21359 5695 21525 5729
rect 21559 5695 21725 5729
rect 21759 5695 21925 5729
rect 21959 5695 22125 5729
rect 22159 5695 22325 5729
rect 22359 5695 22525 5729
rect 22559 5695 22782 5729
rect 20342 5682 22782 5695
rect 23086 5729 25526 5742
rect 23086 5695 23269 5729
rect 23303 5695 23469 5729
rect 23503 5695 23669 5729
rect 23703 5695 23869 5729
rect 23903 5695 24069 5729
rect 24103 5695 24269 5729
rect 24303 5695 24469 5729
rect 24503 5695 24669 5729
rect 24703 5695 24869 5729
rect 24903 5695 25069 5729
rect 25103 5695 25269 5729
rect 25303 5695 25526 5729
rect 23086 5682 25526 5695
rect 25830 5729 28270 5742
rect 25830 5695 26013 5729
rect 26047 5695 26213 5729
rect 26247 5695 26413 5729
rect 26447 5695 26613 5729
rect 26647 5695 26813 5729
rect 26847 5695 27013 5729
rect 27047 5695 27213 5729
rect 27247 5695 27413 5729
rect 27447 5695 27613 5729
rect 27647 5695 27813 5729
rect 27847 5695 28013 5729
rect 28047 5695 28270 5729
rect 25830 5682 28270 5695
rect 28574 5729 31014 5742
rect 28574 5695 28757 5729
rect 28791 5695 28957 5729
rect 28991 5695 29157 5729
rect 29191 5695 29357 5729
rect 29391 5695 29557 5729
rect 29591 5695 29757 5729
rect 29791 5695 29957 5729
rect 29991 5695 30157 5729
rect 30191 5695 30357 5729
rect 30391 5695 30557 5729
rect 30591 5695 30757 5729
rect 30791 5695 31014 5729
rect 28574 5682 31014 5695
rect 31318 5729 33758 5742
rect 31318 5695 31501 5729
rect 31535 5695 31701 5729
rect 31735 5695 31901 5729
rect 31935 5695 32101 5729
rect 32135 5695 32301 5729
rect 32335 5695 32501 5729
rect 32535 5695 32701 5729
rect 32735 5695 32901 5729
rect 32935 5695 33101 5729
rect 33135 5695 33301 5729
rect 33335 5695 33501 5729
rect 33535 5695 33758 5729
rect 31318 5682 33758 5695
rect 35140 5729 37580 5742
rect 35140 5695 35323 5729
rect 35357 5695 35523 5729
rect 35557 5695 35723 5729
rect 35757 5695 35923 5729
rect 35957 5695 36123 5729
rect 36157 5695 36323 5729
rect 36357 5695 36523 5729
rect 36557 5695 36723 5729
rect 36757 5695 36923 5729
rect 36957 5695 37123 5729
rect 37157 5695 37323 5729
rect 37357 5695 37580 5729
rect 35140 5682 37580 5695
rect 37884 5729 40324 5742
rect 37884 5695 38067 5729
rect 38101 5695 38267 5729
rect 38301 5695 38467 5729
rect 38501 5695 38667 5729
rect 38701 5695 38867 5729
rect 38901 5695 39067 5729
rect 39101 5695 39267 5729
rect 39301 5695 39467 5729
rect 39501 5695 39667 5729
rect 39701 5695 39867 5729
rect 39901 5695 40067 5729
rect 40101 5695 40324 5729
rect 37884 5682 40324 5695
<< viali >>
rect 6167 41415 6201 41449
rect 6983 41415 7017 41449
rect 7383 41415 7417 41449
rect 7783 41415 7817 41449
rect 8183 41415 8217 41449
rect 8583 41415 8617 41449
rect 8983 41415 9017 41449
rect 9383 41415 9417 41449
rect 9783 41415 9817 41449
rect 10183 41415 10217 41449
rect 10583 41415 10617 41449
rect 10983 41415 11017 41449
rect 11383 41415 11417 41449
rect 11783 41415 11817 41449
rect 12183 41415 12217 41449
rect 12583 41415 12617 41449
rect 12983 41415 13017 41449
rect 13383 41415 13417 41449
rect 13783 41415 13817 41449
rect 15213 41415 15247 41449
rect 15613 41415 15647 41449
rect 16013 41415 16047 41449
rect 16413 41415 16447 41449
rect 16813 41415 16847 41449
rect 17213 41415 17247 41449
rect 17613 41415 17647 41449
rect 18013 41415 18047 41449
rect 18413 41415 18447 41449
rect 18813 41415 18847 41449
rect 19213 41415 19247 41449
rect 19613 41415 19647 41449
rect 20013 41415 20047 41449
rect 20413 41415 20447 41449
rect 20813 41415 20847 41449
rect 21213 41415 21247 41449
rect 21613 41415 21647 41449
rect 22013 41415 22047 41449
rect 22413 41415 22447 41449
rect 22813 41415 22847 41449
rect 23213 41415 23247 41449
rect 23613 41415 23647 41449
rect 24013 41415 24047 41449
rect 24413 41415 24447 41449
rect 24813 41415 24847 41449
rect 25213 41415 25247 41449
rect 25613 41415 25647 41449
rect 26013 41415 26047 41449
rect 26413 41415 26447 41449
rect 26813 41415 26847 41449
rect 27213 41415 27247 41449
rect 27613 41415 27647 41449
rect 28013 41415 28047 41449
rect 28413 41415 28447 41449
rect 28813 41415 28847 41449
rect 29213 41415 29247 41449
rect 29613 41415 29647 41449
rect 30013 41415 30047 41449
rect 30413 41415 30447 41449
rect 30813 41415 30847 41449
rect 31213 41415 31247 41449
rect 31613 41415 31647 41449
rect 32013 41415 32047 41449
rect 32413 41415 32447 41449
rect 32813 41415 32847 41449
rect 33213 41415 33247 41449
rect 33613 41415 33647 41449
rect 34013 41415 34047 41449
rect 34413 41415 34447 41449
rect 34813 41415 34847 41449
rect 35213 41415 35247 41449
rect 35613 41415 35647 41449
rect 36013 41415 36047 41449
rect 36413 41415 36447 41449
rect 36813 41415 36847 41449
rect 37213 41415 37247 41449
rect 37613 41415 37647 41449
rect 38013 41415 38047 41449
rect 38413 41415 38447 41449
rect 38813 41415 38847 41449
rect 39213 41415 39247 41449
rect 39613 41415 39647 41449
rect 40013 41415 40047 41449
rect 40413 41415 40447 41449
rect 40813 41415 40847 41449
rect 41213 41415 41247 41449
rect 41613 41415 41647 41449
rect 42013 41415 42047 41449
rect 42413 41415 42447 41449
rect 15077 41147 15111 41181
rect 15077 41079 15111 41109
rect 15077 41075 15111 41079
rect 15077 41011 15111 41037
rect 15077 41003 15111 41011
rect 5996 40909 6030 40929
rect 5996 40895 6030 40909
rect 5996 40841 6030 40857
rect 5996 40823 6030 40841
rect 5996 40773 6030 40785
rect 5996 40751 6030 40773
rect 5996 40705 6030 40713
rect 5996 40679 6030 40705
rect 5996 40637 6030 40641
rect 5996 40607 6030 40637
rect 5996 40535 6030 40569
rect 5996 40467 6030 40497
rect 5996 40463 6030 40467
rect 5996 40399 6030 40425
rect 5996 40391 6030 40399
rect 5996 40331 6030 40353
rect 5996 40319 6030 40331
rect 5996 40263 6030 40281
rect 5996 40247 6030 40263
rect 5996 40195 6030 40209
rect 5996 40175 6030 40195
rect 6454 40909 6488 40929
rect 6454 40895 6488 40909
rect 6454 40841 6488 40857
rect 6454 40823 6488 40841
rect 6454 40773 6488 40785
rect 6454 40751 6488 40773
rect 6454 40705 6488 40713
rect 6454 40679 6488 40705
rect 6454 40637 6488 40641
rect 6454 40607 6488 40637
rect 6454 40535 6488 40569
rect 6454 40467 6488 40497
rect 6454 40463 6488 40467
rect 6454 40399 6488 40425
rect 6454 40391 6488 40399
rect 6454 40331 6488 40353
rect 6454 40319 6488 40331
rect 6454 40263 6488 40281
rect 6454 40247 6488 40263
rect 6454 40195 6488 40209
rect 6454 40175 6488 40195
rect 15077 40943 15111 40965
rect 15077 40931 15111 40943
rect 15077 40875 15111 40893
rect 15077 40859 15111 40875
rect 15077 40807 15111 40821
rect 15077 40787 15111 40807
rect 15077 40739 15111 40749
rect 15077 40715 15111 40739
rect 15077 40671 15111 40677
rect 15077 40643 15111 40671
rect 15077 40603 15111 40605
rect 15077 40571 15111 40603
rect 15077 40501 15111 40533
rect 15077 40499 15111 40501
rect 15077 40433 15111 40461
rect 15077 40427 15111 40433
rect 15077 40365 15111 40389
rect 15077 40355 15111 40365
rect 15077 40297 15111 40317
rect 15077 40283 15111 40297
rect 15077 40229 15111 40245
rect 15077 40211 15111 40229
rect 15077 40161 15111 40173
rect 15077 40139 15111 40161
rect 15077 40093 15111 40101
rect 15077 40067 15111 40093
rect 15077 40025 15111 40029
rect 15077 39995 15111 40025
rect 6469 39933 6503 39967
rect 15077 39923 15111 39957
rect 15535 41147 15569 41181
rect 15535 41079 15569 41109
rect 15535 41075 15569 41079
rect 15535 41011 15569 41037
rect 15535 41003 15569 41011
rect 15535 40943 15569 40965
rect 15535 40931 15569 40943
rect 15535 40875 15569 40893
rect 15535 40859 15569 40875
rect 15535 40807 15569 40821
rect 15535 40787 15569 40807
rect 15535 40739 15569 40749
rect 15535 40715 15569 40739
rect 15535 40671 15569 40677
rect 15535 40643 15569 40671
rect 15535 40603 15569 40605
rect 15535 40571 15569 40603
rect 15535 40501 15569 40533
rect 15535 40499 15569 40501
rect 15535 40433 15569 40461
rect 15535 40427 15569 40433
rect 15535 40365 15569 40389
rect 15535 40355 15569 40365
rect 15535 40297 15569 40317
rect 15535 40283 15569 40297
rect 15535 40229 15569 40245
rect 15535 40211 15569 40229
rect 15535 40161 15569 40173
rect 15535 40139 15569 40161
rect 15535 40093 15569 40101
rect 15535 40067 15569 40093
rect 15535 40025 15569 40029
rect 15535 39995 15569 40025
rect 15535 39923 15569 39957
rect 15993 41147 16027 41181
rect 15993 41079 16027 41109
rect 15993 41075 16027 41079
rect 15993 41011 16027 41037
rect 15993 41003 16027 41011
rect 15993 40943 16027 40965
rect 15993 40931 16027 40943
rect 15993 40875 16027 40893
rect 15993 40859 16027 40875
rect 15993 40807 16027 40821
rect 15993 40787 16027 40807
rect 15993 40739 16027 40749
rect 15993 40715 16027 40739
rect 15993 40671 16027 40677
rect 15993 40643 16027 40671
rect 15993 40603 16027 40605
rect 15993 40571 16027 40603
rect 15993 40501 16027 40533
rect 15993 40499 16027 40501
rect 15993 40433 16027 40461
rect 15993 40427 16027 40433
rect 15993 40365 16027 40389
rect 15993 40355 16027 40365
rect 15993 40297 16027 40317
rect 15993 40283 16027 40297
rect 15993 40229 16027 40245
rect 15993 40211 16027 40229
rect 15993 40161 16027 40173
rect 15993 40139 16027 40161
rect 15993 40093 16027 40101
rect 15993 40067 16027 40093
rect 15993 40025 16027 40029
rect 15993 39995 16027 40025
rect 15993 39923 16027 39957
rect 16451 41147 16485 41181
rect 16451 41079 16485 41109
rect 16451 41075 16485 41079
rect 16451 41011 16485 41037
rect 16451 41003 16485 41011
rect 16451 40943 16485 40965
rect 16451 40931 16485 40943
rect 16451 40875 16485 40893
rect 16451 40859 16485 40875
rect 16451 40807 16485 40821
rect 16451 40787 16485 40807
rect 16451 40739 16485 40749
rect 16451 40715 16485 40739
rect 16451 40671 16485 40677
rect 16451 40643 16485 40671
rect 16451 40603 16485 40605
rect 16451 40571 16485 40603
rect 16451 40501 16485 40533
rect 16451 40499 16485 40501
rect 16451 40433 16485 40461
rect 16451 40427 16485 40433
rect 16451 40365 16485 40389
rect 16451 40355 16485 40365
rect 16451 40297 16485 40317
rect 16451 40283 16485 40297
rect 16451 40229 16485 40245
rect 16451 40211 16485 40229
rect 16451 40161 16485 40173
rect 16451 40139 16485 40161
rect 16451 40093 16485 40101
rect 16451 40067 16485 40093
rect 16451 40025 16485 40029
rect 16451 39995 16485 40025
rect 16451 39923 16485 39957
rect 16909 41147 16943 41181
rect 16909 41079 16943 41109
rect 16909 41075 16943 41079
rect 16909 41011 16943 41037
rect 16909 41003 16943 41011
rect 16909 40943 16943 40965
rect 16909 40931 16943 40943
rect 16909 40875 16943 40893
rect 16909 40859 16943 40875
rect 16909 40807 16943 40821
rect 16909 40787 16943 40807
rect 16909 40739 16943 40749
rect 16909 40715 16943 40739
rect 16909 40671 16943 40677
rect 16909 40643 16943 40671
rect 16909 40603 16943 40605
rect 16909 40571 16943 40603
rect 16909 40501 16943 40533
rect 16909 40499 16943 40501
rect 16909 40433 16943 40461
rect 16909 40427 16943 40433
rect 16909 40365 16943 40389
rect 16909 40355 16943 40365
rect 16909 40297 16943 40317
rect 16909 40283 16943 40297
rect 16909 40229 16943 40245
rect 16909 40211 16943 40229
rect 16909 40161 16943 40173
rect 16909 40139 16943 40161
rect 16909 40093 16943 40101
rect 16909 40067 16943 40093
rect 16909 40025 16943 40029
rect 16909 39995 16943 40025
rect 16909 39923 16943 39957
rect 17367 41147 17401 41181
rect 17367 41079 17401 41109
rect 17367 41075 17401 41079
rect 17367 41011 17401 41037
rect 17367 41003 17401 41011
rect 17367 40943 17401 40965
rect 17367 40931 17401 40943
rect 17367 40875 17401 40893
rect 17367 40859 17401 40875
rect 17367 40807 17401 40821
rect 17367 40787 17401 40807
rect 17367 40739 17401 40749
rect 17367 40715 17401 40739
rect 17367 40671 17401 40677
rect 17367 40643 17401 40671
rect 17367 40603 17401 40605
rect 17367 40571 17401 40603
rect 17367 40501 17401 40533
rect 17367 40499 17401 40501
rect 17367 40433 17401 40461
rect 17367 40427 17401 40433
rect 17367 40365 17401 40389
rect 17367 40355 17401 40365
rect 17367 40297 17401 40317
rect 17367 40283 17401 40297
rect 17367 40229 17401 40245
rect 17367 40211 17401 40229
rect 17367 40161 17401 40173
rect 17367 40139 17401 40161
rect 17367 40093 17401 40101
rect 17367 40067 17401 40093
rect 17367 40025 17401 40029
rect 17367 39995 17401 40025
rect 17367 39923 17401 39957
rect 17825 41147 17859 41181
rect 17825 41079 17859 41109
rect 17825 41075 17859 41079
rect 17825 41011 17859 41037
rect 17825 41003 17859 41011
rect 17825 40943 17859 40965
rect 17825 40931 17859 40943
rect 17825 40875 17859 40893
rect 17825 40859 17859 40875
rect 17825 40807 17859 40821
rect 17825 40787 17859 40807
rect 17825 40739 17859 40749
rect 17825 40715 17859 40739
rect 17825 40671 17859 40677
rect 17825 40643 17859 40671
rect 17825 40603 17859 40605
rect 17825 40571 17859 40603
rect 17825 40501 17859 40533
rect 17825 40499 17859 40501
rect 17825 40433 17859 40461
rect 17825 40427 17859 40433
rect 17825 40365 17859 40389
rect 17825 40355 17859 40365
rect 17825 40297 17859 40317
rect 17825 40283 17859 40297
rect 17825 40229 17859 40245
rect 17825 40211 17859 40229
rect 17825 40161 17859 40173
rect 17825 40139 17859 40161
rect 17825 40093 17859 40101
rect 17825 40067 17859 40093
rect 17825 40025 17859 40029
rect 17825 39995 17859 40025
rect 17825 39923 17859 39957
rect 18283 41147 18317 41181
rect 18283 41079 18317 41109
rect 18283 41075 18317 41079
rect 18283 41011 18317 41037
rect 18283 41003 18317 41011
rect 18283 40943 18317 40965
rect 18283 40931 18317 40943
rect 18283 40875 18317 40893
rect 18283 40859 18317 40875
rect 18283 40807 18317 40821
rect 18283 40787 18317 40807
rect 18283 40739 18317 40749
rect 18283 40715 18317 40739
rect 18283 40671 18317 40677
rect 18283 40643 18317 40671
rect 18283 40603 18317 40605
rect 18283 40571 18317 40603
rect 18283 40501 18317 40533
rect 18283 40499 18317 40501
rect 18283 40433 18317 40461
rect 18283 40427 18317 40433
rect 18283 40365 18317 40389
rect 18283 40355 18317 40365
rect 18283 40297 18317 40317
rect 18283 40283 18317 40297
rect 18283 40229 18317 40245
rect 18283 40211 18317 40229
rect 18283 40161 18317 40173
rect 18283 40139 18317 40161
rect 18283 40093 18317 40101
rect 18283 40067 18317 40093
rect 18283 40025 18317 40029
rect 18283 39995 18317 40025
rect 18283 39923 18317 39957
rect 18741 41147 18775 41181
rect 18741 41079 18775 41109
rect 18741 41075 18775 41079
rect 18741 41011 18775 41037
rect 18741 41003 18775 41011
rect 18741 40943 18775 40965
rect 18741 40931 18775 40943
rect 18741 40875 18775 40893
rect 18741 40859 18775 40875
rect 18741 40807 18775 40821
rect 18741 40787 18775 40807
rect 18741 40739 18775 40749
rect 18741 40715 18775 40739
rect 18741 40671 18775 40677
rect 18741 40643 18775 40671
rect 18741 40603 18775 40605
rect 18741 40571 18775 40603
rect 18741 40501 18775 40533
rect 18741 40499 18775 40501
rect 18741 40433 18775 40461
rect 18741 40427 18775 40433
rect 18741 40365 18775 40389
rect 18741 40355 18775 40365
rect 18741 40297 18775 40317
rect 18741 40283 18775 40297
rect 18741 40229 18775 40245
rect 18741 40211 18775 40229
rect 18741 40161 18775 40173
rect 18741 40139 18775 40161
rect 18741 40093 18775 40101
rect 18741 40067 18775 40093
rect 18741 40025 18775 40029
rect 18741 39995 18775 40025
rect 18741 39923 18775 39957
rect 19199 41147 19233 41181
rect 19199 41079 19233 41109
rect 19199 41075 19233 41079
rect 19199 41011 19233 41037
rect 19199 41003 19233 41011
rect 19199 40943 19233 40965
rect 19199 40931 19233 40943
rect 19199 40875 19233 40893
rect 19199 40859 19233 40875
rect 19199 40807 19233 40821
rect 19199 40787 19233 40807
rect 19199 40739 19233 40749
rect 19199 40715 19233 40739
rect 19199 40671 19233 40677
rect 19199 40643 19233 40671
rect 19199 40603 19233 40605
rect 19199 40571 19233 40603
rect 19199 40501 19233 40533
rect 19199 40499 19233 40501
rect 19199 40433 19233 40461
rect 19199 40427 19233 40433
rect 19199 40365 19233 40389
rect 19199 40355 19233 40365
rect 19199 40297 19233 40317
rect 19199 40283 19233 40297
rect 19199 40229 19233 40245
rect 19199 40211 19233 40229
rect 19199 40161 19233 40173
rect 19199 40139 19233 40161
rect 19199 40093 19233 40101
rect 19199 40067 19233 40093
rect 19199 40025 19233 40029
rect 19199 39995 19233 40025
rect 19199 39923 19233 39957
rect 19657 41147 19691 41181
rect 19657 41079 19691 41109
rect 19657 41075 19691 41079
rect 19657 41011 19691 41037
rect 19657 41003 19691 41011
rect 19657 40943 19691 40965
rect 19657 40931 19691 40943
rect 19657 40875 19691 40893
rect 19657 40859 19691 40875
rect 19657 40807 19691 40821
rect 19657 40787 19691 40807
rect 19657 40739 19691 40749
rect 19657 40715 19691 40739
rect 19657 40671 19691 40677
rect 19657 40643 19691 40671
rect 19657 40603 19691 40605
rect 19657 40571 19691 40603
rect 19657 40501 19691 40533
rect 19657 40499 19691 40501
rect 19657 40433 19691 40461
rect 19657 40427 19691 40433
rect 19657 40365 19691 40389
rect 19657 40355 19691 40365
rect 19657 40297 19691 40317
rect 19657 40283 19691 40297
rect 19657 40229 19691 40245
rect 19657 40211 19691 40229
rect 19657 40161 19691 40173
rect 19657 40139 19691 40161
rect 19657 40093 19691 40101
rect 19657 40067 19691 40093
rect 19657 40025 19691 40029
rect 19657 39995 19691 40025
rect 19657 39923 19691 39957
rect 20115 41147 20149 41181
rect 20115 41079 20149 41109
rect 20115 41075 20149 41079
rect 20115 41011 20149 41037
rect 20115 41003 20149 41011
rect 20115 40943 20149 40965
rect 20115 40931 20149 40943
rect 20115 40875 20149 40893
rect 20115 40859 20149 40875
rect 20115 40807 20149 40821
rect 20115 40787 20149 40807
rect 20115 40739 20149 40749
rect 20115 40715 20149 40739
rect 20115 40671 20149 40677
rect 20115 40643 20149 40671
rect 20115 40603 20149 40605
rect 20115 40571 20149 40603
rect 20115 40501 20149 40533
rect 20115 40499 20149 40501
rect 20115 40433 20149 40461
rect 20115 40427 20149 40433
rect 20115 40365 20149 40389
rect 20115 40355 20149 40365
rect 20115 40297 20149 40317
rect 20115 40283 20149 40297
rect 20115 40229 20149 40245
rect 20115 40211 20149 40229
rect 20115 40161 20149 40173
rect 20115 40139 20149 40161
rect 20115 40093 20149 40101
rect 20115 40067 20149 40093
rect 20115 40025 20149 40029
rect 20115 39995 20149 40025
rect 20115 39923 20149 39957
rect 20573 41147 20607 41181
rect 20573 41079 20607 41109
rect 20573 41075 20607 41079
rect 20573 41011 20607 41037
rect 20573 41003 20607 41011
rect 20573 40943 20607 40965
rect 20573 40931 20607 40943
rect 20573 40875 20607 40893
rect 20573 40859 20607 40875
rect 20573 40807 20607 40821
rect 20573 40787 20607 40807
rect 20573 40739 20607 40749
rect 20573 40715 20607 40739
rect 20573 40671 20607 40677
rect 20573 40643 20607 40671
rect 20573 40603 20607 40605
rect 20573 40571 20607 40603
rect 20573 40501 20607 40533
rect 20573 40499 20607 40501
rect 20573 40433 20607 40461
rect 20573 40427 20607 40433
rect 20573 40365 20607 40389
rect 20573 40355 20607 40365
rect 20573 40297 20607 40317
rect 20573 40283 20607 40297
rect 20573 40229 20607 40245
rect 20573 40211 20607 40229
rect 20573 40161 20607 40173
rect 20573 40139 20607 40161
rect 20573 40093 20607 40101
rect 20573 40067 20607 40093
rect 20573 40025 20607 40029
rect 20573 39995 20607 40025
rect 20573 39923 20607 39957
rect 21031 41147 21065 41181
rect 21031 41079 21065 41109
rect 21031 41075 21065 41079
rect 21031 41011 21065 41037
rect 21031 41003 21065 41011
rect 21031 40943 21065 40965
rect 21031 40931 21065 40943
rect 21031 40875 21065 40893
rect 21031 40859 21065 40875
rect 21031 40807 21065 40821
rect 21031 40787 21065 40807
rect 21031 40739 21065 40749
rect 21031 40715 21065 40739
rect 21031 40671 21065 40677
rect 21031 40643 21065 40671
rect 21031 40603 21065 40605
rect 21031 40571 21065 40603
rect 21031 40501 21065 40533
rect 21031 40499 21065 40501
rect 21031 40433 21065 40461
rect 21031 40427 21065 40433
rect 21031 40365 21065 40389
rect 21031 40355 21065 40365
rect 21031 40297 21065 40317
rect 21031 40283 21065 40297
rect 21031 40229 21065 40245
rect 21031 40211 21065 40229
rect 21031 40161 21065 40173
rect 21031 40139 21065 40161
rect 21031 40093 21065 40101
rect 21031 40067 21065 40093
rect 21031 40025 21065 40029
rect 21031 39995 21065 40025
rect 21031 39923 21065 39957
rect 21489 41147 21523 41181
rect 21489 41079 21523 41109
rect 21489 41075 21523 41079
rect 21489 41011 21523 41037
rect 21489 41003 21523 41011
rect 21489 40943 21523 40965
rect 21489 40931 21523 40943
rect 21489 40875 21523 40893
rect 21489 40859 21523 40875
rect 21489 40807 21523 40821
rect 21489 40787 21523 40807
rect 21489 40739 21523 40749
rect 21489 40715 21523 40739
rect 21489 40671 21523 40677
rect 21489 40643 21523 40671
rect 21489 40603 21523 40605
rect 21489 40571 21523 40603
rect 21489 40501 21523 40533
rect 21489 40499 21523 40501
rect 21489 40433 21523 40461
rect 21489 40427 21523 40433
rect 21489 40365 21523 40389
rect 21489 40355 21523 40365
rect 21489 40297 21523 40317
rect 21489 40283 21523 40297
rect 21489 40229 21523 40245
rect 21489 40211 21523 40229
rect 21489 40161 21523 40173
rect 21489 40139 21523 40161
rect 21489 40093 21523 40101
rect 21489 40067 21523 40093
rect 21489 40025 21523 40029
rect 21489 39995 21523 40025
rect 21489 39923 21523 39957
rect 21947 41147 21981 41181
rect 21947 41079 21981 41109
rect 21947 41075 21981 41079
rect 21947 41011 21981 41037
rect 21947 41003 21981 41011
rect 21947 40943 21981 40965
rect 21947 40931 21981 40943
rect 21947 40875 21981 40893
rect 21947 40859 21981 40875
rect 21947 40807 21981 40821
rect 21947 40787 21981 40807
rect 21947 40739 21981 40749
rect 21947 40715 21981 40739
rect 21947 40671 21981 40677
rect 21947 40643 21981 40671
rect 21947 40603 21981 40605
rect 21947 40571 21981 40603
rect 21947 40501 21981 40533
rect 21947 40499 21981 40501
rect 21947 40433 21981 40461
rect 21947 40427 21981 40433
rect 21947 40365 21981 40389
rect 21947 40355 21981 40365
rect 21947 40297 21981 40317
rect 21947 40283 21981 40297
rect 21947 40229 21981 40245
rect 21947 40211 21981 40229
rect 21947 40161 21981 40173
rect 21947 40139 21981 40161
rect 21947 40093 21981 40101
rect 21947 40067 21981 40093
rect 21947 40025 21981 40029
rect 21947 39995 21981 40025
rect 21947 39923 21981 39957
rect 22405 41147 22439 41181
rect 22405 41079 22439 41109
rect 22405 41075 22439 41079
rect 22405 41011 22439 41037
rect 22405 41003 22439 41011
rect 22405 40943 22439 40965
rect 22405 40931 22439 40943
rect 22405 40875 22439 40893
rect 22405 40859 22439 40875
rect 22405 40807 22439 40821
rect 22405 40787 22439 40807
rect 22405 40739 22439 40749
rect 22405 40715 22439 40739
rect 22405 40671 22439 40677
rect 22405 40643 22439 40671
rect 22405 40603 22439 40605
rect 22405 40571 22439 40603
rect 22405 40501 22439 40533
rect 22405 40499 22439 40501
rect 22405 40433 22439 40461
rect 22405 40427 22439 40433
rect 22405 40365 22439 40389
rect 22405 40355 22439 40365
rect 22405 40297 22439 40317
rect 22405 40283 22439 40297
rect 22405 40229 22439 40245
rect 22405 40211 22439 40229
rect 22405 40161 22439 40173
rect 22405 40139 22439 40161
rect 22405 40093 22439 40101
rect 22405 40067 22439 40093
rect 22405 40025 22439 40029
rect 22405 39995 22439 40025
rect 22405 39923 22439 39957
rect 22863 41147 22897 41181
rect 22863 41079 22897 41109
rect 22863 41075 22897 41079
rect 22863 41011 22897 41037
rect 22863 41003 22897 41011
rect 22863 40943 22897 40965
rect 22863 40931 22897 40943
rect 22863 40875 22897 40893
rect 22863 40859 22897 40875
rect 22863 40807 22897 40821
rect 22863 40787 22897 40807
rect 22863 40739 22897 40749
rect 22863 40715 22897 40739
rect 22863 40671 22897 40677
rect 22863 40643 22897 40671
rect 22863 40603 22897 40605
rect 22863 40571 22897 40603
rect 22863 40501 22897 40533
rect 22863 40499 22897 40501
rect 22863 40433 22897 40461
rect 22863 40427 22897 40433
rect 22863 40365 22897 40389
rect 22863 40355 22897 40365
rect 22863 40297 22897 40317
rect 22863 40283 22897 40297
rect 22863 40229 22897 40245
rect 22863 40211 22897 40229
rect 22863 40161 22897 40173
rect 22863 40139 22897 40161
rect 22863 40093 22897 40101
rect 22863 40067 22897 40093
rect 22863 40025 22897 40029
rect 22863 39995 22897 40025
rect 22863 39923 22897 39957
rect 23321 41147 23355 41181
rect 23321 41079 23355 41109
rect 23321 41075 23355 41079
rect 23321 41011 23355 41037
rect 23321 41003 23355 41011
rect 23321 40943 23355 40965
rect 23321 40931 23355 40943
rect 23321 40875 23355 40893
rect 23321 40859 23355 40875
rect 23321 40807 23355 40821
rect 23321 40787 23355 40807
rect 23321 40739 23355 40749
rect 23321 40715 23355 40739
rect 23321 40671 23355 40677
rect 23321 40643 23355 40671
rect 23321 40603 23355 40605
rect 23321 40571 23355 40603
rect 23321 40501 23355 40533
rect 23321 40499 23355 40501
rect 23321 40433 23355 40461
rect 23321 40427 23355 40433
rect 23321 40365 23355 40389
rect 23321 40355 23355 40365
rect 23321 40297 23355 40317
rect 23321 40283 23355 40297
rect 23321 40229 23355 40245
rect 23321 40211 23355 40229
rect 23321 40161 23355 40173
rect 23321 40139 23355 40161
rect 23321 40093 23355 40101
rect 23321 40067 23355 40093
rect 23321 40025 23355 40029
rect 23321 39995 23355 40025
rect 23321 39923 23355 39957
rect 23779 41147 23813 41181
rect 23779 41079 23813 41109
rect 23779 41075 23813 41079
rect 23779 41011 23813 41037
rect 23779 41003 23813 41011
rect 23779 40943 23813 40965
rect 23779 40931 23813 40943
rect 23779 40875 23813 40893
rect 23779 40859 23813 40875
rect 23779 40807 23813 40821
rect 23779 40787 23813 40807
rect 23779 40739 23813 40749
rect 23779 40715 23813 40739
rect 23779 40671 23813 40677
rect 23779 40643 23813 40671
rect 23779 40603 23813 40605
rect 23779 40571 23813 40603
rect 23779 40501 23813 40533
rect 23779 40499 23813 40501
rect 23779 40433 23813 40461
rect 23779 40427 23813 40433
rect 23779 40365 23813 40389
rect 23779 40355 23813 40365
rect 23779 40297 23813 40317
rect 23779 40283 23813 40297
rect 23779 40229 23813 40245
rect 23779 40211 23813 40229
rect 23779 40161 23813 40173
rect 23779 40139 23813 40161
rect 23779 40093 23813 40101
rect 23779 40067 23813 40093
rect 23779 40025 23813 40029
rect 23779 39995 23813 40025
rect 23779 39923 23813 39957
rect 24237 41147 24271 41181
rect 24237 41079 24271 41109
rect 24237 41075 24271 41079
rect 24237 41011 24271 41037
rect 24237 41003 24271 41011
rect 24237 40943 24271 40965
rect 24237 40931 24271 40943
rect 24237 40875 24271 40893
rect 24237 40859 24271 40875
rect 24237 40807 24271 40821
rect 24237 40787 24271 40807
rect 24237 40739 24271 40749
rect 24237 40715 24271 40739
rect 24237 40671 24271 40677
rect 24237 40643 24271 40671
rect 24237 40603 24271 40605
rect 24237 40571 24271 40603
rect 24237 40501 24271 40533
rect 24237 40499 24271 40501
rect 24237 40433 24271 40461
rect 24237 40427 24271 40433
rect 24237 40365 24271 40389
rect 24237 40355 24271 40365
rect 24237 40297 24271 40317
rect 24237 40283 24271 40297
rect 24237 40229 24271 40245
rect 24237 40211 24271 40229
rect 24237 40161 24271 40173
rect 24237 40139 24271 40161
rect 24237 40093 24271 40101
rect 24237 40067 24271 40093
rect 24237 40025 24271 40029
rect 24237 39995 24271 40025
rect 24237 39923 24271 39957
rect 24695 41147 24729 41181
rect 24695 41079 24729 41109
rect 24695 41075 24729 41079
rect 24695 41011 24729 41037
rect 24695 41003 24729 41011
rect 24695 40943 24729 40965
rect 24695 40931 24729 40943
rect 24695 40875 24729 40893
rect 24695 40859 24729 40875
rect 24695 40807 24729 40821
rect 24695 40787 24729 40807
rect 24695 40739 24729 40749
rect 24695 40715 24729 40739
rect 24695 40671 24729 40677
rect 24695 40643 24729 40671
rect 24695 40603 24729 40605
rect 24695 40571 24729 40603
rect 24695 40501 24729 40533
rect 24695 40499 24729 40501
rect 24695 40433 24729 40461
rect 24695 40427 24729 40433
rect 24695 40365 24729 40389
rect 24695 40355 24729 40365
rect 24695 40297 24729 40317
rect 24695 40283 24729 40297
rect 24695 40229 24729 40245
rect 24695 40211 24729 40229
rect 24695 40161 24729 40173
rect 24695 40139 24729 40161
rect 24695 40093 24729 40101
rect 24695 40067 24729 40093
rect 24695 40025 24729 40029
rect 24695 39995 24729 40025
rect 24695 39923 24729 39957
rect 25153 41147 25187 41181
rect 25153 41079 25187 41109
rect 25153 41075 25187 41079
rect 25153 41011 25187 41037
rect 25153 41003 25187 41011
rect 25153 40943 25187 40965
rect 25153 40931 25187 40943
rect 25153 40875 25187 40893
rect 25153 40859 25187 40875
rect 25153 40807 25187 40821
rect 25153 40787 25187 40807
rect 25153 40739 25187 40749
rect 25153 40715 25187 40739
rect 25153 40671 25187 40677
rect 25153 40643 25187 40671
rect 25153 40603 25187 40605
rect 25153 40571 25187 40603
rect 25153 40501 25187 40533
rect 25153 40499 25187 40501
rect 25153 40433 25187 40461
rect 25153 40427 25187 40433
rect 25153 40365 25187 40389
rect 25153 40355 25187 40365
rect 25153 40297 25187 40317
rect 25153 40283 25187 40297
rect 25153 40229 25187 40245
rect 25153 40211 25187 40229
rect 25153 40161 25187 40173
rect 25153 40139 25187 40161
rect 25153 40093 25187 40101
rect 25153 40067 25187 40093
rect 25153 40025 25187 40029
rect 25153 39995 25187 40025
rect 25153 39923 25187 39957
rect 25611 41147 25645 41181
rect 25611 41079 25645 41109
rect 25611 41075 25645 41079
rect 25611 41011 25645 41037
rect 25611 41003 25645 41011
rect 25611 40943 25645 40965
rect 25611 40931 25645 40943
rect 25611 40875 25645 40893
rect 25611 40859 25645 40875
rect 25611 40807 25645 40821
rect 25611 40787 25645 40807
rect 25611 40739 25645 40749
rect 25611 40715 25645 40739
rect 25611 40671 25645 40677
rect 25611 40643 25645 40671
rect 25611 40603 25645 40605
rect 25611 40571 25645 40603
rect 25611 40501 25645 40533
rect 25611 40499 25645 40501
rect 25611 40433 25645 40461
rect 25611 40427 25645 40433
rect 25611 40365 25645 40389
rect 25611 40355 25645 40365
rect 25611 40297 25645 40317
rect 25611 40283 25645 40297
rect 25611 40229 25645 40245
rect 25611 40211 25645 40229
rect 25611 40161 25645 40173
rect 25611 40139 25645 40161
rect 25611 40093 25645 40101
rect 25611 40067 25645 40093
rect 25611 40025 25645 40029
rect 25611 39995 25645 40025
rect 25611 39923 25645 39957
rect 26069 41147 26103 41181
rect 26069 41079 26103 41109
rect 26069 41075 26103 41079
rect 26069 41011 26103 41037
rect 26069 41003 26103 41011
rect 26069 40943 26103 40965
rect 26069 40931 26103 40943
rect 26069 40875 26103 40893
rect 26069 40859 26103 40875
rect 26069 40807 26103 40821
rect 26069 40787 26103 40807
rect 26069 40739 26103 40749
rect 26069 40715 26103 40739
rect 26069 40671 26103 40677
rect 26069 40643 26103 40671
rect 26069 40603 26103 40605
rect 26069 40571 26103 40603
rect 26069 40501 26103 40533
rect 26069 40499 26103 40501
rect 26069 40433 26103 40461
rect 26069 40427 26103 40433
rect 26069 40365 26103 40389
rect 26069 40355 26103 40365
rect 26069 40297 26103 40317
rect 26069 40283 26103 40297
rect 26069 40229 26103 40245
rect 26069 40211 26103 40229
rect 26069 40161 26103 40173
rect 26069 40139 26103 40161
rect 26069 40093 26103 40101
rect 26069 40067 26103 40093
rect 26069 40025 26103 40029
rect 26069 39995 26103 40025
rect 26069 39923 26103 39957
rect 26527 41147 26561 41181
rect 26527 41079 26561 41109
rect 26527 41075 26561 41079
rect 26527 41011 26561 41037
rect 26527 41003 26561 41011
rect 26527 40943 26561 40965
rect 26527 40931 26561 40943
rect 26527 40875 26561 40893
rect 26527 40859 26561 40875
rect 26527 40807 26561 40821
rect 26527 40787 26561 40807
rect 26527 40739 26561 40749
rect 26527 40715 26561 40739
rect 26527 40671 26561 40677
rect 26527 40643 26561 40671
rect 26527 40603 26561 40605
rect 26527 40571 26561 40603
rect 26527 40501 26561 40533
rect 26527 40499 26561 40501
rect 26527 40433 26561 40461
rect 26527 40427 26561 40433
rect 26527 40365 26561 40389
rect 26527 40355 26561 40365
rect 26527 40297 26561 40317
rect 26527 40283 26561 40297
rect 26527 40229 26561 40245
rect 26527 40211 26561 40229
rect 26527 40161 26561 40173
rect 26527 40139 26561 40161
rect 26527 40093 26561 40101
rect 26527 40067 26561 40093
rect 26527 40025 26561 40029
rect 26527 39995 26561 40025
rect 26527 39923 26561 39957
rect 26985 41147 27019 41181
rect 26985 41079 27019 41109
rect 26985 41075 27019 41079
rect 26985 41011 27019 41037
rect 26985 41003 27019 41011
rect 26985 40943 27019 40965
rect 26985 40931 27019 40943
rect 26985 40875 27019 40893
rect 26985 40859 27019 40875
rect 26985 40807 27019 40821
rect 26985 40787 27019 40807
rect 26985 40739 27019 40749
rect 26985 40715 27019 40739
rect 26985 40671 27019 40677
rect 26985 40643 27019 40671
rect 26985 40603 27019 40605
rect 26985 40571 27019 40603
rect 26985 40501 27019 40533
rect 26985 40499 27019 40501
rect 26985 40433 27019 40461
rect 26985 40427 27019 40433
rect 26985 40365 27019 40389
rect 26985 40355 27019 40365
rect 26985 40297 27019 40317
rect 26985 40283 27019 40297
rect 26985 40229 27019 40245
rect 26985 40211 27019 40229
rect 26985 40161 27019 40173
rect 26985 40139 27019 40161
rect 26985 40093 27019 40101
rect 26985 40067 27019 40093
rect 26985 40025 27019 40029
rect 26985 39995 27019 40025
rect 26985 39923 27019 39957
rect 27443 41147 27477 41181
rect 27443 41079 27477 41109
rect 27443 41075 27477 41079
rect 27443 41011 27477 41037
rect 27443 41003 27477 41011
rect 27443 40943 27477 40965
rect 27443 40931 27477 40943
rect 27443 40875 27477 40893
rect 27443 40859 27477 40875
rect 27443 40807 27477 40821
rect 27443 40787 27477 40807
rect 27443 40739 27477 40749
rect 27443 40715 27477 40739
rect 27443 40671 27477 40677
rect 27443 40643 27477 40671
rect 27443 40603 27477 40605
rect 27443 40571 27477 40603
rect 27443 40501 27477 40533
rect 27443 40499 27477 40501
rect 27443 40433 27477 40461
rect 27443 40427 27477 40433
rect 27443 40365 27477 40389
rect 27443 40355 27477 40365
rect 27443 40297 27477 40317
rect 27443 40283 27477 40297
rect 27443 40229 27477 40245
rect 27443 40211 27477 40229
rect 27443 40161 27477 40173
rect 27443 40139 27477 40161
rect 27443 40093 27477 40101
rect 27443 40067 27477 40093
rect 27443 40025 27477 40029
rect 27443 39995 27477 40025
rect 27443 39923 27477 39957
rect 27901 41147 27935 41181
rect 27901 41079 27935 41109
rect 27901 41075 27935 41079
rect 27901 41011 27935 41037
rect 27901 41003 27935 41011
rect 27901 40943 27935 40965
rect 27901 40931 27935 40943
rect 27901 40875 27935 40893
rect 27901 40859 27935 40875
rect 27901 40807 27935 40821
rect 27901 40787 27935 40807
rect 27901 40739 27935 40749
rect 27901 40715 27935 40739
rect 27901 40671 27935 40677
rect 27901 40643 27935 40671
rect 27901 40603 27935 40605
rect 27901 40571 27935 40603
rect 27901 40501 27935 40533
rect 27901 40499 27935 40501
rect 27901 40433 27935 40461
rect 27901 40427 27935 40433
rect 27901 40365 27935 40389
rect 27901 40355 27935 40365
rect 27901 40297 27935 40317
rect 27901 40283 27935 40297
rect 27901 40229 27935 40245
rect 27901 40211 27935 40229
rect 27901 40161 27935 40173
rect 27901 40139 27935 40161
rect 27901 40093 27935 40101
rect 27901 40067 27935 40093
rect 27901 40025 27935 40029
rect 27901 39995 27935 40025
rect 27901 39923 27935 39957
rect 28359 41147 28393 41181
rect 28359 41079 28393 41109
rect 28359 41075 28393 41079
rect 28359 41011 28393 41037
rect 28359 41003 28393 41011
rect 28359 40943 28393 40965
rect 28359 40931 28393 40943
rect 28359 40875 28393 40893
rect 28359 40859 28393 40875
rect 28359 40807 28393 40821
rect 28359 40787 28393 40807
rect 28359 40739 28393 40749
rect 28359 40715 28393 40739
rect 28359 40671 28393 40677
rect 28359 40643 28393 40671
rect 28359 40603 28393 40605
rect 28359 40571 28393 40603
rect 28359 40501 28393 40533
rect 28359 40499 28393 40501
rect 28359 40433 28393 40461
rect 28359 40427 28393 40433
rect 28359 40365 28393 40389
rect 28359 40355 28393 40365
rect 28359 40297 28393 40317
rect 28359 40283 28393 40297
rect 28359 40229 28393 40245
rect 28359 40211 28393 40229
rect 28359 40161 28393 40173
rect 28359 40139 28393 40161
rect 28359 40093 28393 40101
rect 28359 40067 28393 40093
rect 28359 40025 28393 40029
rect 28359 39995 28393 40025
rect 28359 39923 28393 39957
rect 28817 41147 28851 41181
rect 28817 41079 28851 41109
rect 28817 41075 28851 41079
rect 28817 41011 28851 41037
rect 28817 41003 28851 41011
rect 28817 40943 28851 40965
rect 28817 40931 28851 40943
rect 28817 40875 28851 40893
rect 28817 40859 28851 40875
rect 28817 40807 28851 40821
rect 28817 40787 28851 40807
rect 28817 40739 28851 40749
rect 28817 40715 28851 40739
rect 28817 40671 28851 40677
rect 28817 40643 28851 40671
rect 28817 40603 28851 40605
rect 28817 40571 28851 40603
rect 28817 40501 28851 40533
rect 28817 40499 28851 40501
rect 28817 40433 28851 40461
rect 28817 40427 28851 40433
rect 28817 40365 28851 40389
rect 28817 40355 28851 40365
rect 28817 40297 28851 40317
rect 28817 40283 28851 40297
rect 28817 40229 28851 40245
rect 28817 40211 28851 40229
rect 28817 40161 28851 40173
rect 28817 40139 28851 40161
rect 28817 40093 28851 40101
rect 28817 40067 28851 40093
rect 28817 40025 28851 40029
rect 28817 39995 28851 40025
rect 28817 39923 28851 39957
rect 29275 41147 29309 41181
rect 29275 41079 29309 41109
rect 29275 41075 29309 41079
rect 29275 41011 29309 41037
rect 29275 41003 29309 41011
rect 29275 40943 29309 40965
rect 29275 40931 29309 40943
rect 29275 40875 29309 40893
rect 29275 40859 29309 40875
rect 29275 40807 29309 40821
rect 29275 40787 29309 40807
rect 29275 40739 29309 40749
rect 29275 40715 29309 40739
rect 29275 40671 29309 40677
rect 29275 40643 29309 40671
rect 29275 40603 29309 40605
rect 29275 40571 29309 40603
rect 29275 40501 29309 40533
rect 29275 40499 29309 40501
rect 29275 40433 29309 40461
rect 29275 40427 29309 40433
rect 29275 40365 29309 40389
rect 29275 40355 29309 40365
rect 29275 40297 29309 40317
rect 29275 40283 29309 40297
rect 29275 40229 29309 40245
rect 29275 40211 29309 40229
rect 29275 40161 29309 40173
rect 29275 40139 29309 40161
rect 29275 40093 29309 40101
rect 29275 40067 29309 40093
rect 29275 40025 29309 40029
rect 29275 39995 29309 40025
rect 29275 39923 29309 39957
rect 29733 41147 29767 41181
rect 29733 41079 29767 41109
rect 29733 41075 29767 41079
rect 29733 41011 29767 41037
rect 29733 41003 29767 41011
rect 29733 40943 29767 40965
rect 29733 40931 29767 40943
rect 29733 40875 29767 40893
rect 29733 40859 29767 40875
rect 29733 40807 29767 40821
rect 29733 40787 29767 40807
rect 29733 40739 29767 40749
rect 29733 40715 29767 40739
rect 29733 40671 29767 40677
rect 29733 40643 29767 40671
rect 29733 40603 29767 40605
rect 29733 40571 29767 40603
rect 29733 40501 29767 40533
rect 29733 40499 29767 40501
rect 29733 40433 29767 40461
rect 29733 40427 29767 40433
rect 29733 40365 29767 40389
rect 29733 40355 29767 40365
rect 29733 40297 29767 40317
rect 29733 40283 29767 40297
rect 29733 40229 29767 40245
rect 29733 40211 29767 40229
rect 29733 40161 29767 40173
rect 29733 40139 29767 40161
rect 29733 40093 29767 40101
rect 29733 40067 29767 40093
rect 29733 40025 29767 40029
rect 29733 39995 29767 40025
rect 29733 39923 29767 39957
rect 30191 41147 30225 41181
rect 30191 41079 30225 41109
rect 30191 41075 30225 41079
rect 30191 41011 30225 41037
rect 30191 41003 30225 41011
rect 30191 40943 30225 40965
rect 30191 40931 30225 40943
rect 30191 40875 30225 40893
rect 30191 40859 30225 40875
rect 30191 40807 30225 40821
rect 30191 40787 30225 40807
rect 30191 40739 30225 40749
rect 30191 40715 30225 40739
rect 30191 40671 30225 40677
rect 30191 40643 30225 40671
rect 30191 40603 30225 40605
rect 30191 40571 30225 40603
rect 30191 40501 30225 40533
rect 30191 40499 30225 40501
rect 30191 40433 30225 40461
rect 30191 40427 30225 40433
rect 30191 40365 30225 40389
rect 30191 40355 30225 40365
rect 30191 40297 30225 40317
rect 30191 40283 30225 40297
rect 30191 40229 30225 40245
rect 30191 40211 30225 40229
rect 30191 40161 30225 40173
rect 30191 40139 30225 40161
rect 30191 40093 30225 40101
rect 30191 40067 30225 40093
rect 30191 40025 30225 40029
rect 30191 39995 30225 40025
rect 30191 39923 30225 39957
rect 30649 41147 30683 41181
rect 30649 41079 30683 41109
rect 30649 41075 30683 41079
rect 30649 41011 30683 41037
rect 30649 41003 30683 41011
rect 30649 40943 30683 40965
rect 30649 40931 30683 40943
rect 30649 40875 30683 40893
rect 30649 40859 30683 40875
rect 30649 40807 30683 40821
rect 30649 40787 30683 40807
rect 30649 40739 30683 40749
rect 30649 40715 30683 40739
rect 30649 40671 30683 40677
rect 30649 40643 30683 40671
rect 30649 40603 30683 40605
rect 30649 40571 30683 40603
rect 30649 40501 30683 40533
rect 30649 40499 30683 40501
rect 30649 40433 30683 40461
rect 30649 40427 30683 40433
rect 30649 40365 30683 40389
rect 30649 40355 30683 40365
rect 30649 40297 30683 40317
rect 30649 40283 30683 40297
rect 30649 40229 30683 40245
rect 30649 40211 30683 40229
rect 30649 40161 30683 40173
rect 30649 40139 30683 40161
rect 30649 40093 30683 40101
rect 30649 40067 30683 40093
rect 30649 40025 30683 40029
rect 30649 39995 30683 40025
rect 30649 39923 30683 39957
rect 31107 41147 31141 41181
rect 31107 41079 31141 41109
rect 31107 41075 31141 41079
rect 31107 41011 31141 41037
rect 31107 41003 31141 41011
rect 31107 40943 31141 40965
rect 31107 40931 31141 40943
rect 31107 40875 31141 40893
rect 31107 40859 31141 40875
rect 31107 40807 31141 40821
rect 31107 40787 31141 40807
rect 31107 40739 31141 40749
rect 31107 40715 31141 40739
rect 31107 40671 31141 40677
rect 31107 40643 31141 40671
rect 31107 40603 31141 40605
rect 31107 40571 31141 40603
rect 31107 40501 31141 40533
rect 31107 40499 31141 40501
rect 31107 40433 31141 40461
rect 31107 40427 31141 40433
rect 31107 40365 31141 40389
rect 31107 40355 31141 40365
rect 31107 40297 31141 40317
rect 31107 40283 31141 40297
rect 31107 40229 31141 40245
rect 31107 40211 31141 40229
rect 31107 40161 31141 40173
rect 31107 40139 31141 40161
rect 31107 40093 31141 40101
rect 31107 40067 31141 40093
rect 31107 40025 31141 40029
rect 31107 39995 31141 40025
rect 31107 39923 31141 39957
rect 31565 41147 31599 41181
rect 31565 41079 31599 41109
rect 31565 41075 31599 41079
rect 31565 41011 31599 41037
rect 31565 41003 31599 41011
rect 31565 40943 31599 40965
rect 31565 40931 31599 40943
rect 31565 40875 31599 40893
rect 31565 40859 31599 40875
rect 31565 40807 31599 40821
rect 31565 40787 31599 40807
rect 31565 40739 31599 40749
rect 31565 40715 31599 40739
rect 31565 40671 31599 40677
rect 31565 40643 31599 40671
rect 31565 40603 31599 40605
rect 31565 40571 31599 40603
rect 31565 40501 31599 40533
rect 31565 40499 31599 40501
rect 31565 40433 31599 40461
rect 31565 40427 31599 40433
rect 31565 40365 31599 40389
rect 31565 40355 31599 40365
rect 31565 40297 31599 40317
rect 31565 40283 31599 40297
rect 31565 40229 31599 40245
rect 31565 40211 31599 40229
rect 31565 40161 31599 40173
rect 31565 40139 31599 40161
rect 31565 40093 31599 40101
rect 31565 40067 31599 40093
rect 31565 40025 31599 40029
rect 31565 39995 31599 40025
rect 31565 39923 31599 39957
rect 32023 41147 32057 41181
rect 32023 41079 32057 41109
rect 32023 41075 32057 41079
rect 32023 41011 32057 41037
rect 32023 41003 32057 41011
rect 32023 40943 32057 40965
rect 32023 40931 32057 40943
rect 32023 40875 32057 40893
rect 32023 40859 32057 40875
rect 32023 40807 32057 40821
rect 32023 40787 32057 40807
rect 32023 40739 32057 40749
rect 32023 40715 32057 40739
rect 32023 40671 32057 40677
rect 32023 40643 32057 40671
rect 32023 40603 32057 40605
rect 32023 40571 32057 40603
rect 32023 40501 32057 40533
rect 32023 40499 32057 40501
rect 32023 40433 32057 40461
rect 32023 40427 32057 40433
rect 32023 40365 32057 40389
rect 32023 40355 32057 40365
rect 32023 40297 32057 40317
rect 32023 40283 32057 40297
rect 32023 40229 32057 40245
rect 32023 40211 32057 40229
rect 32023 40161 32057 40173
rect 32023 40139 32057 40161
rect 32023 40093 32057 40101
rect 32023 40067 32057 40093
rect 32023 40025 32057 40029
rect 32023 39995 32057 40025
rect 32023 39923 32057 39957
rect 32481 41147 32515 41181
rect 32481 41079 32515 41109
rect 32481 41075 32515 41079
rect 32481 41011 32515 41037
rect 32481 41003 32515 41011
rect 32481 40943 32515 40965
rect 32481 40931 32515 40943
rect 32481 40875 32515 40893
rect 32481 40859 32515 40875
rect 32481 40807 32515 40821
rect 32481 40787 32515 40807
rect 32481 40739 32515 40749
rect 32481 40715 32515 40739
rect 32481 40671 32515 40677
rect 32481 40643 32515 40671
rect 32481 40603 32515 40605
rect 32481 40571 32515 40603
rect 32481 40501 32515 40533
rect 32481 40499 32515 40501
rect 32481 40433 32515 40461
rect 32481 40427 32515 40433
rect 32481 40365 32515 40389
rect 32481 40355 32515 40365
rect 32481 40297 32515 40317
rect 32481 40283 32515 40297
rect 32481 40229 32515 40245
rect 32481 40211 32515 40229
rect 32481 40161 32515 40173
rect 32481 40139 32515 40161
rect 32481 40093 32515 40101
rect 32481 40067 32515 40093
rect 32481 40025 32515 40029
rect 32481 39995 32515 40025
rect 32481 39923 32515 39957
rect 32939 41147 32973 41181
rect 32939 41079 32973 41109
rect 32939 41075 32973 41079
rect 32939 41011 32973 41037
rect 32939 41003 32973 41011
rect 32939 40943 32973 40965
rect 32939 40931 32973 40943
rect 32939 40875 32973 40893
rect 32939 40859 32973 40875
rect 32939 40807 32973 40821
rect 32939 40787 32973 40807
rect 32939 40739 32973 40749
rect 32939 40715 32973 40739
rect 32939 40671 32973 40677
rect 32939 40643 32973 40671
rect 32939 40603 32973 40605
rect 32939 40571 32973 40603
rect 32939 40501 32973 40533
rect 32939 40499 32973 40501
rect 32939 40433 32973 40461
rect 32939 40427 32973 40433
rect 32939 40365 32973 40389
rect 32939 40355 32973 40365
rect 32939 40297 32973 40317
rect 32939 40283 32973 40297
rect 32939 40229 32973 40245
rect 32939 40211 32973 40229
rect 32939 40161 32973 40173
rect 32939 40139 32973 40161
rect 32939 40093 32973 40101
rect 32939 40067 32973 40093
rect 32939 40025 32973 40029
rect 32939 39995 32973 40025
rect 32939 39923 32973 39957
rect 33397 41147 33431 41181
rect 33397 41079 33431 41109
rect 33397 41075 33431 41079
rect 33397 41011 33431 41037
rect 33397 41003 33431 41011
rect 33397 40943 33431 40965
rect 33397 40931 33431 40943
rect 33397 40875 33431 40893
rect 33397 40859 33431 40875
rect 33397 40807 33431 40821
rect 33397 40787 33431 40807
rect 33397 40739 33431 40749
rect 33397 40715 33431 40739
rect 33397 40671 33431 40677
rect 33397 40643 33431 40671
rect 33397 40603 33431 40605
rect 33397 40571 33431 40603
rect 33397 40501 33431 40533
rect 33397 40499 33431 40501
rect 33397 40433 33431 40461
rect 33397 40427 33431 40433
rect 33397 40365 33431 40389
rect 33397 40355 33431 40365
rect 33397 40297 33431 40317
rect 33397 40283 33431 40297
rect 33397 40229 33431 40245
rect 33397 40211 33431 40229
rect 33397 40161 33431 40173
rect 33397 40139 33431 40161
rect 33397 40093 33431 40101
rect 33397 40067 33431 40093
rect 33397 40025 33431 40029
rect 33397 39995 33431 40025
rect 33397 39923 33431 39957
rect 33855 41147 33889 41181
rect 33855 41079 33889 41109
rect 33855 41075 33889 41079
rect 33855 41011 33889 41037
rect 33855 41003 33889 41011
rect 33855 40943 33889 40965
rect 33855 40931 33889 40943
rect 33855 40875 33889 40893
rect 33855 40859 33889 40875
rect 33855 40807 33889 40821
rect 33855 40787 33889 40807
rect 33855 40739 33889 40749
rect 33855 40715 33889 40739
rect 33855 40671 33889 40677
rect 33855 40643 33889 40671
rect 33855 40603 33889 40605
rect 33855 40571 33889 40603
rect 33855 40501 33889 40533
rect 33855 40499 33889 40501
rect 33855 40433 33889 40461
rect 33855 40427 33889 40433
rect 33855 40365 33889 40389
rect 33855 40355 33889 40365
rect 33855 40297 33889 40317
rect 33855 40283 33889 40297
rect 33855 40229 33889 40245
rect 33855 40211 33889 40229
rect 33855 40161 33889 40173
rect 33855 40139 33889 40161
rect 33855 40093 33889 40101
rect 33855 40067 33889 40093
rect 33855 40025 33889 40029
rect 33855 39995 33889 40025
rect 33855 39923 33889 39957
rect 34313 41147 34347 41181
rect 34313 41079 34347 41109
rect 34313 41075 34347 41079
rect 34313 41011 34347 41037
rect 34313 41003 34347 41011
rect 34313 40943 34347 40965
rect 34313 40931 34347 40943
rect 34313 40875 34347 40893
rect 34313 40859 34347 40875
rect 34313 40807 34347 40821
rect 34313 40787 34347 40807
rect 34313 40739 34347 40749
rect 34313 40715 34347 40739
rect 34313 40671 34347 40677
rect 34313 40643 34347 40671
rect 34313 40603 34347 40605
rect 34313 40571 34347 40603
rect 34313 40501 34347 40533
rect 34313 40499 34347 40501
rect 34313 40433 34347 40461
rect 34313 40427 34347 40433
rect 34313 40365 34347 40389
rect 34313 40355 34347 40365
rect 34313 40297 34347 40317
rect 34313 40283 34347 40297
rect 34313 40229 34347 40245
rect 34313 40211 34347 40229
rect 34313 40161 34347 40173
rect 34313 40139 34347 40161
rect 34313 40093 34347 40101
rect 34313 40067 34347 40093
rect 34313 40025 34347 40029
rect 34313 39995 34347 40025
rect 34313 39923 34347 39957
rect 34771 41147 34805 41181
rect 34771 41079 34805 41109
rect 34771 41075 34805 41079
rect 34771 41011 34805 41037
rect 34771 41003 34805 41011
rect 34771 40943 34805 40965
rect 34771 40931 34805 40943
rect 34771 40875 34805 40893
rect 34771 40859 34805 40875
rect 34771 40807 34805 40821
rect 34771 40787 34805 40807
rect 34771 40739 34805 40749
rect 34771 40715 34805 40739
rect 34771 40671 34805 40677
rect 34771 40643 34805 40671
rect 34771 40603 34805 40605
rect 34771 40571 34805 40603
rect 34771 40501 34805 40533
rect 34771 40499 34805 40501
rect 34771 40433 34805 40461
rect 34771 40427 34805 40433
rect 34771 40365 34805 40389
rect 34771 40355 34805 40365
rect 34771 40297 34805 40317
rect 34771 40283 34805 40297
rect 34771 40229 34805 40245
rect 34771 40211 34805 40229
rect 34771 40161 34805 40173
rect 34771 40139 34805 40161
rect 34771 40093 34805 40101
rect 34771 40067 34805 40093
rect 34771 40025 34805 40029
rect 34771 39995 34805 40025
rect 34771 39923 34805 39957
rect 35229 41147 35263 41181
rect 35229 41079 35263 41109
rect 35229 41075 35263 41079
rect 35229 41011 35263 41037
rect 35229 41003 35263 41011
rect 35229 40943 35263 40965
rect 35229 40931 35263 40943
rect 35229 40875 35263 40893
rect 35229 40859 35263 40875
rect 35229 40807 35263 40821
rect 35229 40787 35263 40807
rect 35229 40739 35263 40749
rect 35229 40715 35263 40739
rect 35229 40671 35263 40677
rect 35229 40643 35263 40671
rect 35229 40603 35263 40605
rect 35229 40571 35263 40603
rect 35229 40501 35263 40533
rect 35229 40499 35263 40501
rect 35229 40433 35263 40461
rect 35229 40427 35263 40433
rect 35229 40365 35263 40389
rect 35229 40355 35263 40365
rect 35229 40297 35263 40317
rect 35229 40283 35263 40297
rect 35229 40229 35263 40245
rect 35229 40211 35263 40229
rect 35229 40161 35263 40173
rect 35229 40139 35263 40161
rect 35229 40093 35263 40101
rect 35229 40067 35263 40093
rect 35229 40025 35263 40029
rect 35229 39995 35263 40025
rect 35229 39923 35263 39957
rect 35687 41147 35721 41181
rect 35687 41079 35721 41109
rect 35687 41075 35721 41079
rect 35687 41011 35721 41037
rect 35687 41003 35721 41011
rect 35687 40943 35721 40965
rect 35687 40931 35721 40943
rect 35687 40875 35721 40893
rect 35687 40859 35721 40875
rect 35687 40807 35721 40821
rect 35687 40787 35721 40807
rect 35687 40739 35721 40749
rect 35687 40715 35721 40739
rect 35687 40671 35721 40677
rect 35687 40643 35721 40671
rect 35687 40603 35721 40605
rect 35687 40571 35721 40603
rect 35687 40501 35721 40533
rect 35687 40499 35721 40501
rect 35687 40433 35721 40461
rect 35687 40427 35721 40433
rect 35687 40365 35721 40389
rect 35687 40355 35721 40365
rect 35687 40297 35721 40317
rect 35687 40283 35721 40297
rect 35687 40229 35721 40245
rect 35687 40211 35721 40229
rect 35687 40161 35721 40173
rect 35687 40139 35721 40161
rect 35687 40093 35721 40101
rect 35687 40067 35721 40093
rect 35687 40025 35721 40029
rect 35687 39995 35721 40025
rect 35687 39923 35721 39957
rect 36145 41147 36179 41181
rect 36145 41079 36179 41109
rect 36145 41075 36179 41079
rect 36145 41011 36179 41037
rect 36145 41003 36179 41011
rect 36145 40943 36179 40965
rect 36145 40931 36179 40943
rect 36145 40875 36179 40893
rect 36145 40859 36179 40875
rect 36145 40807 36179 40821
rect 36145 40787 36179 40807
rect 36145 40739 36179 40749
rect 36145 40715 36179 40739
rect 36145 40671 36179 40677
rect 36145 40643 36179 40671
rect 36145 40603 36179 40605
rect 36145 40571 36179 40603
rect 36145 40501 36179 40533
rect 36145 40499 36179 40501
rect 36145 40433 36179 40461
rect 36145 40427 36179 40433
rect 36145 40365 36179 40389
rect 36145 40355 36179 40365
rect 36145 40297 36179 40317
rect 36145 40283 36179 40297
rect 36145 40229 36179 40245
rect 36145 40211 36179 40229
rect 36145 40161 36179 40173
rect 36145 40139 36179 40161
rect 36145 40093 36179 40101
rect 36145 40067 36179 40093
rect 36145 40025 36179 40029
rect 36145 39995 36179 40025
rect 36145 39923 36179 39957
rect 36603 41147 36637 41181
rect 36603 41079 36637 41109
rect 36603 41075 36637 41079
rect 36603 41011 36637 41037
rect 36603 41003 36637 41011
rect 36603 40943 36637 40965
rect 36603 40931 36637 40943
rect 36603 40875 36637 40893
rect 36603 40859 36637 40875
rect 36603 40807 36637 40821
rect 36603 40787 36637 40807
rect 36603 40739 36637 40749
rect 36603 40715 36637 40739
rect 36603 40671 36637 40677
rect 36603 40643 36637 40671
rect 36603 40603 36637 40605
rect 36603 40571 36637 40603
rect 36603 40501 36637 40533
rect 36603 40499 36637 40501
rect 36603 40433 36637 40461
rect 36603 40427 36637 40433
rect 36603 40365 36637 40389
rect 36603 40355 36637 40365
rect 36603 40297 36637 40317
rect 36603 40283 36637 40297
rect 36603 40229 36637 40245
rect 36603 40211 36637 40229
rect 36603 40161 36637 40173
rect 36603 40139 36637 40161
rect 36603 40093 36637 40101
rect 36603 40067 36637 40093
rect 36603 40025 36637 40029
rect 36603 39995 36637 40025
rect 36603 39923 36637 39957
rect 37061 41147 37095 41181
rect 37061 41079 37095 41109
rect 37061 41075 37095 41079
rect 37061 41011 37095 41037
rect 37061 41003 37095 41011
rect 37061 40943 37095 40965
rect 37061 40931 37095 40943
rect 37061 40875 37095 40893
rect 37061 40859 37095 40875
rect 37061 40807 37095 40821
rect 37061 40787 37095 40807
rect 37061 40739 37095 40749
rect 37061 40715 37095 40739
rect 37061 40671 37095 40677
rect 37061 40643 37095 40671
rect 37061 40603 37095 40605
rect 37061 40571 37095 40603
rect 37061 40501 37095 40533
rect 37061 40499 37095 40501
rect 37061 40433 37095 40461
rect 37061 40427 37095 40433
rect 37061 40365 37095 40389
rect 37061 40355 37095 40365
rect 37061 40297 37095 40317
rect 37061 40283 37095 40297
rect 37061 40229 37095 40245
rect 37061 40211 37095 40229
rect 37061 40161 37095 40173
rect 37061 40139 37095 40161
rect 37061 40093 37095 40101
rect 37061 40067 37095 40093
rect 37061 40025 37095 40029
rect 37061 39995 37095 40025
rect 37061 39923 37095 39957
rect 37519 41147 37553 41181
rect 37519 41079 37553 41109
rect 37519 41075 37553 41079
rect 37519 41011 37553 41037
rect 37519 41003 37553 41011
rect 37519 40943 37553 40965
rect 37519 40931 37553 40943
rect 37519 40875 37553 40893
rect 37519 40859 37553 40875
rect 37519 40807 37553 40821
rect 37519 40787 37553 40807
rect 37519 40739 37553 40749
rect 37519 40715 37553 40739
rect 37519 40671 37553 40677
rect 37519 40643 37553 40671
rect 37519 40603 37553 40605
rect 37519 40571 37553 40603
rect 37519 40501 37553 40533
rect 37519 40499 37553 40501
rect 37519 40433 37553 40461
rect 37519 40427 37553 40433
rect 37519 40365 37553 40389
rect 37519 40355 37553 40365
rect 37519 40297 37553 40317
rect 37519 40283 37553 40297
rect 37519 40229 37553 40245
rect 37519 40211 37553 40229
rect 37519 40161 37553 40173
rect 37519 40139 37553 40161
rect 37519 40093 37553 40101
rect 37519 40067 37553 40093
rect 37519 40025 37553 40029
rect 37519 39995 37553 40025
rect 37519 39923 37553 39957
rect 37977 41147 38011 41181
rect 37977 41079 38011 41109
rect 37977 41075 38011 41079
rect 37977 41011 38011 41037
rect 37977 41003 38011 41011
rect 37977 40943 38011 40965
rect 37977 40931 38011 40943
rect 37977 40875 38011 40893
rect 37977 40859 38011 40875
rect 37977 40807 38011 40821
rect 37977 40787 38011 40807
rect 37977 40739 38011 40749
rect 37977 40715 38011 40739
rect 37977 40671 38011 40677
rect 37977 40643 38011 40671
rect 37977 40603 38011 40605
rect 37977 40571 38011 40603
rect 37977 40501 38011 40533
rect 37977 40499 38011 40501
rect 37977 40433 38011 40461
rect 37977 40427 38011 40433
rect 37977 40365 38011 40389
rect 37977 40355 38011 40365
rect 37977 40297 38011 40317
rect 37977 40283 38011 40297
rect 37977 40229 38011 40245
rect 37977 40211 38011 40229
rect 37977 40161 38011 40173
rect 37977 40139 38011 40161
rect 37977 40093 38011 40101
rect 37977 40067 38011 40093
rect 37977 40025 38011 40029
rect 37977 39995 38011 40025
rect 37977 39923 38011 39957
rect 38435 41147 38469 41181
rect 38435 41079 38469 41109
rect 38435 41075 38469 41079
rect 38435 41011 38469 41037
rect 38435 41003 38469 41011
rect 38435 40943 38469 40965
rect 38435 40931 38469 40943
rect 38435 40875 38469 40893
rect 38435 40859 38469 40875
rect 38435 40807 38469 40821
rect 38435 40787 38469 40807
rect 38435 40739 38469 40749
rect 38435 40715 38469 40739
rect 38435 40671 38469 40677
rect 38435 40643 38469 40671
rect 38435 40603 38469 40605
rect 38435 40571 38469 40603
rect 38435 40501 38469 40533
rect 38435 40499 38469 40501
rect 38435 40433 38469 40461
rect 38435 40427 38469 40433
rect 38435 40365 38469 40389
rect 38435 40355 38469 40365
rect 38435 40297 38469 40317
rect 38435 40283 38469 40297
rect 38435 40229 38469 40245
rect 38435 40211 38469 40229
rect 38435 40161 38469 40173
rect 38435 40139 38469 40161
rect 38435 40093 38469 40101
rect 38435 40067 38469 40093
rect 38435 40025 38469 40029
rect 38435 39995 38469 40025
rect 38435 39923 38469 39957
rect 38893 41147 38927 41181
rect 38893 41079 38927 41109
rect 38893 41075 38927 41079
rect 38893 41011 38927 41037
rect 38893 41003 38927 41011
rect 38893 40943 38927 40965
rect 38893 40931 38927 40943
rect 38893 40875 38927 40893
rect 38893 40859 38927 40875
rect 38893 40807 38927 40821
rect 38893 40787 38927 40807
rect 38893 40739 38927 40749
rect 38893 40715 38927 40739
rect 38893 40671 38927 40677
rect 38893 40643 38927 40671
rect 38893 40603 38927 40605
rect 38893 40571 38927 40603
rect 38893 40501 38927 40533
rect 38893 40499 38927 40501
rect 38893 40433 38927 40461
rect 38893 40427 38927 40433
rect 38893 40365 38927 40389
rect 38893 40355 38927 40365
rect 38893 40297 38927 40317
rect 38893 40283 38927 40297
rect 38893 40229 38927 40245
rect 38893 40211 38927 40229
rect 38893 40161 38927 40173
rect 38893 40139 38927 40161
rect 38893 40093 38927 40101
rect 38893 40067 38927 40093
rect 38893 40025 38927 40029
rect 38893 39995 38927 40025
rect 38893 39923 38927 39957
rect 38669 39797 38703 39831
rect 39351 41147 39385 41181
rect 39351 41079 39385 41109
rect 39351 41075 39385 41079
rect 39351 41011 39385 41037
rect 39351 41003 39385 41011
rect 39351 40943 39385 40965
rect 39351 40931 39385 40943
rect 39351 40875 39385 40893
rect 39351 40859 39385 40875
rect 39351 40807 39385 40821
rect 39351 40787 39385 40807
rect 39351 40739 39385 40749
rect 39351 40715 39385 40739
rect 39351 40671 39385 40677
rect 39351 40643 39385 40671
rect 39351 40603 39385 40605
rect 39351 40571 39385 40603
rect 39351 40501 39385 40533
rect 39351 40499 39385 40501
rect 39351 40433 39385 40461
rect 39351 40427 39385 40433
rect 39351 40365 39385 40389
rect 39351 40355 39385 40365
rect 39351 40297 39385 40317
rect 39351 40283 39385 40297
rect 39351 40229 39385 40245
rect 39351 40211 39385 40229
rect 39351 40161 39385 40173
rect 39351 40139 39385 40161
rect 39351 40093 39385 40101
rect 39351 40067 39385 40093
rect 39351 40025 39385 40029
rect 39351 39995 39385 40025
rect 39351 39923 39385 39957
rect 39809 41147 39843 41181
rect 39809 41079 39843 41109
rect 39809 41075 39843 41079
rect 39809 41011 39843 41037
rect 39809 41003 39843 41011
rect 39809 40943 39843 40965
rect 39809 40931 39843 40943
rect 39809 40875 39843 40893
rect 39809 40859 39843 40875
rect 39809 40807 39843 40821
rect 39809 40787 39843 40807
rect 39809 40739 39843 40749
rect 39809 40715 39843 40739
rect 39809 40671 39843 40677
rect 39809 40643 39843 40671
rect 39809 40603 39843 40605
rect 39809 40571 39843 40603
rect 39809 40501 39843 40533
rect 39809 40499 39843 40501
rect 39809 40433 39843 40461
rect 39809 40427 39843 40433
rect 39809 40365 39843 40389
rect 39809 40355 39843 40365
rect 39809 40297 39843 40317
rect 39809 40283 39843 40297
rect 39809 40229 39843 40245
rect 39809 40211 39843 40229
rect 39809 40161 39843 40173
rect 39809 40139 39843 40161
rect 39809 40093 39843 40101
rect 39809 40067 39843 40093
rect 39809 40025 39843 40029
rect 39809 39995 39843 40025
rect 39809 39923 39843 39957
rect 40267 41147 40301 41181
rect 40267 41079 40301 41109
rect 40267 41075 40301 41079
rect 40267 41011 40301 41037
rect 40267 41003 40301 41011
rect 40267 40943 40301 40965
rect 40267 40931 40301 40943
rect 40267 40875 40301 40893
rect 40267 40859 40301 40875
rect 40267 40807 40301 40821
rect 40267 40787 40301 40807
rect 40267 40739 40301 40749
rect 40267 40715 40301 40739
rect 40267 40671 40301 40677
rect 40267 40643 40301 40671
rect 40267 40603 40301 40605
rect 40267 40571 40301 40603
rect 40267 40501 40301 40533
rect 40267 40499 40301 40501
rect 40267 40433 40301 40461
rect 40267 40427 40301 40433
rect 40267 40365 40301 40389
rect 40267 40355 40301 40365
rect 40267 40297 40301 40317
rect 40267 40283 40301 40297
rect 40267 40229 40301 40245
rect 40267 40211 40301 40229
rect 40267 40161 40301 40173
rect 40267 40139 40301 40161
rect 40267 40093 40301 40101
rect 40267 40067 40301 40093
rect 40267 40025 40301 40029
rect 40267 39995 40301 40025
rect 40267 39923 40301 39957
rect 40725 41147 40759 41181
rect 40725 41079 40759 41109
rect 40725 41075 40759 41079
rect 40725 41011 40759 41037
rect 40725 41003 40759 41011
rect 40725 40943 40759 40965
rect 40725 40931 40759 40943
rect 40725 40875 40759 40893
rect 40725 40859 40759 40875
rect 40725 40807 40759 40821
rect 40725 40787 40759 40807
rect 40725 40739 40759 40749
rect 40725 40715 40759 40739
rect 40725 40671 40759 40677
rect 40725 40643 40759 40671
rect 40725 40603 40759 40605
rect 40725 40571 40759 40603
rect 40725 40501 40759 40533
rect 40725 40499 40759 40501
rect 40725 40433 40759 40461
rect 40725 40427 40759 40433
rect 40725 40365 40759 40389
rect 40725 40355 40759 40365
rect 40725 40297 40759 40317
rect 40725 40283 40759 40297
rect 40725 40229 40759 40245
rect 40725 40211 40759 40229
rect 40725 40161 40759 40173
rect 40725 40139 40759 40161
rect 40725 40093 40759 40101
rect 40725 40067 40759 40093
rect 40725 40025 40759 40029
rect 40725 39995 40759 40025
rect 40725 39923 40759 39957
rect 41183 41147 41217 41181
rect 41183 41079 41217 41109
rect 41183 41075 41217 41079
rect 41183 41011 41217 41037
rect 41183 41003 41217 41011
rect 41183 40943 41217 40965
rect 41183 40931 41217 40943
rect 41183 40875 41217 40893
rect 41183 40859 41217 40875
rect 41183 40807 41217 40821
rect 41183 40787 41217 40807
rect 41183 40739 41217 40749
rect 41183 40715 41217 40739
rect 41183 40671 41217 40677
rect 41183 40643 41217 40671
rect 41183 40603 41217 40605
rect 41183 40571 41217 40603
rect 41183 40501 41217 40533
rect 41183 40499 41217 40501
rect 41183 40433 41217 40461
rect 41183 40427 41217 40433
rect 41183 40365 41217 40389
rect 41183 40355 41217 40365
rect 41183 40297 41217 40317
rect 41183 40283 41217 40297
rect 41183 40229 41217 40245
rect 41183 40211 41217 40229
rect 41183 40161 41217 40173
rect 41183 40139 41217 40161
rect 41183 40093 41217 40101
rect 41183 40067 41217 40093
rect 41183 40025 41217 40029
rect 41183 39995 41217 40025
rect 41183 39923 41217 39957
rect 41641 41147 41675 41181
rect 41641 41079 41675 41109
rect 41641 41075 41675 41079
rect 41641 41011 41675 41037
rect 41641 41003 41675 41011
rect 41641 40943 41675 40965
rect 41641 40931 41675 40943
rect 41641 40875 41675 40893
rect 41641 40859 41675 40875
rect 41641 40807 41675 40821
rect 41641 40787 41675 40807
rect 41641 40739 41675 40749
rect 41641 40715 41675 40739
rect 41641 40671 41675 40677
rect 41641 40643 41675 40671
rect 41641 40603 41675 40605
rect 41641 40571 41675 40603
rect 41641 40501 41675 40533
rect 41641 40499 41675 40501
rect 41641 40433 41675 40461
rect 41641 40427 41675 40433
rect 41641 40365 41675 40389
rect 41641 40355 41675 40365
rect 41641 40297 41675 40317
rect 41641 40283 41675 40297
rect 41641 40229 41675 40245
rect 41641 40211 41675 40229
rect 41641 40161 41675 40173
rect 41641 40139 41675 40161
rect 41641 40093 41675 40101
rect 41641 40067 41675 40093
rect 41641 40025 41675 40029
rect 41641 39995 41675 40025
rect 41641 39923 41675 39957
rect 42099 41147 42133 41181
rect 42099 41079 42133 41109
rect 42099 41075 42133 41079
rect 42099 41011 42133 41037
rect 42099 41003 42133 41011
rect 42099 40943 42133 40965
rect 42099 40931 42133 40943
rect 42099 40875 42133 40893
rect 42099 40859 42133 40875
rect 42099 40807 42133 40821
rect 42099 40787 42133 40807
rect 42099 40739 42133 40749
rect 42099 40715 42133 40739
rect 42099 40671 42133 40677
rect 42099 40643 42133 40671
rect 42099 40603 42133 40605
rect 42099 40571 42133 40603
rect 42099 40501 42133 40533
rect 42099 40499 42133 40501
rect 42099 40433 42133 40461
rect 42099 40427 42133 40433
rect 42099 40365 42133 40389
rect 42099 40355 42133 40365
rect 42099 40297 42133 40317
rect 42099 40283 42133 40297
rect 42099 40229 42133 40245
rect 42099 40211 42133 40229
rect 42099 40161 42133 40173
rect 42099 40139 42133 40161
rect 42099 40093 42133 40101
rect 42099 40067 42133 40093
rect 42099 40025 42133 40029
rect 42099 39995 42133 40025
rect 42099 39923 42133 39957
rect 42557 41147 42591 41181
rect 42557 41079 42591 41109
rect 42557 41075 42591 41079
rect 42557 41011 42591 41037
rect 42557 41003 42591 41011
rect 42557 40943 42591 40965
rect 42557 40931 42591 40943
rect 42557 40875 42591 40893
rect 42557 40859 42591 40875
rect 42557 40807 42591 40821
rect 42557 40787 42591 40807
rect 42557 40739 42591 40749
rect 42557 40715 42591 40739
rect 42557 40671 42591 40677
rect 42557 40643 42591 40671
rect 42557 40603 42591 40605
rect 42557 40571 42591 40603
rect 42557 40501 42591 40533
rect 42557 40499 42591 40501
rect 42557 40433 42591 40461
rect 42557 40427 42591 40433
rect 42557 40365 42591 40389
rect 42557 40355 42591 40365
rect 42557 40297 42591 40317
rect 42557 40283 42591 40297
rect 42557 40229 42591 40245
rect 42557 40211 42591 40229
rect 42557 40161 42591 40173
rect 42557 40139 42591 40161
rect 42557 40093 42591 40101
rect 42557 40067 42591 40093
rect 42557 40025 42591 40029
rect 42557 39995 42591 40025
rect 42557 39923 42591 39957
rect 6469 39729 6503 39763
rect 15025 39661 15059 39695
rect 27629 39669 27647 39695
rect 27647 39669 27663 39695
rect 27629 39661 27663 39669
rect 6167 39535 6201 39569
rect 6983 39535 7017 39569
rect 7383 39535 7417 39569
rect 7783 39535 7817 39569
rect 8183 39535 8217 39569
rect 8583 39535 8617 39569
rect 8983 39535 9017 39569
rect 9383 39535 9417 39569
rect 9783 39535 9817 39569
rect 10183 39535 10217 39569
rect 10583 39535 10617 39569
rect 10983 39535 11017 39569
rect 11383 39535 11417 39569
rect 11783 39535 11817 39569
rect 12183 39535 12217 39569
rect 12583 39535 12617 39569
rect 12983 39535 13017 39569
rect 13383 39535 13417 39569
rect 13783 39535 13817 39569
rect 15213 39535 15247 39569
rect 15613 39535 15647 39569
rect 16013 39535 16047 39569
rect 16413 39535 16447 39569
rect 16813 39535 16847 39569
rect 17213 39535 17247 39569
rect 17613 39535 17647 39569
rect 18013 39535 18047 39569
rect 18413 39535 18447 39569
rect 18813 39535 18847 39569
rect 19213 39535 19247 39569
rect 19613 39535 19647 39569
rect 20013 39535 20047 39569
rect 20413 39535 20447 39569
rect 20813 39535 20847 39569
rect 21213 39535 21247 39569
rect 21613 39535 21647 39569
rect 22013 39535 22047 39569
rect 22413 39535 22447 39569
rect 22813 39535 22847 39569
rect 23213 39535 23247 39569
rect 23613 39535 23647 39569
rect 24013 39535 24047 39569
rect 24413 39535 24447 39569
rect 24813 39535 24847 39569
rect 25213 39535 25247 39569
rect 25613 39535 25647 39569
rect 26013 39535 26047 39569
rect 26413 39535 26447 39569
rect 26813 39535 26847 39569
rect 27213 39535 27247 39569
rect 27613 39535 27647 39569
rect 28013 39535 28047 39569
rect 28413 39535 28447 39569
rect 28813 39535 28847 39569
rect 29213 39535 29247 39569
rect 29613 39535 29647 39569
rect 30013 39535 30047 39569
rect 30413 39535 30447 39569
rect 30813 39535 30847 39569
rect 31213 39535 31247 39569
rect 31613 39535 31647 39569
rect 32013 39535 32047 39569
rect 32413 39535 32447 39569
rect 32813 39535 32847 39569
rect 33213 39535 33247 39569
rect 33613 39535 33647 39569
rect 34013 39535 34047 39569
rect 34413 39535 34447 39569
rect 34813 39535 34847 39569
rect 35213 39535 35247 39569
rect 35613 39535 35647 39569
rect 36013 39535 36047 39569
rect 36413 39535 36447 39569
rect 36813 39535 36847 39569
rect 37213 39535 37247 39569
rect 37613 39535 37647 39569
rect 38013 39535 38047 39569
rect 38413 39535 38447 39569
rect 38813 39535 38847 39569
rect 39213 39535 39247 39569
rect 39613 39535 39647 39569
rect 40013 39535 40047 39569
rect 40413 39535 40447 39569
rect 40813 39535 40847 39569
rect 41213 39535 41247 39569
rect 41613 39535 41647 39569
rect 42013 39535 42047 39569
rect 42413 39535 42447 39569
rect 6101 37655 6135 37689
rect 6501 37655 6535 37689
rect 6901 37655 6935 37689
rect 7301 37655 7335 37689
rect 7701 37655 7735 37689
rect 8101 37655 8135 37689
rect 8501 37655 8535 37689
rect 8901 37655 8935 37689
rect 9301 37655 9335 37689
rect 9701 37655 9735 37689
rect 10101 37655 10135 37689
rect 10501 37655 10535 37689
rect 10901 37655 10935 37689
rect 11301 37655 11335 37689
rect 11701 37655 11735 37689
rect 12101 37655 12135 37689
rect 12501 37655 12535 37689
rect 12901 37655 12935 37689
rect 13549 37655 13583 37689
rect 13949 37655 13983 37689
rect 14349 37655 14383 37689
rect 14749 37655 14783 37689
rect 15149 37655 15183 37689
rect 15549 37655 15583 37689
rect 15949 37655 15983 37689
rect 16349 37655 16383 37689
rect 16749 37655 16783 37689
rect 17149 37655 17183 37689
rect 17549 37655 17583 37689
rect 17949 37655 17983 37689
rect 18349 37655 18383 37689
rect 18749 37655 18783 37689
rect 19149 37655 19183 37689
rect 19549 37655 19583 37689
rect 19949 37655 19983 37689
rect 20349 37655 20383 37689
rect 20997 37655 21031 37689
rect 21397 37655 21431 37689
rect 21797 37655 21831 37689
rect 22197 37655 22231 37689
rect 22597 37655 22631 37689
rect 22997 37655 23031 37689
rect 23397 37655 23431 37689
rect 23797 37655 23831 37689
rect 24197 37655 24231 37689
rect 24597 37655 24631 37689
rect 24997 37655 25031 37689
rect 25397 37655 25431 37689
rect 25797 37655 25831 37689
rect 26197 37655 26231 37689
rect 26597 37655 26631 37689
rect 26997 37655 27031 37689
rect 27397 37655 27431 37689
rect 27797 37655 27831 37689
rect 28511 37655 28545 37689
rect 30207 37655 30241 37689
rect 30407 37655 30441 37689
rect 30607 37655 30641 37689
rect 30807 37655 30841 37689
rect 31007 37655 31041 37689
rect 31207 37655 31241 37689
rect 31407 37655 31441 37689
rect 31607 37655 31641 37689
rect 31807 37655 31841 37689
rect 32007 37655 32041 37689
rect 32207 37655 32241 37689
rect 32407 37655 32441 37689
rect 32607 37655 32641 37689
rect 32807 37655 32841 37689
rect 33007 37655 33041 37689
rect 33207 37655 33241 37689
rect 33407 37655 33441 37689
rect 33607 37655 33641 37689
rect 33807 37655 33841 37689
rect 34007 37655 34041 37689
rect 34207 37655 34241 37689
rect 34407 37655 34441 37689
rect 34607 37655 34641 37689
rect 34807 37655 34841 37689
rect 35007 37655 35041 37689
rect 35207 37655 35241 37689
rect 35407 37655 35441 37689
rect 35607 37655 35641 37689
rect 35807 37655 35841 37689
rect 36007 37655 36041 37689
rect 36207 37655 36241 37689
rect 36407 37655 36441 37689
rect 36607 37655 36641 37689
rect 36807 37655 36841 37689
rect 37007 37655 37041 37689
rect 37207 37655 37241 37689
rect 37407 37655 37441 37689
rect 37607 37655 37641 37689
rect 37807 37655 37841 37689
rect 38007 37655 38041 37689
rect 38207 37655 38241 37689
rect 38407 37655 38441 37689
rect 38607 37655 38641 37689
rect 38807 37655 38841 37689
rect 39007 37655 39041 37689
rect 39207 37655 39241 37689
rect 39929 37655 39963 37689
rect 40129 37655 40163 37689
rect 40329 37655 40363 37689
rect 40529 37655 40563 37689
rect 40729 37655 40763 37689
rect 40929 37655 40963 37689
rect 41129 37655 41163 37689
rect 41329 37655 41363 37689
rect 41529 37655 41563 37689
rect 41729 37655 41763 37689
rect 41929 37655 41963 37689
rect 28825 37485 28859 37519
rect 30070 37322 30104 37356
rect 30160 37341 30194 37356
rect 30250 37341 30284 37356
rect 30340 37341 30374 37356
rect 30430 37341 30464 37356
rect 30520 37341 30554 37356
rect 30610 37341 30644 37356
rect 30700 37341 30734 37356
rect 30790 37341 30824 37356
rect 30880 37341 30914 37356
rect 30970 37341 31004 37356
rect 31060 37341 31094 37356
rect 31150 37341 31184 37356
rect 30160 37322 30180 37341
rect 30180 37322 30194 37341
rect 30250 37322 30270 37341
rect 30270 37322 30284 37341
rect 30340 37322 30360 37341
rect 30360 37322 30374 37341
rect 30430 37322 30450 37341
rect 30450 37322 30464 37341
rect 30520 37322 30540 37341
rect 30540 37322 30554 37341
rect 30610 37322 30630 37341
rect 30630 37322 30644 37341
rect 30700 37322 30720 37341
rect 30720 37322 30734 37341
rect 30790 37322 30810 37341
rect 30810 37322 30824 37341
rect 30880 37322 30900 37341
rect 30900 37322 30914 37341
rect 30970 37322 30990 37341
rect 30990 37322 31004 37341
rect 31060 37322 31080 37341
rect 31080 37322 31094 37341
rect 31150 37322 31170 37341
rect 31170 37322 31184 37341
rect 31240 37322 31274 37356
rect 31410 37322 31444 37356
rect 31500 37341 31534 37356
rect 31590 37341 31624 37356
rect 31680 37341 31714 37356
rect 31770 37341 31804 37356
rect 31860 37341 31894 37356
rect 31950 37341 31984 37356
rect 32040 37341 32074 37356
rect 32130 37341 32164 37356
rect 32220 37341 32254 37356
rect 32310 37341 32344 37356
rect 32400 37341 32434 37356
rect 32490 37341 32524 37356
rect 31500 37322 31520 37341
rect 31520 37322 31534 37341
rect 31590 37322 31610 37341
rect 31610 37322 31624 37341
rect 31680 37322 31700 37341
rect 31700 37322 31714 37341
rect 31770 37322 31790 37341
rect 31790 37322 31804 37341
rect 31860 37322 31880 37341
rect 31880 37322 31894 37341
rect 31950 37322 31970 37341
rect 31970 37322 31984 37341
rect 32040 37322 32060 37341
rect 32060 37322 32074 37341
rect 32130 37322 32150 37341
rect 32150 37322 32164 37341
rect 32220 37322 32240 37341
rect 32240 37322 32254 37341
rect 32310 37322 32330 37341
rect 32330 37322 32344 37341
rect 32400 37322 32420 37341
rect 32420 37322 32434 37341
rect 32490 37322 32510 37341
rect 32510 37322 32524 37341
rect 32580 37322 32614 37356
rect 32750 37322 32784 37356
rect 32840 37341 32874 37356
rect 32930 37341 32964 37356
rect 33020 37341 33054 37356
rect 33110 37341 33144 37356
rect 33200 37341 33234 37356
rect 33290 37341 33324 37356
rect 33380 37341 33414 37356
rect 33470 37341 33504 37356
rect 33560 37341 33594 37356
rect 33650 37341 33684 37356
rect 33740 37341 33774 37356
rect 33830 37341 33864 37356
rect 32840 37322 32860 37341
rect 32860 37322 32874 37341
rect 32930 37322 32950 37341
rect 32950 37322 32964 37341
rect 33020 37322 33040 37341
rect 33040 37322 33054 37341
rect 33110 37322 33130 37341
rect 33130 37322 33144 37341
rect 33200 37322 33220 37341
rect 33220 37322 33234 37341
rect 33290 37322 33310 37341
rect 33310 37322 33324 37341
rect 33380 37322 33400 37341
rect 33400 37322 33414 37341
rect 33470 37322 33490 37341
rect 33490 37322 33504 37341
rect 33560 37322 33580 37341
rect 33580 37322 33594 37341
rect 33650 37322 33670 37341
rect 33670 37322 33684 37341
rect 33740 37322 33760 37341
rect 33760 37322 33774 37341
rect 33830 37322 33850 37341
rect 33850 37322 33864 37341
rect 33920 37322 33954 37356
rect 34090 37322 34124 37356
rect 34180 37341 34214 37356
rect 34270 37341 34304 37356
rect 34360 37341 34394 37356
rect 34450 37341 34484 37356
rect 34540 37341 34574 37356
rect 34630 37341 34664 37356
rect 34720 37341 34754 37356
rect 34810 37341 34844 37356
rect 34900 37341 34934 37356
rect 34990 37341 35024 37356
rect 35080 37341 35114 37356
rect 35170 37341 35204 37356
rect 34180 37322 34200 37341
rect 34200 37322 34214 37341
rect 34270 37322 34290 37341
rect 34290 37322 34304 37341
rect 34360 37322 34380 37341
rect 34380 37322 34394 37341
rect 34450 37322 34470 37341
rect 34470 37322 34484 37341
rect 34540 37322 34560 37341
rect 34560 37322 34574 37341
rect 34630 37322 34650 37341
rect 34650 37322 34664 37341
rect 34720 37322 34740 37341
rect 34740 37322 34754 37341
rect 34810 37322 34830 37341
rect 34830 37322 34844 37341
rect 34900 37322 34920 37341
rect 34920 37322 34934 37341
rect 34990 37322 35010 37341
rect 35010 37322 35024 37341
rect 35080 37322 35100 37341
rect 35100 37322 35114 37341
rect 35170 37322 35190 37341
rect 35190 37322 35204 37341
rect 35260 37322 35294 37356
rect 35430 37322 35464 37356
rect 35520 37341 35554 37356
rect 35610 37341 35644 37356
rect 35700 37341 35734 37356
rect 35790 37341 35824 37356
rect 35880 37341 35914 37356
rect 35970 37341 36004 37356
rect 36060 37341 36094 37356
rect 36150 37341 36184 37356
rect 36240 37341 36274 37356
rect 36330 37341 36364 37356
rect 36420 37341 36454 37356
rect 36510 37341 36544 37356
rect 35520 37322 35540 37341
rect 35540 37322 35554 37341
rect 35610 37322 35630 37341
rect 35630 37322 35644 37341
rect 35700 37322 35720 37341
rect 35720 37322 35734 37341
rect 35790 37322 35810 37341
rect 35810 37322 35824 37341
rect 35880 37322 35900 37341
rect 35900 37322 35914 37341
rect 35970 37322 35990 37341
rect 35990 37322 36004 37341
rect 36060 37322 36080 37341
rect 36080 37322 36094 37341
rect 36150 37322 36170 37341
rect 36170 37322 36184 37341
rect 36240 37322 36260 37341
rect 36260 37322 36274 37341
rect 36330 37322 36350 37341
rect 36350 37322 36364 37341
rect 36420 37322 36440 37341
rect 36440 37322 36454 37341
rect 36510 37322 36530 37341
rect 36530 37322 36544 37341
rect 36600 37322 36634 37356
rect 36770 37322 36804 37356
rect 36860 37341 36894 37356
rect 36950 37341 36984 37356
rect 37040 37341 37074 37356
rect 37130 37341 37164 37356
rect 37220 37341 37254 37356
rect 37310 37341 37344 37356
rect 37400 37341 37434 37356
rect 37490 37341 37524 37356
rect 37580 37341 37614 37356
rect 37670 37341 37704 37356
rect 37760 37341 37794 37356
rect 37850 37341 37884 37356
rect 36860 37322 36880 37341
rect 36880 37322 36894 37341
rect 36950 37322 36970 37341
rect 36970 37322 36984 37341
rect 37040 37322 37060 37341
rect 37060 37322 37074 37341
rect 37130 37322 37150 37341
rect 37150 37322 37164 37341
rect 37220 37322 37240 37341
rect 37240 37322 37254 37341
rect 37310 37322 37330 37341
rect 37330 37322 37344 37341
rect 37400 37322 37420 37341
rect 37420 37322 37434 37341
rect 37490 37322 37510 37341
rect 37510 37322 37524 37341
rect 37580 37322 37600 37341
rect 37600 37322 37614 37341
rect 37670 37322 37690 37341
rect 37690 37322 37704 37341
rect 37760 37322 37780 37341
rect 37780 37322 37794 37341
rect 37850 37322 37870 37341
rect 37870 37322 37884 37341
rect 37940 37322 37974 37356
rect 38110 37322 38144 37356
rect 38200 37341 38234 37356
rect 38290 37341 38324 37356
rect 38380 37341 38414 37356
rect 38470 37341 38504 37356
rect 38560 37341 38594 37356
rect 38650 37341 38684 37356
rect 38740 37341 38774 37356
rect 38830 37341 38864 37356
rect 38920 37341 38954 37356
rect 39010 37341 39044 37356
rect 39100 37341 39134 37356
rect 39190 37341 39224 37356
rect 38200 37322 38220 37341
rect 38220 37322 38234 37341
rect 38290 37322 38310 37341
rect 38310 37322 38324 37341
rect 38380 37322 38400 37341
rect 38400 37322 38414 37341
rect 38470 37322 38490 37341
rect 38490 37322 38504 37341
rect 38560 37322 38580 37341
rect 38580 37322 38594 37341
rect 38650 37322 38670 37341
rect 38670 37322 38684 37341
rect 38740 37322 38760 37341
rect 38760 37322 38774 37341
rect 38830 37322 38850 37341
rect 38850 37322 38864 37341
rect 38920 37322 38940 37341
rect 38940 37322 38954 37341
rect 39010 37322 39030 37341
rect 39030 37322 39044 37341
rect 39100 37322 39120 37341
rect 39120 37322 39134 37341
rect 39190 37322 39210 37341
rect 39210 37322 39224 37341
rect 39280 37322 39314 37356
rect 28340 37149 28374 37169
rect 28340 37135 28374 37149
rect 28340 37081 28374 37097
rect 28340 37063 28374 37081
rect 28340 37013 28374 37025
rect 28340 36991 28374 37013
rect 28340 36945 28374 36953
rect 28340 36919 28374 36945
rect 28340 36877 28374 36881
rect 28340 36847 28374 36877
rect 28340 36775 28374 36809
rect 28340 36707 28374 36737
rect 28340 36703 28374 36707
rect 28340 36639 28374 36665
rect 28340 36631 28374 36639
rect 28340 36571 28374 36593
rect 28340 36559 28374 36571
rect 28340 36503 28374 36521
rect 28340 36487 28374 36503
rect 28340 36435 28374 36449
rect 28340 36415 28374 36435
rect 28798 37149 28832 37169
rect 28798 37135 28832 37149
rect 28798 37081 28832 37097
rect 28798 37063 28832 37081
rect 28798 37013 28832 37025
rect 28798 36991 28832 37013
rect 28798 36945 28832 36953
rect 28798 36919 28832 36945
rect 28798 36877 28832 36881
rect 28798 36847 28832 36877
rect 28798 36775 28832 36809
rect 28798 36707 28832 36737
rect 28798 36703 28832 36707
rect 28798 36639 28832 36665
rect 28798 36631 28832 36639
rect 28798 36571 28832 36593
rect 28798 36559 28832 36571
rect 28798 36503 28832 36521
rect 28798 36487 28832 36503
rect 28798 36435 28832 36449
rect 28798 36415 28832 36435
rect 30234 37162 30268 37196
rect 30324 37194 30358 37196
rect 30414 37194 30448 37196
rect 30504 37194 30538 37196
rect 30594 37194 30628 37196
rect 30684 37194 30718 37196
rect 30774 37194 30808 37196
rect 30864 37194 30898 37196
rect 30954 37194 30988 37196
rect 31044 37194 31078 37196
rect 30324 37162 30344 37194
rect 30344 37162 30358 37194
rect 30414 37162 30434 37194
rect 30434 37162 30448 37194
rect 30504 37162 30524 37194
rect 30524 37162 30538 37194
rect 30594 37162 30614 37194
rect 30614 37162 30628 37194
rect 30684 37162 30704 37194
rect 30704 37162 30718 37194
rect 30774 37162 30794 37194
rect 30794 37162 30808 37194
rect 30864 37162 30884 37194
rect 30884 37162 30898 37194
rect 30954 37162 30974 37194
rect 30974 37162 30988 37194
rect 31044 37162 31064 37194
rect 31064 37162 31078 37194
rect 31134 37162 31168 37196
rect 30420 36986 30442 36992
rect 30442 36986 30454 36992
rect 30520 36986 30532 36992
rect 30532 36986 30554 36992
rect 30620 36986 30622 36992
rect 30622 36986 30654 36992
rect 30420 36958 30454 36986
rect 30520 36958 30554 36986
rect 30620 36958 30654 36986
rect 30720 36958 30754 36992
rect 30820 36958 30854 36992
rect 30920 36986 30948 36992
rect 30948 36986 30954 36992
rect 30920 36958 30954 36986
rect 30420 36858 30454 36892
rect 30520 36858 30554 36892
rect 30620 36858 30654 36892
rect 30720 36858 30754 36892
rect 30820 36858 30854 36892
rect 30920 36858 30954 36892
rect 30420 36758 30454 36792
rect 30520 36758 30554 36792
rect 30620 36758 30654 36792
rect 30720 36758 30754 36792
rect 30820 36758 30854 36792
rect 30920 36758 30954 36792
rect 30420 36660 30454 36692
rect 30520 36660 30554 36692
rect 30620 36660 30654 36692
rect 30420 36658 30442 36660
rect 30442 36658 30454 36660
rect 30520 36658 30532 36660
rect 30532 36658 30554 36660
rect 30620 36658 30622 36660
rect 30622 36658 30654 36660
rect 30720 36658 30754 36692
rect 30820 36658 30854 36692
rect 30920 36660 30954 36692
rect 30920 36658 30948 36660
rect 30948 36658 30954 36660
rect 30420 36570 30454 36592
rect 30520 36570 30554 36592
rect 30620 36570 30654 36592
rect 30420 36558 30442 36570
rect 30442 36558 30454 36570
rect 30520 36558 30532 36570
rect 30532 36558 30554 36570
rect 30620 36558 30622 36570
rect 30622 36558 30654 36570
rect 30720 36558 30754 36592
rect 30820 36558 30854 36592
rect 30920 36570 30954 36592
rect 30920 36558 30948 36570
rect 30948 36558 30954 36570
rect 30420 36480 30454 36492
rect 30520 36480 30554 36492
rect 30620 36480 30654 36492
rect 30420 36458 30442 36480
rect 30442 36458 30454 36480
rect 30520 36458 30532 36480
rect 30532 36458 30554 36480
rect 30620 36458 30622 36480
rect 30622 36458 30654 36480
rect 30720 36458 30754 36492
rect 30820 36458 30854 36492
rect 30920 36480 30954 36492
rect 30920 36458 30948 36480
rect 30948 36458 30954 36480
rect 28365 36193 28399 36227
rect 31574 37162 31608 37196
rect 31664 37194 31698 37196
rect 31754 37194 31788 37196
rect 31844 37194 31878 37196
rect 31934 37194 31968 37196
rect 32024 37194 32058 37196
rect 32114 37194 32148 37196
rect 32204 37194 32238 37196
rect 32294 37194 32328 37196
rect 32384 37194 32418 37196
rect 31664 37162 31684 37194
rect 31684 37162 31698 37194
rect 31754 37162 31774 37194
rect 31774 37162 31788 37194
rect 31844 37162 31864 37194
rect 31864 37162 31878 37194
rect 31934 37162 31954 37194
rect 31954 37162 31968 37194
rect 32024 37162 32044 37194
rect 32044 37162 32058 37194
rect 32114 37162 32134 37194
rect 32134 37162 32148 37194
rect 32204 37162 32224 37194
rect 32224 37162 32238 37194
rect 32294 37162 32314 37194
rect 32314 37162 32328 37194
rect 32384 37162 32404 37194
rect 32404 37162 32418 37194
rect 32474 37162 32508 37196
rect 31760 36986 31782 36992
rect 31782 36986 31794 36992
rect 31860 36986 31872 36992
rect 31872 36986 31894 36992
rect 31960 36986 31962 36992
rect 31962 36986 31994 36992
rect 31760 36958 31794 36986
rect 31860 36958 31894 36986
rect 31960 36958 31994 36986
rect 32060 36958 32094 36992
rect 32160 36958 32194 36992
rect 32260 36986 32288 36992
rect 32288 36986 32294 36992
rect 32260 36958 32294 36986
rect 31760 36858 31794 36892
rect 31860 36858 31894 36892
rect 31960 36858 31994 36892
rect 32060 36858 32094 36892
rect 32160 36858 32194 36892
rect 32260 36858 32294 36892
rect 31760 36758 31794 36792
rect 31860 36758 31894 36792
rect 31960 36758 31994 36792
rect 32060 36758 32094 36792
rect 32160 36758 32194 36792
rect 32260 36758 32294 36792
rect 31760 36660 31794 36692
rect 31860 36660 31894 36692
rect 31960 36660 31994 36692
rect 31760 36658 31782 36660
rect 31782 36658 31794 36660
rect 31860 36658 31872 36660
rect 31872 36658 31894 36660
rect 31960 36658 31962 36660
rect 31962 36658 31994 36660
rect 32060 36658 32094 36692
rect 32160 36658 32194 36692
rect 32260 36660 32294 36692
rect 32260 36658 32288 36660
rect 32288 36658 32294 36660
rect 31760 36570 31794 36592
rect 31860 36570 31894 36592
rect 31960 36570 31994 36592
rect 31760 36558 31782 36570
rect 31782 36558 31794 36570
rect 31860 36558 31872 36570
rect 31872 36558 31894 36570
rect 31960 36558 31962 36570
rect 31962 36558 31994 36570
rect 32060 36558 32094 36592
rect 32160 36558 32194 36592
rect 32260 36570 32294 36592
rect 32260 36558 32288 36570
rect 32288 36558 32294 36570
rect 31760 36480 31794 36492
rect 31860 36480 31894 36492
rect 31960 36480 31994 36492
rect 31760 36458 31782 36480
rect 31782 36458 31794 36480
rect 31860 36458 31872 36480
rect 31872 36458 31894 36480
rect 31960 36458 31962 36480
rect 31962 36458 31994 36480
rect 32060 36458 32094 36492
rect 32160 36458 32194 36492
rect 32260 36480 32294 36492
rect 32260 36458 32288 36480
rect 32288 36458 32294 36480
rect 32914 37162 32948 37196
rect 33004 37194 33038 37196
rect 33094 37194 33128 37196
rect 33184 37194 33218 37196
rect 33274 37194 33308 37196
rect 33364 37194 33398 37196
rect 33454 37194 33488 37196
rect 33544 37194 33578 37196
rect 33634 37194 33668 37196
rect 33724 37194 33758 37196
rect 33004 37162 33024 37194
rect 33024 37162 33038 37194
rect 33094 37162 33114 37194
rect 33114 37162 33128 37194
rect 33184 37162 33204 37194
rect 33204 37162 33218 37194
rect 33274 37162 33294 37194
rect 33294 37162 33308 37194
rect 33364 37162 33384 37194
rect 33384 37162 33398 37194
rect 33454 37162 33474 37194
rect 33474 37162 33488 37194
rect 33544 37162 33564 37194
rect 33564 37162 33578 37194
rect 33634 37162 33654 37194
rect 33654 37162 33668 37194
rect 33724 37162 33744 37194
rect 33744 37162 33758 37194
rect 33814 37162 33848 37196
rect 33100 36986 33122 36992
rect 33122 36986 33134 36992
rect 33200 36986 33212 36992
rect 33212 36986 33234 36992
rect 33300 36986 33302 36992
rect 33302 36986 33334 36992
rect 33100 36958 33134 36986
rect 33200 36958 33234 36986
rect 33300 36958 33334 36986
rect 33400 36958 33434 36992
rect 33500 36958 33534 36992
rect 33600 36986 33628 36992
rect 33628 36986 33634 36992
rect 33600 36958 33634 36986
rect 33100 36858 33134 36892
rect 33200 36858 33234 36892
rect 33300 36858 33334 36892
rect 33400 36858 33434 36892
rect 33500 36858 33534 36892
rect 33600 36858 33634 36892
rect 33100 36758 33134 36792
rect 33200 36758 33234 36792
rect 33300 36758 33334 36792
rect 33400 36758 33434 36792
rect 33500 36758 33534 36792
rect 33600 36758 33634 36792
rect 33100 36660 33134 36692
rect 33200 36660 33234 36692
rect 33300 36660 33334 36692
rect 33100 36658 33122 36660
rect 33122 36658 33134 36660
rect 33200 36658 33212 36660
rect 33212 36658 33234 36660
rect 33300 36658 33302 36660
rect 33302 36658 33334 36660
rect 33400 36658 33434 36692
rect 33500 36658 33534 36692
rect 33600 36660 33634 36692
rect 33600 36658 33628 36660
rect 33628 36658 33634 36660
rect 33100 36570 33134 36592
rect 33200 36570 33234 36592
rect 33300 36570 33334 36592
rect 33100 36558 33122 36570
rect 33122 36558 33134 36570
rect 33200 36558 33212 36570
rect 33212 36558 33234 36570
rect 33300 36558 33302 36570
rect 33302 36558 33334 36570
rect 33400 36558 33434 36592
rect 33500 36558 33534 36592
rect 33600 36570 33634 36592
rect 33600 36558 33628 36570
rect 33628 36558 33634 36570
rect 33100 36480 33134 36492
rect 33200 36480 33234 36492
rect 33300 36480 33334 36492
rect 33100 36458 33122 36480
rect 33122 36458 33134 36480
rect 33200 36458 33212 36480
rect 33212 36458 33234 36480
rect 33300 36458 33302 36480
rect 33302 36458 33334 36480
rect 33400 36458 33434 36492
rect 33500 36458 33534 36492
rect 33600 36480 33634 36492
rect 33600 36458 33628 36480
rect 33628 36458 33634 36480
rect 34254 37162 34288 37196
rect 34344 37194 34378 37196
rect 34434 37194 34468 37196
rect 34524 37194 34558 37196
rect 34614 37194 34648 37196
rect 34704 37194 34738 37196
rect 34794 37194 34828 37196
rect 34884 37194 34918 37196
rect 34974 37194 35008 37196
rect 35064 37194 35098 37196
rect 34344 37162 34364 37194
rect 34364 37162 34378 37194
rect 34434 37162 34454 37194
rect 34454 37162 34468 37194
rect 34524 37162 34544 37194
rect 34544 37162 34558 37194
rect 34614 37162 34634 37194
rect 34634 37162 34648 37194
rect 34704 37162 34724 37194
rect 34724 37162 34738 37194
rect 34794 37162 34814 37194
rect 34814 37162 34828 37194
rect 34884 37162 34904 37194
rect 34904 37162 34918 37194
rect 34974 37162 34994 37194
rect 34994 37162 35008 37194
rect 35064 37162 35084 37194
rect 35084 37162 35098 37194
rect 35154 37162 35188 37196
rect 34440 36986 34462 36992
rect 34462 36986 34474 36992
rect 34540 36986 34552 36992
rect 34552 36986 34574 36992
rect 34640 36986 34642 36992
rect 34642 36986 34674 36992
rect 34440 36958 34474 36986
rect 34540 36958 34574 36986
rect 34640 36958 34674 36986
rect 34740 36958 34774 36992
rect 34840 36958 34874 36992
rect 34940 36986 34968 36992
rect 34968 36986 34974 36992
rect 34940 36958 34974 36986
rect 34440 36858 34474 36892
rect 34540 36858 34574 36892
rect 34640 36858 34674 36892
rect 34740 36858 34774 36892
rect 34840 36858 34874 36892
rect 34940 36858 34974 36892
rect 34440 36758 34474 36792
rect 34540 36758 34574 36792
rect 34640 36758 34674 36792
rect 34740 36758 34774 36792
rect 34840 36758 34874 36792
rect 34940 36758 34974 36792
rect 34440 36660 34474 36692
rect 34540 36660 34574 36692
rect 34640 36660 34674 36692
rect 34440 36658 34462 36660
rect 34462 36658 34474 36660
rect 34540 36658 34552 36660
rect 34552 36658 34574 36660
rect 34640 36658 34642 36660
rect 34642 36658 34674 36660
rect 34740 36658 34774 36692
rect 34840 36658 34874 36692
rect 34940 36660 34974 36692
rect 34940 36658 34968 36660
rect 34968 36658 34974 36660
rect 34440 36570 34474 36592
rect 34540 36570 34574 36592
rect 34640 36570 34674 36592
rect 34440 36558 34462 36570
rect 34462 36558 34474 36570
rect 34540 36558 34552 36570
rect 34552 36558 34574 36570
rect 34640 36558 34642 36570
rect 34642 36558 34674 36570
rect 34740 36558 34774 36592
rect 34840 36558 34874 36592
rect 34940 36570 34974 36592
rect 34940 36558 34968 36570
rect 34968 36558 34974 36570
rect 34440 36480 34474 36492
rect 34540 36480 34574 36492
rect 34640 36480 34674 36492
rect 34440 36458 34462 36480
rect 34462 36458 34474 36480
rect 34540 36458 34552 36480
rect 34552 36458 34574 36480
rect 34640 36458 34642 36480
rect 34642 36458 34674 36480
rect 34740 36458 34774 36492
rect 34840 36458 34874 36492
rect 34940 36480 34974 36492
rect 34940 36458 34968 36480
rect 34968 36458 34974 36480
rect 35594 37162 35628 37196
rect 35684 37194 35718 37196
rect 35774 37194 35808 37196
rect 35864 37194 35898 37196
rect 35954 37194 35988 37196
rect 36044 37194 36078 37196
rect 36134 37194 36168 37196
rect 36224 37194 36258 37196
rect 36314 37194 36348 37196
rect 36404 37194 36438 37196
rect 35684 37162 35704 37194
rect 35704 37162 35718 37194
rect 35774 37162 35794 37194
rect 35794 37162 35808 37194
rect 35864 37162 35884 37194
rect 35884 37162 35898 37194
rect 35954 37162 35974 37194
rect 35974 37162 35988 37194
rect 36044 37162 36064 37194
rect 36064 37162 36078 37194
rect 36134 37162 36154 37194
rect 36154 37162 36168 37194
rect 36224 37162 36244 37194
rect 36244 37162 36258 37194
rect 36314 37162 36334 37194
rect 36334 37162 36348 37194
rect 36404 37162 36424 37194
rect 36424 37162 36438 37194
rect 36494 37162 36528 37196
rect 35780 36986 35802 36992
rect 35802 36986 35814 36992
rect 35880 36986 35892 36992
rect 35892 36986 35914 36992
rect 35980 36986 35982 36992
rect 35982 36986 36014 36992
rect 35780 36958 35814 36986
rect 35880 36958 35914 36986
rect 35980 36958 36014 36986
rect 36080 36958 36114 36992
rect 36180 36958 36214 36992
rect 36280 36986 36308 36992
rect 36308 36986 36314 36992
rect 36280 36958 36314 36986
rect 35780 36858 35814 36892
rect 35880 36858 35914 36892
rect 35980 36858 36014 36892
rect 36080 36858 36114 36892
rect 36180 36858 36214 36892
rect 36280 36858 36314 36892
rect 35780 36758 35814 36792
rect 35880 36758 35914 36792
rect 35980 36758 36014 36792
rect 36080 36758 36114 36792
rect 36180 36758 36214 36792
rect 36280 36758 36314 36792
rect 35780 36660 35814 36692
rect 35880 36660 35914 36692
rect 35980 36660 36014 36692
rect 35780 36658 35802 36660
rect 35802 36658 35814 36660
rect 35880 36658 35892 36660
rect 35892 36658 35914 36660
rect 35980 36658 35982 36660
rect 35982 36658 36014 36660
rect 36080 36658 36114 36692
rect 36180 36658 36214 36692
rect 36280 36660 36314 36692
rect 36280 36658 36308 36660
rect 36308 36658 36314 36660
rect 35780 36570 35814 36592
rect 35880 36570 35914 36592
rect 35980 36570 36014 36592
rect 35780 36558 35802 36570
rect 35802 36558 35814 36570
rect 35880 36558 35892 36570
rect 35892 36558 35914 36570
rect 35980 36558 35982 36570
rect 35982 36558 36014 36570
rect 36080 36558 36114 36592
rect 36180 36558 36214 36592
rect 36280 36570 36314 36592
rect 36280 36558 36308 36570
rect 36308 36558 36314 36570
rect 35780 36480 35814 36492
rect 35880 36480 35914 36492
rect 35980 36480 36014 36492
rect 35780 36458 35802 36480
rect 35802 36458 35814 36480
rect 35880 36458 35892 36480
rect 35892 36458 35914 36480
rect 35980 36458 35982 36480
rect 35982 36458 36014 36480
rect 36080 36458 36114 36492
rect 36180 36458 36214 36492
rect 36280 36480 36314 36492
rect 36280 36458 36308 36480
rect 36308 36458 36314 36480
rect 36934 37162 36968 37196
rect 37024 37194 37058 37196
rect 37114 37194 37148 37196
rect 37204 37194 37238 37196
rect 37294 37194 37328 37196
rect 37384 37194 37418 37196
rect 37474 37194 37508 37196
rect 37564 37194 37598 37196
rect 37654 37194 37688 37196
rect 37744 37194 37778 37196
rect 37024 37162 37044 37194
rect 37044 37162 37058 37194
rect 37114 37162 37134 37194
rect 37134 37162 37148 37194
rect 37204 37162 37224 37194
rect 37224 37162 37238 37194
rect 37294 37162 37314 37194
rect 37314 37162 37328 37194
rect 37384 37162 37404 37194
rect 37404 37162 37418 37194
rect 37474 37162 37494 37194
rect 37494 37162 37508 37194
rect 37564 37162 37584 37194
rect 37584 37162 37598 37194
rect 37654 37162 37674 37194
rect 37674 37162 37688 37194
rect 37744 37162 37764 37194
rect 37764 37162 37778 37194
rect 37834 37162 37868 37196
rect 37120 36986 37142 36992
rect 37142 36986 37154 36992
rect 37220 36986 37232 36992
rect 37232 36986 37254 36992
rect 37320 36986 37322 36992
rect 37322 36986 37354 36992
rect 37120 36958 37154 36986
rect 37220 36958 37254 36986
rect 37320 36958 37354 36986
rect 37420 36958 37454 36992
rect 37520 36958 37554 36992
rect 37620 36986 37648 36992
rect 37648 36986 37654 36992
rect 37620 36958 37654 36986
rect 37120 36858 37154 36892
rect 37220 36858 37254 36892
rect 37320 36858 37354 36892
rect 37420 36858 37454 36892
rect 37520 36858 37554 36892
rect 37620 36858 37654 36892
rect 37120 36758 37154 36792
rect 37220 36758 37254 36792
rect 37320 36758 37354 36792
rect 37420 36758 37454 36792
rect 37520 36758 37554 36792
rect 37620 36758 37654 36792
rect 37120 36660 37154 36692
rect 37220 36660 37254 36692
rect 37320 36660 37354 36692
rect 37120 36658 37142 36660
rect 37142 36658 37154 36660
rect 37220 36658 37232 36660
rect 37232 36658 37254 36660
rect 37320 36658 37322 36660
rect 37322 36658 37354 36660
rect 37420 36658 37454 36692
rect 37520 36658 37554 36692
rect 37620 36660 37654 36692
rect 37620 36658 37648 36660
rect 37648 36658 37654 36660
rect 37120 36570 37154 36592
rect 37220 36570 37254 36592
rect 37320 36570 37354 36592
rect 37120 36558 37142 36570
rect 37142 36558 37154 36570
rect 37220 36558 37232 36570
rect 37232 36558 37254 36570
rect 37320 36558 37322 36570
rect 37322 36558 37354 36570
rect 37420 36558 37454 36592
rect 37520 36558 37554 36592
rect 37620 36570 37654 36592
rect 37620 36558 37648 36570
rect 37648 36558 37654 36570
rect 37120 36480 37154 36492
rect 37220 36480 37254 36492
rect 37320 36480 37354 36492
rect 37120 36458 37142 36480
rect 37142 36458 37154 36480
rect 37220 36458 37232 36480
rect 37232 36458 37254 36480
rect 37320 36458 37322 36480
rect 37322 36458 37354 36480
rect 37420 36458 37454 36492
rect 37520 36458 37554 36492
rect 37620 36480 37654 36492
rect 37620 36458 37648 36480
rect 37648 36458 37654 36480
rect 38274 37162 38308 37196
rect 38364 37194 38398 37196
rect 38454 37194 38488 37196
rect 38544 37194 38578 37196
rect 38634 37194 38668 37196
rect 38724 37194 38758 37196
rect 38814 37194 38848 37196
rect 38904 37194 38938 37196
rect 38994 37194 39028 37196
rect 39084 37194 39118 37196
rect 38364 37162 38384 37194
rect 38384 37162 38398 37194
rect 38454 37162 38474 37194
rect 38474 37162 38488 37194
rect 38544 37162 38564 37194
rect 38564 37162 38578 37194
rect 38634 37162 38654 37194
rect 38654 37162 38668 37194
rect 38724 37162 38744 37194
rect 38744 37162 38758 37194
rect 38814 37162 38834 37194
rect 38834 37162 38848 37194
rect 38904 37162 38924 37194
rect 38924 37162 38938 37194
rect 38994 37162 39014 37194
rect 39014 37162 39028 37194
rect 39084 37162 39104 37194
rect 39104 37162 39118 37194
rect 39174 37162 39208 37196
rect 38460 36986 38482 36992
rect 38482 36986 38494 36992
rect 38560 36986 38572 36992
rect 38572 36986 38594 36992
rect 38660 36986 38662 36992
rect 38662 36986 38694 36992
rect 38460 36958 38494 36986
rect 38560 36958 38594 36986
rect 38660 36958 38694 36986
rect 38760 36958 38794 36992
rect 38860 36958 38894 36992
rect 38960 36986 38988 36992
rect 38988 36986 38994 36992
rect 38960 36958 38994 36986
rect 38460 36858 38494 36892
rect 38560 36858 38594 36892
rect 38660 36858 38694 36892
rect 38760 36858 38794 36892
rect 38860 36858 38894 36892
rect 38960 36858 38994 36892
rect 38460 36758 38494 36792
rect 38560 36758 38594 36792
rect 38660 36758 38694 36792
rect 38760 36758 38794 36792
rect 38860 36758 38894 36792
rect 38960 36758 38994 36792
rect 38460 36660 38494 36692
rect 38560 36660 38594 36692
rect 38660 36660 38694 36692
rect 38460 36658 38482 36660
rect 38482 36658 38494 36660
rect 38560 36658 38572 36660
rect 38572 36658 38594 36660
rect 38660 36658 38662 36660
rect 38662 36658 38694 36660
rect 38760 36658 38794 36692
rect 38860 36658 38894 36692
rect 38960 36660 38994 36692
rect 38960 36658 38988 36660
rect 38988 36658 38994 36660
rect 38460 36570 38494 36592
rect 38560 36570 38594 36592
rect 38660 36570 38694 36592
rect 38460 36558 38482 36570
rect 38482 36558 38494 36570
rect 38560 36558 38572 36570
rect 38572 36558 38594 36570
rect 38660 36558 38662 36570
rect 38662 36558 38694 36570
rect 38760 36558 38794 36592
rect 38860 36558 38894 36592
rect 38960 36570 38994 36592
rect 38960 36558 38988 36570
rect 38988 36558 38994 36570
rect 38460 36480 38494 36492
rect 38560 36480 38594 36492
rect 38660 36480 38694 36492
rect 38460 36458 38482 36480
rect 38482 36458 38494 36480
rect 38560 36458 38572 36480
rect 38572 36458 38594 36480
rect 38660 36458 38662 36480
rect 38662 36458 38694 36480
rect 38760 36458 38794 36492
rect 38860 36458 38894 36492
rect 38960 36480 38994 36492
rect 38960 36458 38988 36480
rect 38988 36458 38994 36480
rect 39765 36883 40159 37421
rect 41772 36883 42166 37421
rect 28457 35921 28491 35955
rect 39765 35923 40159 36461
rect 41772 35923 42166 36461
rect 6101 35775 6135 35809
rect 6501 35775 6535 35809
rect 6901 35775 6935 35809
rect 7301 35775 7335 35809
rect 7701 35775 7735 35809
rect 8101 35775 8135 35809
rect 8501 35775 8535 35809
rect 8901 35775 8935 35809
rect 9301 35775 9335 35809
rect 9701 35775 9735 35809
rect 10101 35775 10135 35809
rect 10501 35775 10535 35809
rect 10901 35775 10935 35809
rect 11301 35775 11335 35809
rect 11701 35775 11735 35809
rect 12101 35775 12135 35809
rect 12501 35775 12535 35809
rect 12901 35775 12935 35809
rect 13549 35775 13583 35809
rect 13949 35775 13983 35809
rect 14349 35775 14383 35809
rect 14749 35775 14783 35809
rect 15149 35775 15183 35809
rect 15549 35775 15583 35809
rect 15949 35775 15983 35809
rect 16349 35775 16383 35809
rect 16749 35775 16783 35809
rect 17149 35775 17183 35809
rect 17549 35775 17583 35809
rect 17949 35775 17983 35809
rect 18349 35775 18383 35809
rect 18749 35775 18783 35809
rect 19149 35775 19183 35809
rect 19549 35775 19583 35809
rect 19949 35775 19983 35809
rect 20349 35775 20383 35809
rect 20997 35775 21031 35809
rect 21397 35775 21431 35809
rect 21797 35775 21831 35809
rect 22197 35775 22231 35809
rect 22597 35775 22631 35809
rect 22997 35775 23031 35809
rect 23397 35775 23431 35809
rect 23797 35775 23831 35809
rect 24197 35775 24231 35809
rect 24597 35775 24631 35809
rect 24997 35775 25031 35809
rect 25397 35775 25431 35809
rect 25797 35775 25831 35809
rect 26197 35775 26231 35809
rect 26597 35775 26631 35809
rect 26997 35775 27031 35809
rect 27397 35775 27431 35809
rect 27797 35775 27831 35809
rect 28511 35775 28545 35809
rect 30207 35775 30241 35809
rect 30407 35775 30441 35809
rect 30607 35775 30641 35809
rect 30807 35775 30841 35809
rect 31007 35775 31041 35809
rect 31207 35775 31241 35809
rect 31407 35775 31441 35809
rect 31607 35775 31641 35809
rect 31807 35775 31841 35809
rect 32007 35775 32041 35809
rect 32207 35775 32241 35809
rect 32407 35775 32441 35809
rect 32607 35775 32641 35809
rect 32807 35775 32841 35809
rect 33007 35775 33041 35809
rect 33207 35775 33241 35809
rect 33407 35775 33441 35809
rect 33607 35775 33641 35809
rect 33807 35775 33841 35809
rect 34007 35775 34041 35809
rect 34207 35775 34241 35809
rect 34407 35775 34441 35809
rect 34607 35775 34641 35809
rect 34807 35775 34841 35809
rect 35007 35775 35041 35809
rect 35207 35775 35241 35809
rect 35407 35775 35441 35809
rect 35607 35775 35641 35809
rect 35807 35775 35841 35809
rect 36007 35775 36041 35809
rect 36207 35775 36241 35809
rect 36407 35775 36441 35809
rect 36607 35775 36641 35809
rect 36807 35775 36841 35809
rect 37007 35775 37041 35809
rect 37207 35775 37241 35809
rect 37407 35775 37441 35809
rect 37607 35775 37641 35809
rect 37807 35775 37841 35809
rect 38007 35775 38041 35809
rect 38207 35775 38241 35809
rect 38407 35775 38441 35809
rect 38607 35775 38641 35809
rect 38807 35775 38841 35809
rect 39007 35775 39041 35809
rect 39207 35775 39241 35809
rect 39929 35775 39963 35809
rect 40129 35775 40163 35809
rect 40329 35775 40363 35809
rect 40529 35775 40563 35809
rect 40729 35775 40763 35809
rect 40929 35775 40963 35809
rect 41129 35775 41163 35809
rect 41329 35775 41363 35809
rect 41529 35775 41563 35809
rect 41729 35775 41763 35809
rect 41929 35775 41963 35809
rect 6787 33895 6821 33929
rect 7187 33895 7221 33929
rect 7587 33895 7621 33929
rect 7987 33895 8021 33929
rect 8387 33895 8421 33929
rect 8787 33895 8821 33929
rect 9187 33895 9221 33929
rect 9587 33895 9621 33929
rect 9987 33895 10021 33929
rect 10387 33895 10421 33929
rect 10787 33895 10821 33929
rect 11187 33895 11221 33929
rect 11587 33895 11621 33929
rect 11987 33895 12021 33929
rect 12387 33895 12421 33929
rect 12787 33895 12821 33929
rect 13187 33895 13221 33929
rect 13587 33895 13621 33929
rect 14331 33895 14365 33929
rect 14731 33895 14765 33929
rect 15131 33895 15165 33929
rect 15531 33895 15565 33929
rect 15931 33895 15965 33929
rect 16331 33895 16365 33929
rect 16731 33895 16765 33929
rect 17131 33895 17165 33929
rect 17531 33895 17565 33929
rect 17931 33895 17965 33929
rect 18331 33895 18365 33929
rect 18731 33895 18765 33929
rect 19131 33895 19165 33929
rect 19531 33895 19565 33929
rect 19931 33895 19965 33929
rect 20331 33895 20365 33929
rect 20731 33895 20765 33929
rect 21131 33895 21165 33929
rect 21531 33895 21565 33929
rect 21931 33895 21965 33929
rect 22331 33895 22365 33929
rect 22731 33895 22765 33929
rect 23131 33895 23165 33929
rect 23531 33895 23565 33929
rect 23931 33895 23965 33929
rect 24331 33895 24365 33929
rect 24731 33895 24765 33929
rect 25131 33895 25165 33929
rect 25531 33895 25565 33929
rect 25931 33895 25965 33929
rect 26331 33895 26365 33929
rect 26731 33895 26765 33929
rect 27131 33895 27165 33929
rect 27531 33895 27565 33929
rect 27931 33895 27965 33929
rect 28331 33895 28365 33929
rect 28731 33895 28765 33929
rect 29131 33895 29165 33929
rect 29531 33895 29565 33929
rect 29931 33895 29965 33929
rect 30331 33895 30365 33929
rect 30731 33895 30765 33929
rect 31131 33895 31165 33929
rect 31531 33895 31565 33929
rect 31931 33895 31965 33929
rect 32331 33895 32365 33929
rect 32731 33895 32765 33929
rect 33131 33895 33165 33929
rect 33531 33895 33565 33929
rect 33931 33895 33965 33929
rect 34331 33895 34365 33929
rect 34731 33895 34765 33929
rect 35131 33895 35165 33929
rect 35531 33895 35565 33929
rect 35931 33895 35965 33929
rect 36331 33895 36365 33929
rect 36731 33895 36765 33929
rect 37131 33895 37165 33929
rect 37531 33895 37565 33929
rect 37931 33895 37965 33929
rect 38331 33895 38365 33929
rect 38731 33895 38765 33929
rect 39131 33895 39165 33929
rect 39531 33895 39565 33929
rect 39931 33895 39965 33929
rect 40331 33895 40365 33929
rect 40731 33895 40765 33929
rect 41131 33895 41165 33929
rect 41531 33895 41565 33929
rect 14195 33627 14229 33661
rect 14195 33559 14229 33589
rect 14195 33555 14229 33559
rect 14195 33491 14229 33517
rect 14195 33483 14229 33491
rect 14195 33423 14229 33445
rect 14195 33411 14229 33423
rect 14195 33355 14229 33373
rect 14195 33339 14229 33355
rect 14195 33287 14229 33301
rect 14195 33267 14229 33287
rect 14195 33219 14229 33229
rect 14195 33195 14229 33219
rect 14195 33151 14229 33157
rect 14195 33123 14229 33151
rect 14195 33083 14229 33085
rect 14195 33051 14229 33083
rect 14195 32981 14229 33013
rect 14195 32979 14229 32981
rect 14195 32913 14229 32941
rect 14195 32907 14229 32913
rect 14195 32845 14229 32869
rect 14195 32835 14229 32845
rect 14195 32777 14229 32797
rect 14195 32763 14229 32777
rect 14195 32709 14229 32725
rect 14195 32691 14229 32709
rect 14195 32641 14229 32653
rect 14195 32619 14229 32641
rect 14195 32573 14229 32581
rect 14195 32547 14229 32573
rect 14195 32505 14229 32509
rect 14195 32475 14229 32505
rect 14195 32403 14229 32437
rect 14653 33627 14687 33661
rect 14653 33559 14687 33589
rect 14653 33555 14687 33559
rect 14653 33491 14687 33517
rect 14653 33483 14687 33491
rect 14653 33423 14687 33445
rect 14653 33411 14687 33423
rect 14653 33355 14687 33373
rect 14653 33339 14687 33355
rect 14653 33287 14687 33301
rect 14653 33267 14687 33287
rect 14653 33219 14687 33229
rect 14653 33195 14687 33219
rect 14653 33151 14687 33157
rect 14653 33123 14687 33151
rect 14653 33083 14687 33085
rect 14653 33051 14687 33083
rect 14653 32981 14687 33013
rect 14653 32979 14687 32981
rect 14653 32913 14687 32941
rect 14653 32907 14687 32913
rect 14653 32845 14687 32869
rect 14653 32835 14687 32845
rect 14653 32777 14687 32797
rect 14653 32763 14687 32777
rect 14653 32709 14687 32725
rect 14653 32691 14687 32709
rect 14653 32641 14687 32653
rect 14653 32619 14687 32641
rect 14653 32573 14687 32581
rect 14653 32547 14687 32573
rect 14653 32505 14687 32509
rect 14653 32475 14687 32505
rect 14653 32403 14687 32437
rect 15111 33627 15145 33661
rect 15111 33559 15145 33589
rect 15111 33555 15145 33559
rect 15111 33491 15145 33517
rect 15111 33483 15145 33491
rect 15111 33423 15145 33445
rect 15111 33411 15145 33423
rect 15111 33355 15145 33373
rect 15111 33339 15145 33355
rect 15111 33287 15145 33301
rect 15111 33267 15145 33287
rect 15111 33219 15145 33229
rect 15111 33195 15145 33219
rect 15111 33151 15145 33157
rect 15111 33123 15145 33151
rect 15111 33083 15145 33085
rect 15111 33051 15145 33083
rect 15111 32981 15145 33013
rect 15111 32979 15145 32981
rect 15111 32913 15145 32941
rect 15111 32907 15145 32913
rect 15111 32845 15145 32869
rect 15111 32835 15145 32845
rect 15111 32777 15145 32797
rect 15111 32763 15145 32777
rect 15111 32709 15145 32725
rect 15111 32691 15145 32709
rect 15111 32641 15145 32653
rect 15111 32619 15145 32641
rect 15111 32573 15145 32581
rect 15111 32547 15145 32573
rect 15111 32505 15145 32509
rect 15111 32475 15145 32505
rect 15111 32403 15145 32437
rect 15569 33627 15603 33661
rect 15569 33559 15603 33589
rect 15569 33555 15603 33559
rect 15569 33491 15603 33517
rect 15569 33483 15603 33491
rect 15569 33423 15603 33445
rect 15569 33411 15603 33423
rect 15569 33355 15603 33373
rect 15569 33339 15603 33355
rect 15569 33287 15603 33301
rect 15569 33267 15603 33287
rect 15569 33219 15603 33229
rect 15569 33195 15603 33219
rect 15569 33151 15603 33157
rect 15569 33123 15603 33151
rect 15569 33083 15603 33085
rect 15569 33051 15603 33083
rect 15569 32981 15603 33013
rect 15569 32979 15603 32981
rect 15569 32913 15603 32941
rect 15569 32907 15603 32913
rect 15569 32845 15603 32869
rect 15569 32835 15603 32845
rect 15569 32777 15603 32797
rect 15569 32763 15603 32777
rect 15569 32709 15603 32725
rect 15569 32691 15603 32709
rect 15569 32641 15603 32653
rect 15569 32619 15603 32641
rect 15569 32573 15603 32581
rect 15569 32547 15603 32573
rect 15569 32505 15603 32509
rect 15569 32475 15603 32505
rect 15569 32403 15603 32437
rect 16027 33627 16061 33661
rect 16027 33559 16061 33589
rect 16027 33555 16061 33559
rect 16027 33491 16061 33517
rect 16027 33483 16061 33491
rect 16027 33423 16061 33445
rect 16027 33411 16061 33423
rect 16027 33355 16061 33373
rect 16027 33339 16061 33355
rect 16027 33287 16061 33301
rect 16027 33267 16061 33287
rect 16027 33219 16061 33229
rect 16027 33195 16061 33219
rect 16027 33151 16061 33157
rect 16027 33123 16061 33151
rect 16027 33083 16061 33085
rect 16027 33051 16061 33083
rect 16027 32981 16061 33013
rect 16027 32979 16061 32981
rect 16027 32913 16061 32941
rect 16027 32907 16061 32913
rect 16027 32845 16061 32869
rect 16027 32835 16061 32845
rect 16027 32777 16061 32797
rect 16027 32763 16061 32777
rect 16027 32709 16061 32725
rect 16027 32691 16061 32709
rect 16027 32641 16061 32653
rect 16027 32619 16061 32641
rect 16027 32573 16061 32581
rect 16027 32547 16061 32573
rect 16027 32505 16061 32509
rect 16027 32475 16061 32505
rect 16027 32403 16061 32437
rect 16485 33627 16519 33661
rect 16485 33559 16519 33589
rect 16485 33555 16519 33559
rect 16485 33491 16519 33517
rect 16485 33483 16519 33491
rect 16485 33423 16519 33445
rect 16485 33411 16519 33423
rect 16485 33355 16519 33373
rect 16485 33339 16519 33355
rect 16485 33287 16519 33301
rect 16485 33267 16519 33287
rect 16485 33219 16519 33229
rect 16485 33195 16519 33219
rect 16485 33151 16519 33157
rect 16485 33123 16519 33151
rect 16485 33083 16519 33085
rect 16485 33051 16519 33083
rect 16485 32981 16519 33013
rect 16485 32979 16519 32981
rect 16485 32913 16519 32941
rect 16485 32907 16519 32913
rect 16485 32845 16519 32869
rect 16485 32835 16519 32845
rect 16485 32777 16519 32797
rect 16485 32763 16519 32777
rect 16485 32709 16519 32725
rect 16485 32691 16519 32709
rect 16485 32641 16519 32653
rect 16485 32619 16519 32641
rect 16485 32573 16519 32581
rect 16485 32547 16519 32573
rect 16485 32505 16519 32509
rect 16485 32475 16519 32505
rect 16485 32403 16519 32437
rect 16943 33627 16977 33661
rect 16943 33559 16977 33589
rect 16943 33555 16977 33559
rect 16943 33491 16977 33517
rect 16943 33483 16977 33491
rect 16943 33423 16977 33445
rect 16943 33411 16977 33423
rect 16943 33355 16977 33373
rect 16943 33339 16977 33355
rect 16943 33287 16977 33301
rect 16943 33267 16977 33287
rect 16943 33219 16977 33229
rect 16943 33195 16977 33219
rect 16943 33151 16977 33157
rect 16943 33123 16977 33151
rect 16943 33083 16977 33085
rect 16943 33051 16977 33083
rect 16943 32981 16977 33013
rect 16943 32979 16977 32981
rect 16943 32913 16977 32941
rect 16943 32907 16977 32913
rect 16943 32845 16977 32869
rect 16943 32835 16977 32845
rect 16943 32777 16977 32797
rect 16943 32763 16977 32777
rect 16943 32709 16977 32725
rect 16943 32691 16977 32709
rect 16943 32641 16977 32653
rect 16943 32619 16977 32641
rect 16943 32573 16977 32581
rect 16943 32547 16977 32573
rect 16943 32505 16977 32509
rect 16943 32475 16977 32505
rect 16943 32403 16977 32437
rect 17401 33627 17435 33661
rect 17401 33559 17435 33589
rect 17401 33555 17435 33559
rect 17401 33491 17435 33517
rect 17401 33483 17435 33491
rect 17401 33423 17435 33445
rect 17401 33411 17435 33423
rect 17401 33355 17435 33373
rect 17401 33339 17435 33355
rect 17401 33287 17435 33301
rect 17401 33267 17435 33287
rect 17401 33219 17435 33229
rect 17401 33195 17435 33219
rect 17401 33151 17435 33157
rect 17401 33123 17435 33151
rect 17401 33083 17435 33085
rect 17401 33051 17435 33083
rect 17401 32981 17435 33013
rect 17401 32979 17435 32981
rect 17401 32913 17435 32941
rect 17401 32907 17435 32913
rect 17401 32845 17435 32869
rect 17401 32835 17435 32845
rect 17401 32777 17435 32797
rect 17401 32763 17435 32777
rect 17401 32709 17435 32725
rect 17401 32691 17435 32709
rect 17401 32641 17435 32653
rect 17401 32619 17435 32641
rect 17401 32573 17435 32581
rect 17401 32547 17435 32573
rect 17401 32505 17435 32509
rect 17401 32475 17435 32505
rect 17401 32403 17435 32437
rect 17859 33627 17893 33661
rect 17859 33559 17893 33589
rect 17859 33555 17893 33559
rect 17859 33491 17893 33517
rect 17859 33483 17893 33491
rect 17859 33423 17893 33445
rect 17859 33411 17893 33423
rect 17859 33355 17893 33373
rect 17859 33339 17893 33355
rect 17859 33287 17893 33301
rect 17859 33267 17893 33287
rect 17859 33219 17893 33229
rect 17859 33195 17893 33219
rect 17859 33151 17893 33157
rect 17859 33123 17893 33151
rect 17859 33083 17893 33085
rect 17859 33051 17893 33083
rect 17859 32981 17893 33013
rect 17859 32979 17893 32981
rect 17859 32913 17893 32941
rect 17859 32907 17893 32913
rect 17859 32845 17893 32869
rect 17859 32835 17893 32845
rect 17859 32777 17893 32797
rect 17859 32763 17893 32777
rect 17859 32709 17893 32725
rect 17859 32691 17893 32709
rect 17859 32641 17893 32653
rect 17859 32619 17893 32641
rect 17859 32573 17893 32581
rect 17859 32547 17893 32573
rect 17859 32505 17893 32509
rect 17859 32475 17893 32505
rect 17859 32403 17893 32437
rect 18317 33627 18351 33661
rect 18317 33559 18351 33589
rect 18317 33555 18351 33559
rect 18317 33491 18351 33517
rect 18317 33483 18351 33491
rect 18317 33423 18351 33445
rect 18317 33411 18351 33423
rect 18317 33355 18351 33373
rect 18317 33339 18351 33355
rect 18317 33287 18351 33301
rect 18317 33267 18351 33287
rect 18317 33219 18351 33229
rect 18317 33195 18351 33219
rect 18317 33151 18351 33157
rect 18317 33123 18351 33151
rect 18317 33083 18351 33085
rect 18317 33051 18351 33083
rect 18317 32981 18351 33013
rect 18317 32979 18351 32981
rect 18317 32913 18351 32941
rect 18317 32907 18351 32913
rect 18317 32845 18351 32869
rect 18317 32835 18351 32845
rect 18317 32777 18351 32797
rect 18317 32763 18351 32777
rect 18317 32709 18351 32725
rect 18317 32691 18351 32709
rect 18317 32641 18351 32653
rect 18317 32619 18351 32641
rect 18317 32573 18351 32581
rect 18317 32547 18351 32573
rect 18317 32505 18351 32509
rect 18317 32475 18351 32505
rect 18317 32403 18351 32437
rect 18775 33627 18809 33661
rect 18775 33559 18809 33589
rect 18775 33555 18809 33559
rect 18775 33491 18809 33517
rect 18775 33483 18809 33491
rect 18775 33423 18809 33445
rect 18775 33411 18809 33423
rect 18775 33355 18809 33373
rect 18775 33339 18809 33355
rect 18775 33287 18809 33301
rect 18775 33267 18809 33287
rect 18775 33219 18809 33229
rect 18775 33195 18809 33219
rect 18775 33151 18809 33157
rect 18775 33123 18809 33151
rect 18775 33083 18809 33085
rect 18775 33051 18809 33083
rect 18775 32981 18809 33013
rect 18775 32979 18809 32981
rect 18775 32913 18809 32941
rect 18775 32907 18809 32913
rect 18775 32845 18809 32869
rect 18775 32835 18809 32845
rect 18775 32777 18809 32797
rect 18775 32763 18809 32777
rect 18775 32709 18809 32725
rect 18775 32691 18809 32709
rect 18775 32641 18809 32653
rect 18775 32619 18809 32641
rect 18775 32573 18809 32581
rect 18775 32547 18809 32573
rect 18775 32505 18809 32509
rect 18775 32475 18809 32505
rect 18775 32403 18809 32437
rect 19233 33627 19267 33661
rect 19233 33559 19267 33589
rect 19233 33555 19267 33559
rect 19233 33491 19267 33517
rect 19233 33483 19267 33491
rect 19233 33423 19267 33445
rect 19233 33411 19267 33423
rect 19233 33355 19267 33373
rect 19233 33339 19267 33355
rect 19233 33287 19267 33301
rect 19233 33267 19267 33287
rect 19233 33219 19267 33229
rect 19233 33195 19267 33219
rect 19233 33151 19267 33157
rect 19233 33123 19267 33151
rect 19233 33083 19267 33085
rect 19233 33051 19267 33083
rect 19233 32981 19267 33013
rect 19233 32979 19267 32981
rect 19233 32913 19267 32941
rect 19233 32907 19267 32913
rect 19233 32845 19267 32869
rect 19233 32835 19267 32845
rect 19233 32777 19267 32797
rect 19233 32763 19267 32777
rect 19233 32709 19267 32725
rect 19233 32691 19267 32709
rect 19233 32641 19267 32653
rect 19233 32619 19267 32641
rect 19233 32573 19267 32581
rect 19233 32547 19267 32573
rect 19233 32505 19267 32509
rect 19233 32475 19267 32505
rect 19233 32403 19267 32437
rect 19691 33627 19725 33661
rect 19691 33559 19725 33589
rect 19691 33555 19725 33559
rect 19691 33491 19725 33517
rect 19691 33483 19725 33491
rect 19691 33423 19725 33445
rect 19691 33411 19725 33423
rect 19691 33355 19725 33373
rect 19691 33339 19725 33355
rect 19691 33287 19725 33301
rect 19691 33267 19725 33287
rect 19691 33219 19725 33229
rect 19691 33195 19725 33219
rect 19691 33151 19725 33157
rect 19691 33123 19725 33151
rect 19691 33083 19725 33085
rect 19691 33051 19725 33083
rect 19691 32981 19725 33013
rect 19691 32979 19725 32981
rect 19691 32913 19725 32941
rect 19691 32907 19725 32913
rect 19691 32845 19725 32869
rect 19691 32835 19725 32845
rect 19691 32777 19725 32797
rect 19691 32763 19725 32777
rect 19691 32709 19725 32725
rect 19691 32691 19725 32709
rect 19691 32641 19725 32653
rect 19691 32619 19725 32641
rect 19691 32573 19725 32581
rect 19691 32547 19725 32573
rect 19691 32505 19725 32509
rect 19691 32475 19725 32505
rect 19691 32403 19725 32437
rect 20149 33627 20183 33661
rect 20149 33559 20183 33589
rect 20149 33555 20183 33559
rect 20149 33491 20183 33517
rect 20149 33483 20183 33491
rect 20149 33423 20183 33445
rect 20149 33411 20183 33423
rect 20149 33355 20183 33373
rect 20149 33339 20183 33355
rect 20149 33287 20183 33301
rect 20149 33267 20183 33287
rect 20149 33219 20183 33229
rect 20149 33195 20183 33219
rect 20149 33151 20183 33157
rect 20149 33123 20183 33151
rect 20149 33083 20183 33085
rect 20149 33051 20183 33083
rect 20149 32981 20183 33013
rect 20149 32979 20183 32981
rect 20149 32913 20183 32941
rect 20149 32907 20183 32913
rect 20149 32845 20183 32869
rect 20149 32835 20183 32845
rect 20149 32777 20183 32797
rect 20149 32763 20183 32777
rect 20149 32709 20183 32725
rect 20149 32691 20183 32709
rect 20149 32641 20183 32653
rect 20149 32619 20183 32641
rect 20149 32573 20183 32581
rect 20149 32547 20183 32573
rect 20149 32505 20183 32509
rect 20149 32475 20183 32505
rect 20149 32403 20183 32437
rect 20607 33627 20641 33661
rect 20607 33559 20641 33589
rect 20607 33555 20641 33559
rect 20607 33491 20641 33517
rect 20607 33483 20641 33491
rect 20607 33423 20641 33445
rect 20607 33411 20641 33423
rect 20607 33355 20641 33373
rect 20607 33339 20641 33355
rect 20607 33287 20641 33301
rect 20607 33267 20641 33287
rect 20607 33219 20641 33229
rect 20607 33195 20641 33219
rect 20607 33151 20641 33157
rect 20607 33123 20641 33151
rect 20607 33083 20641 33085
rect 20607 33051 20641 33083
rect 20607 32981 20641 33013
rect 20607 32979 20641 32981
rect 20607 32913 20641 32941
rect 20607 32907 20641 32913
rect 20607 32845 20641 32869
rect 20607 32835 20641 32845
rect 20607 32777 20641 32797
rect 20607 32763 20641 32777
rect 20607 32709 20641 32725
rect 20607 32691 20641 32709
rect 20607 32641 20641 32653
rect 20607 32619 20641 32641
rect 20607 32573 20641 32581
rect 20607 32547 20641 32573
rect 20607 32505 20641 32509
rect 20607 32475 20641 32505
rect 20607 32403 20641 32437
rect 21065 33627 21099 33661
rect 21065 33559 21099 33589
rect 21065 33555 21099 33559
rect 21065 33491 21099 33517
rect 21065 33483 21099 33491
rect 21065 33423 21099 33445
rect 21065 33411 21099 33423
rect 21065 33355 21099 33373
rect 21065 33339 21099 33355
rect 21065 33287 21099 33301
rect 21065 33267 21099 33287
rect 21065 33219 21099 33229
rect 21065 33195 21099 33219
rect 21065 33151 21099 33157
rect 21065 33123 21099 33151
rect 21065 33083 21099 33085
rect 21065 33051 21099 33083
rect 21065 32981 21099 33013
rect 21065 32979 21099 32981
rect 21065 32913 21099 32941
rect 21065 32907 21099 32913
rect 21065 32845 21099 32869
rect 21065 32835 21099 32845
rect 21065 32777 21099 32797
rect 21065 32763 21099 32777
rect 21065 32709 21099 32725
rect 21065 32691 21099 32709
rect 21065 32641 21099 32653
rect 21065 32619 21099 32641
rect 21065 32573 21099 32581
rect 21065 32547 21099 32573
rect 21065 32505 21099 32509
rect 21065 32475 21099 32505
rect 21065 32403 21099 32437
rect 21523 33627 21557 33661
rect 21523 33559 21557 33589
rect 21523 33555 21557 33559
rect 21523 33491 21557 33517
rect 21523 33483 21557 33491
rect 21523 33423 21557 33445
rect 21523 33411 21557 33423
rect 21523 33355 21557 33373
rect 21523 33339 21557 33355
rect 21523 33287 21557 33301
rect 21523 33267 21557 33287
rect 21523 33219 21557 33229
rect 21523 33195 21557 33219
rect 21523 33151 21557 33157
rect 21523 33123 21557 33151
rect 21523 33083 21557 33085
rect 21523 33051 21557 33083
rect 21523 32981 21557 33013
rect 21523 32979 21557 32981
rect 21523 32913 21557 32941
rect 21523 32907 21557 32913
rect 21523 32845 21557 32869
rect 21523 32835 21557 32845
rect 21523 32777 21557 32797
rect 21523 32763 21557 32777
rect 21523 32709 21557 32725
rect 21523 32691 21557 32709
rect 21523 32641 21557 32653
rect 21523 32619 21557 32641
rect 21523 32573 21557 32581
rect 21523 32547 21557 32573
rect 21523 32505 21557 32509
rect 21523 32475 21557 32505
rect 21523 32403 21557 32437
rect 21981 33627 22015 33661
rect 21981 33559 22015 33589
rect 21981 33555 22015 33559
rect 21981 33491 22015 33517
rect 21981 33483 22015 33491
rect 21981 33423 22015 33445
rect 21981 33411 22015 33423
rect 21981 33355 22015 33373
rect 21981 33339 22015 33355
rect 21981 33287 22015 33301
rect 21981 33267 22015 33287
rect 21981 33219 22015 33229
rect 21981 33195 22015 33219
rect 21981 33151 22015 33157
rect 21981 33123 22015 33151
rect 21981 33083 22015 33085
rect 21981 33051 22015 33083
rect 21981 32981 22015 33013
rect 21981 32979 22015 32981
rect 21981 32913 22015 32941
rect 21981 32907 22015 32913
rect 21981 32845 22015 32869
rect 21981 32835 22015 32845
rect 21981 32777 22015 32797
rect 21981 32763 22015 32777
rect 21981 32709 22015 32725
rect 21981 32691 22015 32709
rect 21981 32641 22015 32653
rect 21981 32619 22015 32641
rect 21981 32573 22015 32581
rect 21981 32547 22015 32573
rect 21981 32505 22015 32509
rect 21981 32475 22015 32505
rect 21981 32403 22015 32437
rect 22439 33627 22473 33661
rect 22439 33559 22473 33589
rect 22439 33555 22473 33559
rect 22439 33491 22473 33517
rect 22439 33483 22473 33491
rect 22439 33423 22473 33445
rect 22439 33411 22473 33423
rect 22439 33355 22473 33373
rect 22439 33339 22473 33355
rect 22439 33287 22473 33301
rect 22439 33267 22473 33287
rect 22439 33219 22473 33229
rect 22439 33195 22473 33219
rect 22439 33151 22473 33157
rect 22439 33123 22473 33151
rect 22439 33083 22473 33085
rect 22439 33051 22473 33083
rect 22439 32981 22473 33013
rect 22439 32979 22473 32981
rect 22439 32913 22473 32941
rect 22439 32907 22473 32913
rect 22439 32845 22473 32869
rect 22439 32835 22473 32845
rect 22439 32777 22473 32797
rect 22439 32763 22473 32777
rect 22439 32709 22473 32725
rect 22439 32691 22473 32709
rect 22439 32641 22473 32653
rect 22439 32619 22473 32641
rect 22439 32573 22473 32581
rect 22439 32547 22473 32573
rect 22439 32505 22473 32509
rect 22439 32475 22473 32505
rect 22439 32403 22473 32437
rect 22897 33627 22931 33661
rect 22897 33559 22931 33589
rect 22897 33555 22931 33559
rect 22897 33491 22931 33517
rect 22897 33483 22931 33491
rect 22897 33423 22931 33445
rect 22897 33411 22931 33423
rect 22897 33355 22931 33373
rect 22897 33339 22931 33355
rect 22897 33287 22931 33301
rect 22897 33267 22931 33287
rect 22897 33219 22931 33229
rect 22897 33195 22931 33219
rect 22897 33151 22931 33157
rect 22897 33123 22931 33151
rect 22897 33083 22931 33085
rect 22897 33051 22931 33083
rect 22897 32981 22931 33013
rect 22897 32979 22931 32981
rect 22897 32913 22931 32941
rect 22897 32907 22931 32913
rect 22897 32845 22931 32869
rect 22897 32835 22931 32845
rect 22897 32777 22931 32797
rect 22897 32763 22931 32777
rect 22897 32709 22931 32725
rect 22897 32691 22931 32709
rect 22897 32641 22931 32653
rect 22897 32619 22931 32641
rect 22897 32573 22931 32581
rect 22897 32547 22931 32573
rect 22897 32505 22931 32509
rect 22897 32475 22931 32505
rect 22897 32403 22931 32437
rect 23355 33627 23389 33661
rect 23355 33559 23389 33589
rect 23355 33555 23389 33559
rect 23355 33491 23389 33517
rect 23355 33483 23389 33491
rect 23355 33423 23389 33445
rect 23355 33411 23389 33423
rect 23355 33355 23389 33373
rect 23355 33339 23389 33355
rect 23355 33287 23389 33301
rect 23355 33267 23389 33287
rect 23355 33219 23389 33229
rect 23355 33195 23389 33219
rect 23355 33151 23389 33157
rect 23355 33123 23389 33151
rect 23355 33083 23389 33085
rect 23355 33051 23389 33083
rect 23355 32981 23389 33013
rect 23355 32979 23389 32981
rect 23355 32913 23389 32941
rect 23355 32907 23389 32913
rect 23355 32845 23389 32869
rect 23355 32835 23389 32845
rect 23355 32777 23389 32797
rect 23355 32763 23389 32777
rect 23355 32709 23389 32725
rect 23355 32691 23389 32709
rect 23355 32641 23389 32653
rect 23355 32619 23389 32641
rect 23355 32573 23389 32581
rect 23355 32547 23389 32573
rect 23355 32505 23389 32509
rect 23355 32475 23389 32505
rect 23355 32403 23389 32437
rect 23813 33627 23847 33661
rect 23813 33559 23847 33589
rect 23813 33555 23847 33559
rect 23813 33491 23847 33517
rect 23813 33483 23847 33491
rect 23813 33423 23847 33445
rect 23813 33411 23847 33423
rect 23813 33355 23847 33373
rect 23813 33339 23847 33355
rect 23813 33287 23847 33301
rect 23813 33267 23847 33287
rect 23813 33219 23847 33229
rect 23813 33195 23847 33219
rect 23813 33151 23847 33157
rect 23813 33123 23847 33151
rect 23813 33083 23847 33085
rect 23813 33051 23847 33083
rect 23813 32981 23847 33013
rect 23813 32979 23847 32981
rect 23813 32913 23847 32941
rect 23813 32907 23847 32913
rect 23813 32845 23847 32869
rect 23813 32835 23847 32845
rect 23813 32777 23847 32797
rect 23813 32763 23847 32777
rect 23813 32709 23847 32725
rect 23813 32691 23847 32709
rect 23813 32641 23847 32653
rect 23813 32619 23847 32641
rect 23813 32573 23847 32581
rect 23813 32547 23847 32573
rect 23813 32505 23847 32509
rect 23813 32475 23847 32505
rect 23813 32403 23847 32437
rect 24271 33627 24305 33661
rect 24271 33559 24305 33589
rect 24271 33555 24305 33559
rect 24271 33491 24305 33517
rect 24271 33483 24305 33491
rect 24271 33423 24305 33445
rect 24271 33411 24305 33423
rect 24271 33355 24305 33373
rect 24271 33339 24305 33355
rect 24271 33287 24305 33301
rect 24271 33267 24305 33287
rect 24271 33219 24305 33229
rect 24271 33195 24305 33219
rect 24271 33151 24305 33157
rect 24271 33123 24305 33151
rect 24271 33083 24305 33085
rect 24271 33051 24305 33083
rect 24271 32981 24305 33013
rect 24271 32979 24305 32981
rect 24271 32913 24305 32941
rect 24271 32907 24305 32913
rect 24271 32845 24305 32869
rect 24271 32835 24305 32845
rect 24271 32777 24305 32797
rect 24271 32763 24305 32777
rect 24271 32709 24305 32725
rect 24271 32691 24305 32709
rect 24271 32641 24305 32653
rect 24271 32619 24305 32641
rect 24271 32573 24305 32581
rect 24271 32547 24305 32573
rect 24271 32505 24305 32509
rect 24271 32475 24305 32505
rect 24271 32403 24305 32437
rect 24729 33627 24763 33661
rect 24729 33559 24763 33589
rect 24729 33555 24763 33559
rect 24729 33491 24763 33517
rect 24729 33483 24763 33491
rect 24729 33423 24763 33445
rect 24729 33411 24763 33423
rect 24729 33355 24763 33373
rect 24729 33339 24763 33355
rect 24729 33287 24763 33301
rect 24729 33267 24763 33287
rect 24729 33219 24763 33229
rect 24729 33195 24763 33219
rect 24729 33151 24763 33157
rect 24729 33123 24763 33151
rect 24729 33083 24763 33085
rect 24729 33051 24763 33083
rect 24729 32981 24763 33013
rect 24729 32979 24763 32981
rect 24729 32913 24763 32941
rect 24729 32907 24763 32913
rect 24729 32845 24763 32869
rect 24729 32835 24763 32845
rect 24729 32777 24763 32797
rect 24729 32763 24763 32777
rect 24729 32709 24763 32725
rect 24729 32691 24763 32709
rect 24729 32641 24763 32653
rect 24729 32619 24763 32641
rect 24729 32573 24763 32581
rect 24729 32547 24763 32573
rect 24729 32505 24763 32509
rect 24729 32475 24763 32505
rect 24729 32403 24763 32437
rect 25187 33627 25221 33661
rect 25187 33559 25221 33589
rect 25187 33555 25221 33559
rect 25187 33491 25221 33517
rect 25187 33483 25221 33491
rect 25187 33423 25221 33445
rect 25187 33411 25221 33423
rect 25187 33355 25221 33373
rect 25187 33339 25221 33355
rect 25187 33287 25221 33301
rect 25187 33267 25221 33287
rect 25187 33219 25221 33229
rect 25187 33195 25221 33219
rect 25187 33151 25221 33157
rect 25187 33123 25221 33151
rect 25187 33083 25221 33085
rect 25187 33051 25221 33083
rect 25187 32981 25221 33013
rect 25187 32979 25221 32981
rect 25187 32913 25221 32941
rect 25187 32907 25221 32913
rect 25187 32845 25221 32869
rect 25187 32835 25221 32845
rect 25187 32777 25221 32797
rect 25187 32763 25221 32777
rect 25187 32709 25221 32725
rect 25187 32691 25221 32709
rect 25187 32641 25221 32653
rect 25187 32619 25221 32641
rect 25187 32573 25221 32581
rect 25187 32547 25221 32573
rect 25187 32505 25221 32509
rect 25187 32475 25221 32505
rect 25187 32403 25221 32437
rect 25645 33627 25679 33661
rect 25645 33559 25679 33589
rect 25645 33555 25679 33559
rect 25645 33491 25679 33517
rect 25645 33483 25679 33491
rect 25645 33423 25679 33445
rect 25645 33411 25679 33423
rect 25645 33355 25679 33373
rect 25645 33339 25679 33355
rect 25645 33287 25679 33301
rect 25645 33267 25679 33287
rect 25645 33219 25679 33229
rect 25645 33195 25679 33219
rect 25645 33151 25679 33157
rect 25645 33123 25679 33151
rect 25645 33083 25679 33085
rect 25645 33051 25679 33083
rect 25645 32981 25679 33013
rect 25645 32979 25679 32981
rect 25645 32913 25679 32941
rect 25645 32907 25679 32913
rect 25645 32845 25679 32869
rect 25645 32835 25679 32845
rect 25645 32777 25679 32797
rect 25645 32763 25679 32777
rect 25645 32709 25679 32725
rect 25645 32691 25679 32709
rect 25645 32641 25679 32653
rect 25645 32619 25679 32641
rect 25645 32573 25679 32581
rect 25645 32547 25679 32573
rect 25645 32505 25679 32509
rect 25645 32475 25679 32505
rect 25645 32403 25679 32437
rect 26103 33627 26137 33661
rect 26103 33559 26137 33589
rect 26103 33555 26137 33559
rect 26103 33491 26137 33517
rect 26103 33483 26137 33491
rect 26103 33423 26137 33445
rect 26103 33411 26137 33423
rect 26103 33355 26137 33373
rect 26103 33339 26137 33355
rect 26103 33287 26137 33301
rect 26103 33267 26137 33287
rect 26103 33219 26137 33229
rect 26103 33195 26137 33219
rect 26103 33151 26137 33157
rect 26103 33123 26137 33151
rect 26103 33083 26137 33085
rect 26103 33051 26137 33083
rect 26103 32981 26137 33013
rect 26103 32979 26137 32981
rect 26103 32913 26137 32941
rect 26103 32907 26137 32913
rect 26103 32845 26137 32869
rect 26103 32835 26137 32845
rect 26103 32777 26137 32797
rect 26103 32763 26137 32777
rect 26103 32709 26137 32725
rect 26103 32691 26137 32709
rect 26103 32641 26137 32653
rect 26103 32619 26137 32641
rect 26103 32573 26137 32581
rect 26103 32547 26137 32573
rect 26103 32505 26137 32509
rect 26103 32475 26137 32505
rect 26103 32403 26137 32437
rect 26561 33627 26595 33661
rect 26561 33559 26595 33589
rect 26561 33555 26595 33559
rect 26561 33491 26595 33517
rect 26561 33483 26595 33491
rect 26561 33423 26595 33445
rect 26561 33411 26595 33423
rect 26561 33355 26595 33373
rect 26561 33339 26595 33355
rect 26561 33287 26595 33301
rect 26561 33267 26595 33287
rect 26561 33219 26595 33229
rect 26561 33195 26595 33219
rect 26561 33151 26595 33157
rect 26561 33123 26595 33151
rect 26561 33083 26595 33085
rect 26561 33051 26595 33083
rect 26561 32981 26595 33013
rect 26561 32979 26595 32981
rect 26561 32913 26595 32941
rect 26561 32907 26595 32913
rect 26561 32845 26595 32869
rect 26561 32835 26595 32845
rect 26561 32777 26595 32797
rect 26561 32763 26595 32777
rect 26561 32709 26595 32725
rect 26561 32691 26595 32709
rect 26561 32641 26595 32653
rect 26561 32619 26595 32641
rect 26561 32573 26595 32581
rect 26561 32547 26595 32573
rect 26561 32505 26595 32509
rect 26561 32475 26595 32505
rect 26561 32403 26595 32437
rect 27019 33627 27053 33661
rect 27019 33559 27053 33589
rect 27019 33555 27053 33559
rect 27019 33491 27053 33517
rect 27019 33483 27053 33491
rect 27019 33423 27053 33445
rect 27019 33411 27053 33423
rect 27019 33355 27053 33373
rect 27019 33339 27053 33355
rect 27019 33287 27053 33301
rect 27019 33267 27053 33287
rect 27019 33219 27053 33229
rect 27019 33195 27053 33219
rect 27019 33151 27053 33157
rect 27019 33123 27053 33151
rect 27019 33083 27053 33085
rect 27019 33051 27053 33083
rect 27019 32981 27053 33013
rect 27019 32979 27053 32981
rect 27019 32913 27053 32941
rect 27019 32907 27053 32913
rect 27019 32845 27053 32869
rect 27019 32835 27053 32845
rect 27019 32777 27053 32797
rect 27019 32763 27053 32777
rect 27019 32709 27053 32725
rect 27019 32691 27053 32709
rect 27019 32641 27053 32653
rect 27019 32619 27053 32641
rect 27019 32573 27053 32581
rect 27019 32547 27053 32573
rect 27019 32505 27053 32509
rect 27019 32475 27053 32505
rect 27019 32403 27053 32437
rect 27477 33627 27511 33661
rect 27477 33559 27511 33589
rect 27477 33555 27511 33559
rect 27477 33491 27511 33517
rect 27477 33483 27511 33491
rect 27477 33423 27511 33445
rect 27477 33411 27511 33423
rect 27477 33355 27511 33373
rect 27477 33339 27511 33355
rect 27477 33287 27511 33301
rect 27477 33267 27511 33287
rect 27477 33219 27511 33229
rect 27477 33195 27511 33219
rect 27477 33151 27511 33157
rect 27477 33123 27511 33151
rect 27477 33083 27511 33085
rect 27477 33051 27511 33083
rect 27477 32981 27511 33013
rect 27477 32979 27511 32981
rect 27477 32913 27511 32941
rect 27477 32907 27511 32913
rect 27477 32845 27511 32869
rect 27477 32835 27511 32845
rect 27477 32777 27511 32797
rect 27477 32763 27511 32777
rect 27477 32709 27511 32725
rect 27477 32691 27511 32709
rect 27477 32641 27511 32653
rect 27477 32619 27511 32641
rect 27477 32573 27511 32581
rect 27477 32547 27511 32573
rect 27477 32505 27511 32509
rect 27477 32475 27511 32505
rect 27477 32403 27511 32437
rect 27935 33627 27969 33661
rect 27935 33559 27969 33589
rect 27935 33555 27969 33559
rect 27935 33491 27969 33517
rect 27935 33483 27969 33491
rect 27935 33423 27969 33445
rect 27935 33411 27969 33423
rect 27935 33355 27969 33373
rect 27935 33339 27969 33355
rect 27935 33287 27969 33301
rect 27935 33267 27969 33287
rect 27935 33219 27969 33229
rect 27935 33195 27969 33219
rect 27935 33151 27969 33157
rect 27935 33123 27969 33151
rect 27935 33083 27969 33085
rect 27935 33051 27969 33083
rect 27935 32981 27969 33013
rect 27935 32979 27969 32981
rect 27935 32913 27969 32941
rect 27935 32907 27969 32913
rect 27935 32845 27969 32869
rect 27935 32835 27969 32845
rect 27935 32777 27969 32797
rect 27935 32763 27969 32777
rect 27935 32709 27969 32725
rect 27935 32691 27969 32709
rect 27935 32641 27969 32653
rect 27935 32619 27969 32641
rect 27935 32573 27969 32581
rect 27935 32547 27969 32573
rect 27935 32505 27969 32509
rect 27935 32475 27969 32505
rect 27935 32403 27969 32437
rect 28393 33627 28427 33661
rect 28393 33559 28427 33589
rect 28393 33555 28427 33559
rect 28393 33491 28427 33517
rect 28393 33483 28427 33491
rect 28393 33423 28427 33445
rect 28393 33411 28427 33423
rect 28393 33355 28427 33373
rect 28393 33339 28427 33355
rect 28393 33287 28427 33301
rect 28393 33267 28427 33287
rect 28393 33219 28427 33229
rect 28393 33195 28427 33219
rect 28393 33151 28427 33157
rect 28393 33123 28427 33151
rect 28393 33083 28427 33085
rect 28393 33051 28427 33083
rect 28393 32981 28427 33013
rect 28393 32979 28427 32981
rect 28393 32913 28427 32941
rect 28393 32907 28427 32913
rect 28393 32845 28427 32869
rect 28393 32835 28427 32845
rect 28393 32777 28427 32797
rect 28393 32763 28427 32777
rect 28393 32709 28427 32725
rect 28393 32691 28427 32709
rect 28393 32641 28427 32653
rect 28393 32619 28427 32641
rect 28393 32573 28427 32581
rect 28393 32547 28427 32573
rect 28393 32505 28427 32509
rect 28393 32475 28427 32505
rect 28393 32403 28427 32437
rect 28851 33627 28885 33661
rect 28851 33559 28885 33589
rect 28851 33555 28885 33559
rect 28851 33491 28885 33517
rect 28851 33483 28885 33491
rect 28851 33423 28885 33445
rect 28851 33411 28885 33423
rect 28851 33355 28885 33373
rect 28851 33339 28885 33355
rect 28851 33287 28885 33301
rect 28851 33267 28885 33287
rect 28851 33219 28885 33229
rect 28851 33195 28885 33219
rect 28851 33151 28885 33157
rect 28851 33123 28885 33151
rect 28851 33083 28885 33085
rect 28851 33051 28885 33083
rect 28851 32981 28885 33013
rect 28851 32979 28885 32981
rect 28851 32913 28885 32941
rect 28851 32907 28885 32913
rect 28851 32845 28885 32869
rect 28851 32835 28885 32845
rect 28851 32777 28885 32797
rect 28851 32763 28885 32777
rect 28851 32709 28885 32725
rect 28851 32691 28885 32709
rect 28851 32641 28885 32653
rect 28851 32619 28885 32641
rect 28851 32573 28885 32581
rect 28851 32547 28885 32573
rect 28851 32505 28885 32509
rect 28851 32475 28885 32505
rect 28851 32403 28885 32437
rect 29309 33627 29343 33661
rect 29309 33559 29343 33589
rect 29309 33555 29343 33559
rect 29309 33491 29343 33517
rect 29309 33483 29343 33491
rect 29309 33423 29343 33445
rect 29309 33411 29343 33423
rect 29309 33355 29343 33373
rect 29309 33339 29343 33355
rect 29309 33287 29343 33301
rect 29309 33267 29343 33287
rect 29309 33219 29343 33229
rect 29309 33195 29343 33219
rect 29309 33151 29343 33157
rect 29309 33123 29343 33151
rect 29309 33083 29343 33085
rect 29309 33051 29343 33083
rect 29309 32981 29343 33013
rect 29309 32979 29343 32981
rect 29309 32913 29343 32941
rect 29309 32907 29343 32913
rect 29309 32845 29343 32869
rect 29309 32835 29343 32845
rect 29309 32777 29343 32797
rect 29309 32763 29343 32777
rect 29309 32709 29343 32725
rect 29309 32691 29343 32709
rect 29309 32641 29343 32653
rect 29309 32619 29343 32641
rect 29309 32573 29343 32581
rect 29309 32547 29343 32573
rect 29309 32505 29343 32509
rect 29309 32475 29343 32505
rect 29309 32403 29343 32437
rect 29767 33627 29801 33661
rect 29767 33559 29801 33589
rect 29767 33555 29801 33559
rect 29767 33491 29801 33517
rect 29767 33483 29801 33491
rect 29767 33423 29801 33445
rect 29767 33411 29801 33423
rect 29767 33355 29801 33373
rect 29767 33339 29801 33355
rect 29767 33287 29801 33301
rect 29767 33267 29801 33287
rect 29767 33219 29801 33229
rect 29767 33195 29801 33219
rect 29767 33151 29801 33157
rect 29767 33123 29801 33151
rect 29767 33083 29801 33085
rect 29767 33051 29801 33083
rect 29767 32981 29801 33013
rect 29767 32979 29801 32981
rect 29767 32913 29801 32941
rect 29767 32907 29801 32913
rect 29767 32845 29801 32869
rect 29767 32835 29801 32845
rect 29767 32777 29801 32797
rect 29767 32763 29801 32777
rect 29767 32709 29801 32725
rect 29767 32691 29801 32709
rect 29767 32641 29801 32653
rect 29767 32619 29801 32641
rect 29767 32573 29801 32581
rect 29767 32547 29801 32573
rect 29767 32505 29801 32509
rect 29767 32475 29801 32505
rect 29767 32403 29801 32437
rect 30225 33627 30259 33661
rect 30225 33559 30259 33589
rect 30225 33555 30259 33559
rect 30225 33491 30259 33517
rect 30225 33483 30259 33491
rect 30225 33423 30259 33445
rect 30225 33411 30259 33423
rect 30225 33355 30259 33373
rect 30225 33339 30259 33355
rect 30225 33287 30259 33301
rect 30225 33267 30259 33287
rect 30225 33219 30259 33229
rect 30225 33195 30259 33219
rect 30225 33151 30259 33157
rect 30225 33123 30259 33151
rect 30225 33083 30259 33085
rect 30225 33051 30259 33083
rect 30225 32981 30259 33013
rect 30225 32979 30259 32981
rect 30225 32913 30259 32941
rect 30225 32907 30259 32913
rect 30225 32845 30259 32869
rect 30225 32835 30259 32845
rect 30225 32777 30259 32797
rect 30225 32763 30259 32777
rect 30225 32709 30259 32725
rect 30225 32691 30259 32709
rect 30225 32641 30259 32653
rect 30225 32619 30259 32641
rect 30225 32573 30259 32581
rect 30225 32547 30259 32573
rect 30225 32505 30259 32509
rect 30225 32475 30259 32505
rect 30225 32403 30259 32437
rect 30683 33627 30717 33661
rect 30683 33559 30717 33589
rect 30683 33555 30717 33559
rect 30683 33491 30717 33517
rect 30683 33483 30717 33491
rect 30683 33423 30717 33445
rect 30683 33411 30717 33423
rect 30683 33355 30717 33373
rect 30683 33339 30717 33355
rect 30683 33287 30717 33301
rect 30683 33267 30717 33287
rect 30683 33219 30717 33229
rect 30683 33195 30717 33219
rect 30683 33151 30717 33157
rect 30683 33123 30717 33151
rect 30683 33083 30717 33085
rect 30683 33051 30717 33083
rect 30683 32981 30717 33013
rect 30683 32979 30717 32981
rect 30683 32913 30717 32941
rect 30683 32907 30717 32913
rect 30683 32845 30717 32869
rect 30683 32835 30717 32845
rect 30683 32777 30717 32797
rect 30683 32763 30717 32777
rect 30683 32709 30717 32725
rect 30683 32691 30717 32709
rect 30683 32641 30717 32653
rect 30683 32619 30717 32641
rect 30683 32573 30717 32581
rect 30683 32547 30717 32573
rect 30683 32505 30717 32509
rect 30683 32475 30717 32505
rect 30683 32403 30717 32437
rect 31141 33627 31175 33661
rect 31141 33559 31175 33589
rect 31141 33555 31175 33559
rect 31141 33491 31175 33517
rect 31141 33483 31175 33491
rect 31141 33423 31175 33445
rect 31141 33411 31175 33423
rect 31141 33355 31175 33373
rect 31141 33339 31175 33355
rect 31141 33287 31175 33301
rect 31141 33267 31175 33287
rect 31141 33219 31175 33229
rect 31141 33195 31175 33219
rect 31141 33151 31175 33157
rect 31141 33123 31175 33151
rect 31141 33083 31175 33085
rect 31141 33051 31175 33083
rect 31141 32981 31175 33013
rect 31141 32979 31175 32981
rect 31141 32913 31175 32941
rect 31141 32907 31175 32913
rect 31141 32845 31175 32869
rect 31141 32835 31175 32845
rect 31141 32777 31175 32797
rect 31141 32763 31175 32777
rect 31141 32709 31175 32725
rect 31141 32691 31175 32709
rect 31141 32641 31175 32653
rect 31141 32619 31175 32641
rect 31141 32573 31175 32581
rect 31141 32547 31175 32573
rect 31141 32505 31175 32509
rect 31141 32475 31175 32505
rect 31141 32403 31175 32437
rect 31599 33627 31633 33661
rect 31599 33559 31633 33589
rect 31599 33555 31633 33559
rect 31599 33491 31633 33517
rect 31599 33483 31633 33491
rect 31599 33423 31633 33445
rect 31599 33411 31633 33423
rect 31599 33355 31633 33373
rect 31599 33339 31633 33355
rect 31599 33287 31633 33301
rect 31599 33267 31633 33287
rect 31599 33219 31633 33229
rect 31599 33195 31633 33219
rect 31599 33151 31633 33157
rect 31599 33123 31633 33151
rect 31599 33083 31633 33085
rect 31599 33051 31633 33083
rect 31599 32981 31633 33013
rect 31599 32979 31633 32981
rect 31599 32913 31633 32941
rect 31599 32907 31633 32913
rect 31599 32845 31633 32869
rect 31599 32835 31633 32845
rect 31599 32777 31633 32797
rect 31599 32763 31633 32777
rect 31599 32709 31633 32725
rect 31599 32691 31633 32709
rect 31599 32641 31633 32653
rect 31599 32619 31633 32641
rect 31599 32573 31633 32581
rect 31599 32547 31633 32573
rect 31599 32505 31633 32509
rect 31599 32475 31633 32505
rect 31599 32403 31633 32437
rect 32057 33627 32091 33661
rect 32057 33559 32091 33589
rect 32057 33555 32091 33559
rect 32057 33491 32091 33517
rect 32057 33483 32091 33491
rect 32057 33423 32091 33445
rect 32057 33411 32091 33423
rect 32057 33355 32091 33373
rect 32057 33339 32091 33355
rect 32057 33287 32091 33301
rect 32057 33267 32091 33287
rect 32057 33219 32091 33229
rect 32057 33195 32091 33219
rect 32057 33151 32091 33157
rect 32057 33123 32091 33151
rect 32057 33083 32091 33085
rect 32057 33051 32091 33083
rect 32057 32981 32091 33013
rect 32057 32979 32091 32981
rect 32057 32913 32091 32941
rect 32057 32907 32091 32913
rect 32057 32845 32091 32869
rect 32057 32835 32091 32845
rect 32057 32777 32091 32797
rect 32057 32763 32091 32777
rect 32057 32709 32091 32725
rect 32057 32691 32091 32709
rect 32057 32641 32091 32653
rect 32057 32619 32091 32641
rect 32057 32573 32091 32581
rect 32057 32547 32091 32573
rect 32057 32505 32091 32509
rect 32057 32475 32091 32505
rect 32057 32403 32091 32437
rect 32515 33627 32549 33661
rect 32515 33559 32549 33589
rect 32515 33555 32549 33559
rect 32515 33491 32549 33517
rect 32515 33483 32549 33491
rect 32515 33423 32549 33445
rect 32515 33411 32549 33423
rect 32515 33355 32549 33373
rect 32515 33339 32549 33355
rect 32515 33287 32549 33301
rect 32515 33267 32549 33287
rect 32515 33219 32549 33229
rect 32515 33195 32549 33219
rect 32515 33151 32549 33157
rect 32515 33123 32549 33151
rect 32515 33083 32549 33085
rect 32515 33051 32549 33083
rect 32515 32981 32549 33013
rect 32515 32979 32549 32981
rect 32515 32913 32549 32941
rect 32515 32907 32549 32913
rect 32515 32845 32549 32869
rect 32515 32835 32549 32845
rect 32515 32777 32549 32797
rect 32515 32763 32549 32777
rect 32515 32709 32549 32725
rect 32515 32691 32549 32709
rect 32515 32641 32549 32653
rect 32515 32619 32549 32641
rect 32515 32573 32549 32581
rect 32515 32547 32549 32573
rect 32515 32505 32549 32509
rect 32515 32475 32549 32505
rect 32515 32403 32549 32437
rect 32973 33627 33007 33661
rect 32973 33559 33007 33589
rect 32973 33555 33007 33559
rect 32973 33491 33007 33517
rect 32973 33483 33007 33491
rect 32973 33423 33007 33445
rect 32973 33411 33007 33423
rect 32973 33355 33007 33373
rect 32973 33339 33007 33355
rect 32973 33287 33007 33301
rect 32973 33267 33007 33287
rect 32973 33219 33007 33229
rect 32973 33195 33007 33219
rect 32973 33151 33007 33157
rect 32973 33123 33007 33151
rect 32973 33083 33007 33085
rect 32973 33051 33007 33083
rect 32973 32981 33007 33013
rect 32973 32979 33007 32981
rect 32973 32913 33007 32941
rect 32973 32907 33007 32913
rect 32973 32845 33007 32869
rect 32973 32835 33007 32845
rect 32973 32777 33007 32797
rect 32973 32763 33007 32777
rect 32973 32709 33007 32725
rect 32973 32691 33007 32709
rect 32973 32641 33007 32653
rect 32973 32619 33007 32641
rect 32973 32573 33007 32581
rect 32973 32547 33007 32573
rect 32973 32505 33007 32509
rect 32973 32475 33007 32505
rect 32973 32403 33007 32437
rect 33431 33627 33465 33661
rect 33431 33559 33465 33589
rect 33431 33555 33465 33559
rect 33431 33491 33465 33517
rect 33431 33483 33465 33491
rect 33431 33423 33465 33445
rect 33431 33411 33465 33423
rect 33431 33355 33465 33373
rect 33431 33339 33465 33355
rect 33431 33287 33465 33301
rect 33431 33267 33465 33287
rect 33431 33219 33465 33229
rect 33431 33195 33465 33219
rect 33431 33151 33465 33157
rect 33431 33123 33465 33151
rect 33431 33083 33465 33085
rect 33431 33051 33465 33083
rect 33431 32981 33465 33013
rect 33431 32979 33465 32981
rect 33431 32913 33465 32941
rect 33431 32907 33465 32913
rect 33431 32845 33465 32869
rect 33431 32835 33465 32845
rect 33431 32777 33465 32797
rect 33431 32763 33465 32777
rect 33431 32709 33465 32725
rect 33431 32691 33465 32709
rect 33431 32641 33465 32653
rect 33431 32619 33465 32641
rect 33431 32573 33465 32581
rect 33431 32547 33465 32573
rect 33431 32505 33465 32509
rect 33431 32475 33465 32505
rect 33431 32403 33465 32437
rect 33889 33627 33923 33661
rect 33889 33559 33923 33589
rect 33889 33555 33923 33559
rect 33889 33491 33923 33517
rect 33889 33483 33923 33491
rect 33889 33423 33923 33445
rect 33889 33411 33923 33423
rect 33889 33355 33923 33373
rect 33889 33339 33923 33355
rect 33889 33287 33923 33301
rect 33889 33267 33923 33287
rect 33889 33219 33923 33229
rect 33889 33195 33923 33219
rect 33889 33151 33923 33157
rect 33889 33123 33923 33151
rect 33889 33083 33923 33085
rect 33889 33051 33923 33083
rect 33889 32981 33923 33013
rect 33889 32979 33923 32981
rect 33889 32913 33923 32941
rect 33889 32907 33923 32913
rect 33889 32845 33923 32869
rect 33889 32835 33923 32845
rect 33889 32777 33923 32797
rect 33889 32763 33923 32777
rect 33889 32709 33923 32725
rect 33889 32691 33923 32709
rect 33889 32641 33923 32653
rect 33889 32619 33923 32641
rect 33889 32573 33923 32581
rect 33889 32547 33923 32573
rect 33889 32505 33923 32509
rect 33889 32475 33923 32505
rect 33889 32403 33923 32437
rect 34347 33627 34381 33661
rect 34347 33559 34381 33589
rect 34347 33555 34381 33559
rect 34347 33491 34381 33517
rect 34347 33483 34381 33491
rect 34347 33423 34381 33445
rect 34347 33411 34381 33423
rect 34347 33355 34381 33373
rect 34347 33339 34381 33355
rect 34347 33287 34381 33301
rect 34347 33267 34381 33287
rect 34347 33219 34381 33229
rect 34347 33195 34381 33219
rect 34347 33151 34381 33157
rect 34347 33123 34381 33151
rect 34347 33083 34381 33085
rect 34347 33051 34381 33083
rect 34347 32981 34381 33013
rect 34347 32979 34381 32981
rect 34347 32913 34381 32941
rect 34347 32907 34381 32913
rect 34347 32845 34381 32869
rect 34347 32835 34381 32845
rect 34347 32777 34381 32797
rect 34347 32763 34381 32777
rect 34347 32709 34381 32725
rect 34347 32691 34381 32709
rect 34347 32641 34381 32653
rect 34347 32619 34381 32641
rect 34347 32573 34381 32581
rect 34347 32547 34381 32573
rect 34347 32505 34381 32509
rect 34347 32475 34381 32505
rect 34347 32403 34381 32437
rect 34805 33627 34839 33661
rect 34805 33559 34839 33589
rect 34805 33555 34839 33559
rect 34805 33491 34839 33517
rect 34805 33483 34839 33491
rect 34805 33423 34839 33445
rect 34805 33411 34839 33423
rect 34805 33355 34839 33373
rect 34805 33339 34839 33355
rect 34805 33287 34839 33301
rect 34805 33267 34839 33287
rect 34805 33219 34839 33229
rect 34805 33195 34839 33219
rect 34805 33151 34839 33157
rect 34805 33123 34839 33151
rect 34805 33083 34839 33085
rect 34805 33051 34839 33083
rect 34805 32981 34839 33013
rect 34805 32979 34839 32981
rect 34805 32913 34839 32941
rect 34805 32907 34839 32913
rect 34805 32845 34839 32869
rect 34805 32835 34839 32845
rect 34805 32777 34839 32797
rect 34805 32763 34839 32777
rect 34805 32709 34839 32725
rect 34805 32691 34839 32709
rect 34805 32641 34839 32653
rect 34805 32619 34839 32641
rect 34805 32573 34839 32581
rect 34805 32547 34839 32573
rect 34805 32505 34839 32509
rect 34805 32475 34839 32505
rect 34805 32403 34839 32437
rect 35263 33627 35297 33661
rect 35263 33559 35297 33589
rect 35263 33555 35297 33559
rect 35263 33491 35297 33517
rect 35263 33483 35297 33491
rect 35263 33423 35297 33445
rect 35263 33411 35297 33423
rect 35263 33355 35297 33373
rect 35263 33339 35297 33355
rect 35263 33287 35297 33301
rect 35263 33267 35297 33287
rect 35263 33219 35297 33229
rect 35263 33195 35297 33219
rect 35263 33151 35297 33157
rect 35263 33123 35297 33151
rect 35263 33083 35297 33085
rect 35263 33051 35297 33083
rect 35263 32981 35297 33013
rect 35263 32979 35297 32981
rect 35263 32913 35297 32941
rect 35263 32907 35297 32913
rect 35263 32845 35297 32869
rect 35263 32835 35297 32845
rect 35263 32777 35297 32797
rect 35263 32763 35297 32777
rect 35263 32709 35297 32725
rect 35263 32691 35297 32709
rect 35263 32641 35297 32653
rect 35263 32619 35297 32641
rect 35263 32573 35297 32581
rect 35263 32547 35297 32573
rect 35263 32505 35297 32509
rect 35263 32475 35297 32505
rect 35263 32403 35297 32437
rect 35721 33627 35755 33661
rect 35721 33559 35755 33589
rect 35721 33555 35755 33559
rect 35721 33491 35755 33517
rect 35721 33483 35755 33491
rect 35721 33423 35755 33445
rect 35721 33411 35755 33423
rect 35721 33355 35755 33373
rect 35721 33339 35755 33355
rect 35721 33287 35755 33301
rect 35721 33267 35755 33287
rect 35721 33219 35755 33229
rect 35721 33195 35755 33219
rect 35721 33151 35755 33157
rect 35721 33123 35755 33151
rect 35721 33083 35755 33085
rect 35721 33051 35755 33083
rect 35721 32981 35755 33013
rect 35721 32979 35755 32981
rect 35721 32913 35755 32941
rect 35721 32907 35755 32913
rect 35721 32845 35755 32869
rect 35721 32835 35755 32845
rect 35721 32777 35755 32797
rect 35721 32763 35755 32777
rect 35721 32709 35755 32725
rect 35721 32691 35755 32709
rect 35721 32641 35755 32653
rect 35721 32619 35755 32641
rect 35721 32573 35755 32581
rect 35721 32547 35755 32573
rect 35721 32505 35755 32509
rect 35721 32475 35755 32505
rect 35721 32403 35755 32437
rect 36179 33627 36213 33661
rect 36179 33559 36213 33589
rect 36179 33555 36213 33559
rect 36179 33491 36213 33517
rect 36179 33483 36213 33491
rect 36179 33423 36213 33445
rect 36179 33411 36213 33423
rect 36179 33355 36213 33373
rect 36179 33339 36213 33355
rect 36179 33287 36213 33301
rect 36179 33267 36213 33287
rect 36179 33219 36213 33229
rect 36179 33195 36213 33219
rect 36179 33151 36213 33157
rect 36179 33123 36213 33151
rect 36179 33083 36213 33085
rect 36179 33051 36213 33083
rect 36179 32981 36213 33013
rect 36179 32979 36213 32981
rect 36179 32913 36213 32941
rect 36179 32907 36213 32913
rect 36179 32845 36213 32869
rect 36179 32835 36213 32845
rect 36179 32777 36213 32797
rect 36179 32763 36213 32777
rect 36179 32709 36213 32725
rect 36179 32691 36213 32709
rect 36179 32641 36213 32653
rect 36179 32619 36213 32641
rect 36179 32573 36213 32581
rect 36179 32547 36213 32573
rect 36179 32505 36213 32509
rect 36179 32475 36213 32505
rect 36179 32403 36213 32437
rect 36637 33627 36671 33661
rect 36637 33559 36671 33589
rect 36637 33555 36671 33559
rect 36637 33491 36671 33517
rect 36637 33483 36671 33491
rect 36637 33423 36671 33445
rect 36637 33411 36671 33423
rect 36637 33355 36671 33373
rect 36637 33339 36671 33355
rect 36637 33287 36671 33301
rect 36637 33267 36671 33287
rect 36637 33219 36671 33229
rect 36637 33195 36671 33219
rect 36637 33151 36671 33157
rect 36637 33123 36671 33151
rect 36637 33083 36671 33085
rect 36637 33051 36671 33083
rect 36637 32981 36671 33013
rect 36637 32979 36671 32981
rect 36637 32913 36671 32941
rect 36637 32907 36671 32913
rect 36637 32845 36671 32869
rect 36637 32835 36671 32845
rect 36637 32777 36671 32797
rect 36637 32763 36671 32777
rect 36637 32709 36671 32725
rect 36637 32691 36671 32709
rect 36637 32641 36671 32653
rect 36637 32619 36671 32641
rect 36637 32573 36671 32581
rect 36637 32547 36671 32573
rect 36637 32505 36671 32509
rect 36637 32475 36671 32505
rect 36637 32403 36671 32437
rect 37095 33627 37129 33661
rect 37095 33559 37129 33589
rect 37095 33555 37129 33559
rect 37095 33491 37129 33517
rect 37095 33483 37129 33491
rect 37095 33423 37129 33445
rect 37095 33411 37129 33423
rect 37095 33355 37129 33373
rect 37095 33339 37129 33355
rect 37095 33287 37129 33301
rect 37095 33267 37129 33287
rect 37095 33219 37129 33229
rect 37095 33195 37129 33219
rect 37095 33151 37129 33157
rect 37095 33123 37129 33151
rect 37095 33083 37129 33085
rect 37095 33051 37129 33083
rect 37095 32981 37129 33013
rect 37095 32979 37129 32981
rect 37095 32913 37129 32941
rect 37095 32907 37129 32913
rect 37095 32845 37129 32869
rect 37095 32835 37129 32845
rect 37095 32777 37129 32797
rect 37095 32763 37129 32777
rect 37095 32709 37129 32725
rect 37095 32691 37129 32709
rect 37095 32641 37129 32653
rect 37095 32619 37129 32641
rect 37095 32573 37129 32581
rect 37095 32547 37129 32573
rect 37095 32505 37129 32509
rect 37095 32475 37129 32505
rect 37095 32403 37129 32437
rect 37553 33627 37587 33661
rect 37553 33559 37587 33589
rect 37553 33555 37587 33559
rect 37553 33491 37587 33517
rect 37553 33483 37587 33491
rect 37553 33423 37587 33445
rect 37553 33411 37587 33423
rect 37553 33355 37587 33373
rect 37553 33339 37587 33355
rect 37553 33287 37587 33301
rect 37553 33267 37587 33287
rect 37553 33219 37587 33229
rect 37553 33195 37587 33219
rect 37553 33151 37587 33157
rect 37553 33123 37587 33151
rect 37553 33083 37587 33085
rect 37553 33051 37587 33083
rect 37553 32981 37587 33013
rect 37553 32979 37587 32981
rect 37553 32913 37587 32941
rect 37553 32907 37587 32913
rect 37553 32845 37587 32869
rect 37553 32835 37587 32845
rect 37553 32777 37587 32797
rect 37553 32763 37587 32777
rect 37553 32709 37587 32725
rect 37553 32691 37587 32709
rect 37553 32641 37587 32653
rect 37553 32619 37587 32641
rect 37553 32573 37587 32581
rect 37553 32547 37587 32573
rect 37553 32505 37587 32509
rect 37553 32475 37587 32505
rect 37553 32403 37587 32437
rect 38011 33627 38045 33661
rect 38011 33559 38045 33589
rect 38011 33555 38045 33559
rect 38011 33491 38045 33517
rect 38011 33483 38045 33491
rect 38011 33423 38045 33445
rect 38011 33411 38045 33423
rect 38011 33355 38045 33373
rect 38011 33339 38045 33355
rect 38011 33287 38045 33301
rect 38011 33267 38045 33287
rect 38011 33219 38045 33229
rect 38011 33195 38045 33219
rect 38011 33151 38045 33157
rect 38011 33123 38045 33151
rect 38011 33083 38045 33085
rect 38011 33051 38045 33083
rect 38011 32981 38045 33013
rect 38011 32979 38045 32981
rect 38011 32913 38045 32941
rect 38011 32907 38045 32913
rect 38011 32845 38045 32869
rect 38011 32835 38045 32845
rect 38011 32777 38045 32797
rect 38011 32763 38045 32777
rect 38011 32709 38045 32725
rect 38011 32691 38045 32709
rect 38011 32641 38045 32653
rect 38011 32619 38045 32641
rect 38011 32573 38045 32581
rect 38011 32547 38045 32573
rect 38011 32505 38045 32509
rect 38011 32475 38045 32505
rect 38011 32403 38045 32437
rect 38469 33627 38503 33661
rect 38469 33559 38503 33589
rect 38469 33555 38503 33559
rect 38469 33491 38503 33517
rect 38469 33483 38503 33491
rect 38469 33423 38503 33445
rect 38469 33411 38503 33423
rect 38469 33355 38503 33373
rect 38469 33339 38503 33355
rect 38469 33287 38503 33301
rect 38469 33267 38503 33287
rect 38469 33219 38503 33229
rect 38469 33195 38503 33219
rect 38469 33151 38503 33157
rect 38469 33123 38503 33151
rect 38469 33083 38503 33085
rect 38469 33051 38503 33083
rect 38469 32981 38503 33013
rect 38469 32979 38503 32981
rect 38469 32913 38503 32941
rect 38469 32907 38503 32913
rect 38469 32845 38503 32869
rect 38469 32835 38503 32845
rect 38469 32777 38503 32797
rect 38469 32763 38503 32777
rect 38469 32709 38503 32725
rect 38469 32691 38503 32709
rect 38469 32641 38503 32653
rect 38469 32619 38503 32641
rect 38469 32573 38503 32581
rect 38469 32547 38503 32573
rect 38469 32505 38503 32509
rect 38469 32475 38503 32505
rect 38469 32403 38503 32437
rect 38927 33627 38961 33661
rect 38927 33559 38961 33589
rect 38927 33555 38961 33559
rect 38927 33491 38961 33517
rect 38927 33483 38961 33491
rect 38927 33423 38961 33445
rect 38927 33411 38961 33423
rect 38927 33355 38961 33373
rect 38927 33339 38961 33355
rect 38927 33287 38961 33301
rect 38927 33267 38961 33287
rect 38927 33219 38961 33229
rect 38927 33195 38961 33219
rect 38927 33151 38961 33157
rect 38927 33123 38961 33151
rect 38927 33083 38961 33085
rect 38927 33051 38961 33083
rect 38927 32981 38961 33013
rect 38927 32979 38961 32981
rect 38927 32913 38961 32941
rect 38927 32907 38961 32913
rect 38927 32845 38961 32869
rect 38927 32835 38961 32845
rect 38927 32777 38961 32797
rect 38927 32763 38961 32777
rect 38927 32709 38961 32725
rect 38927 32691 38961 32709
rect 38927 32641 38961 32653
rect 38927 32619 38961 32641
rect 38927 32573 38961 32581
rect 38927 32547 38961 32573
rect 38927 32505 38961 32509
rect 38927 32475 38961 32505
rect 38927 32403 38961 32437
rect 39385 33627 39419 33661
rect 39385 33559 39419 33589
rect 39385 33555 39419 33559
rect 39385 33491 39419 33517
rect 39385 33483 39419 33491
rect 39385 33423 39419 33445
rect 39385 33411 39419 33423
rect 39385 33355 39419 33373
rect 39385 33339 39419 33355
rect 39385 33287 39419 33301
rect 39385 33267 39419 33287
rect 39385 33219 39419 33229
rect 39385 33195 39419 33219
rect 39385 33151 39419 33157
rect 39385 33123 39419 33151
rect 39385 33083 39419 33085
rect 39385 33051 39419 33083
rect 39385 32981 39419 33013
rect 39385 32979 39419 32981
rect 39385 32913 39419 32941
rect 39385 32907 39419 32913
rect 39385 32845 39419 32869
rect 39385 32835 39419 32845
rect 39385 32777 39419 32797
rect 39385 32763 39419 32777
rect 39385 32709 39419 32725
rect 39385 32691 39419 32709
rect 39385 32641 39419 32653
rect 39385 32619 39419 32641
rect 39385 32573 39419 32581
rect 39385 32547 39419 32573
rect 39385 32505 39419 32509
rect 39385 32475 39419 32505
rect 39385 32403 39419 32437
rect 39843 33627 39877 33661
rect 39843 33559 39877 33589
rect 39843 33555 39877 33559
rect 39843 33491 39877 33517
rect 39843 33483 39877 33491
rect 39843 33423 39877 33445
rect 39843 33411 39877 33423
rect 39843 33355 39877 33373
rect 39843 33339 39877 33355
rect 39843 33287 39877 33301
rect 39843 33267 39877 33287
rect 39843 33219 39877 33229
rect 39843 33195 39877 33219
rect 39843 33151 39877 33157
rect 39843 33123 39877 33151
rect 39843 33083 39877 33085
rect 39843 33051 39877 33083
rect 39843 32981 39877 33013
rect 39843 32979 39877 32981
rect 39843 32913 39877 32941
rect 39843 32907 39877 32913
rect 39843 32845 39877 32869
rect 39843 32835 39877 32845
rect 39843 32777 39877 32797
rect 39843 32763 39877 32777
rect 39843 32709 39877 32725
rect 39843 32691 39877 32709
rect 39843 32641 39877 32653
rect 39843 32619 39877 32641
rect 39843 32573 39877 32581
rect 39843 32547 39877 32573
rect 39843 32505 39877 32509
rect 39843 32475 39877 32505
rect 39843 32403 39877 32437
rect 40301 33627 40335 33661
rect 40301 33559 40335 33589
rect 40301 33555 40335 33559
rect 40301 33491 40335 33517
rect 40301 33483 40335 33491
rect 40301 33423 40335 33445
rect 40301 33411 40335 33423
rect 40301 33355 40335 33373
rect 40301 33339 40335 33355
rect 40301 33287 40335 33301
rect 40301 33267 40335 33287
rect 40301 33219 40335 33229
rect 40301 33195 40335 33219
rect 40301 33151 40335 33157
rect 40301 33123 40335 33151
rect 40301 33083 40335 33085
rect 40301 33051 40335 33083
rect 40301 32981 40335 33013
rect 40301 32979 40335 32981
rect 40301 32913 40335 32941
rect 40301 32907 40335 32913
rect 40301 32845 40335 32869
rect 40301 32835 40335 32845
rect 40301 32777 40335 32797
rect 40301 32763 40335 32777
rect 40301 32709 40335 32725
rect 40301 32691 40335 32709
rect 40301 32641 40335 32653
rect 40301 32619 40335 32641
rect 40301 32573 40335 32581
rect 40301 32547 40335 32573
rect 40301 32505 40335 32509
rect 40301 32475 40335 32505
rect 40301 32403 40335 32437
rect 40759 33627 40793 33661
rect 40759 33559 40793 33589
rect 40759 33555 40793 33559
rect 40759 33491 40793 33517
rect 40759 33483 40793 33491
rect 40759 33423 40793 33445
rect 40759 33411 40793 33423
rect 40759 33355 40793 33373
rect 40759 33339 40793 33355
rect 40759 33287 40793 33301
rect 40759 33267 40793 33287
rect 40759 33219 40793 33229
rect 40759 33195 40793 33219
rect 40759 33151 40793 33157
rect 40759 33123 40793 33151
rect 40759 33083 40793 33085
rect 40759 33051 40793 33083
rect 40759 32981 40793 33013
rect 40759 32979 40793 32981
rect 40759 32913 40793 32941
rect 40759 32907 40793 32913
rect 40759 32845 40793 32869
rect 40759 32835 40793 32845
rect 40759 32777 40793 32797
rect 40759 32763 40793 32777
rect 40759 32709 40793 32725
rect 40759 32691 40793 32709
rect 40759 32641 40793 32653
rect 40759 32619 40793 32641
rect 40759 32573 40793 32581
rect 40759 32547 40793 32573
rect 40759 32505 40793 32509
rect 40759 32475 40793 32505
rect 40759 32403 40793 32437
rect 41217 33627 41251 33661
rect 41217 33559 41251 33589
rect 41217 33555 41251 33559
rect 41217 33491 41251 33517
rect 41217 33483 41251 33491
rect 41217 33423 41251 33445
rect 41217 33411 41251 33423
rect 41217 33355 41251 33373
rect 41217 33339 41251 33355
rect 41217 33287 41251 33301
rect 41217 33267 41251 33287
rect 41217 33219 41251 33229
rect 41217 33195 41251 33219
rect 41217 33151 41251 33157
rect 41217 33123 41251 33151
rect 41217 33083 41251 33085
rect 41217 33051 41251 33083
rect 41217 32981 41251 33013
rect 41217 32979 41251 32981
rect 41217 32913 41251 32941
rect 41217 32907 41251 32913
rect 41217 32845 41251 32869
rect 41217 32835 41251 32845
rect 41217 32777 41251 32797
rect 41217 32763 41251 32777
rect 41217 32709 41251 32725
rect 41217 32691 41251 32709
rect 41217 32641 41251 32653
rect 41217 32619 41251 32641
rect 41217 32573 41251 32581
rect 41217 32547 41251 32573
rect 41217 32505 41251 32509
rect 41217 32475 41251 32505
rect 41217 32403 41251 32437
rect 41675 33627 41709 33661
rect 41675 33559 41709 33589
rect 41675 33555 41709 33559
rect 41675 33491 41709 33517
rect 41675 33483 41709 33491
rect 41675 33423 41709 33445
rect 41675 33411 41709 33423
rect 41675 33355 41709 33373
rect 41675 33339 41709 33355
rect 41675 33287 41709 33301
rect 41675 33267 41709 33287
rect 41675 33219 41709 33229
rect 41675 33195 41709 33219
rect 41675 33151 41709 33157
rect 41675 33123 41709 33151
rect 41675 33083 41709 33085
rect 41675 33051 41709 33083
rect 41675 32981 41709 33013
rect 41675 32979 41709 32981
rect 41675 32913 41709 32941
rect 41675 32907 41709 32913
rect 41675 32845 41709 32869
rect 41675 32835 41709 32845
rect 41675 32777 41709 32797
rect 41675 32763 41709 32777
rect 41675 32709 41709 32725
rect 41675 32691 41709 32709
rect 41675 32641 41709 32653
rect 41675 32619 41709 32641
rect 41675 32573 41709 32581
rect 41675 32547 41709 32573
rect 41675 32505 41709 32509
rect 41675 32475 41709 32505
rect 41675 32403 41709 32437
rect 26893 32249 26927 32283
rect 14197 32147 14231 32181
rect 6787 32015 6821 32049
rect 7187 32015 7221 32049
rect 7587 32015 7621 32049
rect 7987 32015 8021 32049
rect 8387 32015 8421 32049
rect 8787 32015 8821 32049
rect 9187 32015 9221 32049
rect 9587 32015 9621 32049
rect 9987 32015 10021 32049
rect 10387 32015 10421 32049
rect 10787 32015 10821 32049
rect 11187 32015 11221 32049
rect 11587 32015 11621 32049
rect 11987 32015 12021 32049
rect 12387 32015 12421 32049
rect 12787 32015 12821 32049
rect 13187 32015 13221 32049
rect 13587 32015 13621 32049
rect 14331 32015 14365 32049
rect 14731 32015 14765 32049
rect 15131 32015 15165 32049
rect 15531 32015 15565 32049
rect 15931 32015 15965 32049
rect 16331 32015 16365 32049
rect 16731 32015 16765 32049
rect 17131 32015 17165 32049
rect 17531 32015 17565 32049
rect 17931 32015 17965 32049
rect 18331 32015 18365 32049
rect 18731 32015 18765 32049
rect 19131 32015 19165 32049
rect 19531 32015 19565 32049
rect 19931 32015 19965 32049
rect 20331 32015 20365 32049
rect 20731 32015 20765 32049
rect 21131 32015 21165 32049
rect 21531 32015 21565 32049
rect 21931 32015 21965 32049
rect 22331 32015 22365 32049
rect 22731 32015 22765 32049
rect 23131 32015 23165 32049
rect 23531 32015 23565 32049
rect 23931 32015 23965 32049
rect 24331 32015 24365 32049
rect 24731 32015 24765 32049
rect 25131 32015 25165 32049
rect 25531 32015 25565 32049
rect 25931 32015 25965 32049
rect 26331 32015 26365 32049
rect 26731 32015 26765 32049
rect 27131 32015 27165 32049
rect 27531 32015 27565 32049
rect 27931 32015 27965 32049
rect 28331 32015 28365 32049
rect 28731 32015 28765 32049
rect 29131 32015 29165 32049
rect 29531 32015 29565 32049
rect 29931 32015 29965 32049
rect 30331 32015 30365 32049
rect 30731 32015 30765 32049
rect 31131 32015 31165 32049
rect 31531 32015 31565 32049
rect 31931 32015 31965 32049
rect 32331 32015 32365 32049
rect 32731 32015 32765 32049
rect 33131 32015 33165 32049
rect 33531 32015 33565 32049
rect 33931 32015 33965 32049
rect 34331 32015 34365 32049
rect 34731 32015 34765 32049
rect 35131 32015 35165 32049
rect 35531 32015 35565 32049
rect 35931 32015 35965 32049
rect 36331 32015 36365 32049
rect 36731 32015 36765 32049
rect 37131 32015 37165 32049
rect 37531 32015 37565 32049
rect 37931 32015 37965 32049
rect 38331 32015 38365 32049
rect 38731 32015 38765 32049
rect 39131 32015 39165 32049
rect 39531 32015 39565 32049
rect 39931 32015 39965 32049
rect 40331 32015 40365 32049
rect 40731 32015 40765 32049
rect 41131 32015 41165 32049
rect 41531 32015 41565 32049
rect 6197 30135 6231 30169
rect 6597 30135 6631 30169
rect 6997 30135 7031 30169
rect 7397 30135 7431 30169
rect 7797 30135 7831 30169
rect 8197 30135 8231 30169
rect 8597 30135 8631 30169
rect 8997 30135 9031 30169
rect 9397 30135 9431 30169
rect 9797 30135 9831 30169
rect 10197 30135 10231 30169
rect 10597 30135 10631 30169
rect 10997 30135 11031 30169
rect 11397 30135 11431 30169
rect 11797 30135 11831 30169
rect 12197 30135 12231 30169
rect 12597 30135 12631 30169
rect 12997 30135 13031 30169
rect 13397 30135 13431 30169
rect 13797 30135 13831 30169
rect 14197 30135 14231 30169
rect 14597 30135 14631 30169
rect 14997 30135 15031 30169
rect 15397 30135 15431 30169
rect 15797 30135 15831 30169
rect 16197 30135 16231 30169
rect 16597 30135 16631 30169
rect 16997 30135 17031 30169
rect 17397 30135 17431 30169
rect 17797 30135 17831 30169
rect 18197 30135 18231 30169
rect 18597 30135 18631 30169
rect 18997 30135 19031 30169
rect 19397 30135 19431 30169
rect 19797 30135 19831 30169
rect 20197 30135 20231 30169
rect 20597 30135 20631 30169
rect 20997 30135 21031 30169
rect 21397 30135 21431 30169
rect 21797 30135 21831 30169
rect 22197 30135 22231 30169
rect 22597 30135 22631 30169
rect 22997 30135 23031 30169
rect 23397 30135 23431 30169
rect 23797 30135 23831 30169
rect 24197 30135 24231 30169
rect 24597 30135 24631 30169
rect 24997 30135 25031 30169
rect 25397 30135 25431 30169
rect 25797 30135 25831 30169
rect 26197 30135 26231 30169
rect 26597 30135 26631 30169
rect 26997 30135 27031 30169
rect 27397 30135 27431 30169
rect 27797 30135 27831 30169
rect 28197 30135 28231 30169
rect 28597 30135 28631 30169
rect 28997 30135 29031 30169
rect 29397 30135 29431 30169
rect 29797 30135 29831 30169
rect 30197 30135 30231 30169
rect 30597 30135 30631 30169
rect 30997 30135 31031 30169
rect 31397 30135 31431 30169
rect 31797 30135 31831 30169
rect 32197 30135 32231 30169
rect 32597 30135 32631 30169
rect 32997 30135 33031 30169
rect 33397 30135 33431 30169
rect 34225 30135 34259 30169
rect 34625 30135 34659 30169
rect 35025 30135 35059 30169
rect 35425 30135 35459 30169
rect 35825 30135 35859 30169
rect 36225 30135 36259 30169
rect 36625 30135 36659 30169
rect 37577 30135 37611 30169
rect 37777 30135 37811 30169
rect 37977 30135 38011 30169
rect 38177 30135 38211 30169
rect 38377 30135 38411 30169
rect 38577 30135 38611 30169
rect 38777 30135 38811 30169
rect 38977 30135 39011 30169
rect 39177 30135 39211 30169
rect 39377 30135 39411 30169
rect 39577 30135 39611 30169
rect 40321 30135 40355 30169
rect 40521 30135 40555 30169
rect 40721 30135 40755 30169
rect 40921 30135 40955 30169
rect 41121 30135 41155 30169
rect 41321 30135 41355 30169
rect 41521 30135 41555 30169
rect 41721 30135 41755 30169
rect 41921 30135 41955 30169
rect 42121 30135 42155 30169
rect 42321 30135 42355 30169
rect 6061 29867 6095 29901
rect 6061 29799 6095 29829
rect 6061 29795 6095 29799
rect 6061 29731 6095 29757
rect 6061 29723 6095 29731
rect 6061 29663 6095 29685
rect 6061 29651 6095 29663
rect 6061 29595 6095 29613
rect 6061 29579 6095 29595
rect 6061 29527 6095 29541
rect 6061 29507 6095 29527
rect 6061 29459 6095 29469
rect 6061 29435 6095 29459
rect 6061 29391 6095 29397
rect 6061 29363 6095 29391
rect 6061 29323 6095 29325
rect 6061 29291 6095 29323
rect 6061 29221 6095 29253
rect 6061 29219 6095 29221
rect 6061 29153 6095 29181
rect 6061 29147 6095 29153
rect 6061 29085 6095 29109
rect 6061 29075 6095 29085
rect 6061 29017 6095 29037
rect 6061 29003 6095 29017
rect 6061 28949 6095 28965
rect 6061 28931 6095 28949
rect 6061 28881 6095 28893
rect 6061 28859 6095 28881
rect 6061 28813 6095 28821
rect 6061 28787 6095 28813
rect 6061 28745 6095 28749
rect 6061 28715 6095 28745
rect 6061 28643 6095 28677
rect 6519 29867 6553 29901
rect 6519 29799 6553 29829
rect 6519 29795 6553 29799
rect 6519 29731 6553 29757
rect 6519 29723 6553 29731
rect 6519 29663 6553 29685
rect 6519 29651 6553 29663
rect 6519 29595 6553 29613
rect 6519 29579 6553 29595
rect 6519 29527 6553 29541
rect 6519 29507 6553 29527
rect 6519 29459 6553 29469
rect 6519 29435 6553 29459
rect 6519 29391 6553 29397
rect 6519 29363 6553 29391
rect 6519 29323 6553 29325
rect 6519 29291 6553 29323
rect 6519 29221 6553 29253
rect 6519 29219 6553 29221
rect 6519 29153 6553 29181
rect 6519 29147 6553 29153
rect 6519 29085 6553 29109
rect 6519 29075 6553 29085
rect 6519 29017 6553 29037
rect 6519 29003 6553 29017
rect 6519 28949 6553 28965
rect 6519 28931 6553 28949
rect 6519 28881 6553 28893
rect 6519 28859 6553 28881
rect 6519 28813 6553 28821
rect 6519 28787 6553 28813
rect 6519 28745 6553 28749
rect 6519 28715 6553 28745
rect 6519 28643 6553 28677
rect 6977 29867 7011 29901
rect 6977 29799 7011 29829
rect 6977 29795 7011 29799
rect 6977 29731 7011 29757
rect 6977 29723 7011 29731
rect 6977 29663 7011 29685
rect 6977 29651 7011 29663
rect 6977 29595 7011 29613
rect 6977 29579 7011 29595
rect 6977 29527 7011 29541
rect 6977 29507 7011 29527
rect 6977 29459 7011 29469
rect 6977 29435 7011 29459
rect 6977 29391 7011 29397
rect 6977 29363 7011 29391
rect 6977 29323 7011 29325
rect 6977 29291 7011 29323
rect 6977 29221 7011 29253
rect 6977 29219 7011 29221
rect 6977 29153 7011 29181
rect 6977 29147 7011 29153
rect 6977 29085 7011 29109
rect 6977 29075 7011 29085
rect 6977 29017 7011 29037
rect 6977 29003 7011 29017
rect 6977 28949 7011 28965
rect 6977 28931 7011 28949
rect 6977 28881 7011 28893
rect 6977 28859 7011 28881
rect 6977 28813 7011 28821
rect 6977 28787 7011 28813
rect 6977 28745 7011 28749
rect 6977 28715 7011 28745
rect 6977 28643 7011 28677
rect 7435 29867 7469 29901
rect 7435 29799 7469 29829
rect 7435 29795 7469 29799
rect 7435 29731 7469 29757
rect 7435 29723 7469 29731
rect 7435 29663 7469 29685
rect 7435 29651 7469 29663
rect 7435 29595 7469 29613
rect 7435 29579 7469 29595
rect 7435 29527 7469 29541
rect 7435 29507 7469 29527
rect 7435 29459 7469 29469
rect 7435 29435 7469 29459
rect 7435 29391 7469 29397
rect 7435 29363 7469 29391
rect 7435 29323 7469 29325
rect 7435 29291 7469 29323
rect 7435 29221 7469 29253
rect 7435 29219 7469 29221
rect 7435 29153 7469 29181
rect 7435 29147 7469 29153
rect 7435 29085 7469 29109
rect 7435 29075 7469 29085
rect 7435 29017 7469 29037
rect 7435 29003 7469 29017
rect 7435 28949 7469 28965
rect 7435 28931 7469 28949
rect 7435 28881 7469 28893
rect 7435 28859 7469 28881
rect 7435 28813 7469 28821
rect 7435 28787 7469 28813
rect 7435 28745 7469 28749
rect 7435 28715 7469 28745
rect 7435 28643 7469 28677
rect 7893 29867 7927 29901
rect 7893 29799 7927 29829
rect 7893 29795 7927 29799
rect 7893 29731 7927 29757
rect 7893 29723 7927 29731
rect 7893 29663 7927 29685
rect 7893 29651 7927 29663
rect 7893 29595 7927 29613
rect 7893 29579 7927 29595
rect 7893 29527 7927 29541
rect 7893 29507 7927 29527
rect 7893 29459 7927 29469
rect 7893 29435 7927 29459
rect 7893 29391 7927 29397
rect 7893 29363 7927 29391
rect 7893 29323 7927 29325
rect 7893 29291 7927 29323
rect 7893 29221 7927 29253
rect 7893 29219 7927 29221
rect 7893 29153 7927 29181
rect 7893 29147 7927 29153
rect 7893 29085 7927 29109
rect 7893 29075 7927 29085
rect 7893 29017 7927 29037
rect 7893 29003 7927 29017
rect 7893 28949 7927 28965
rect 7893 28931 7927 28949
rect 7893 28881 7927 28893
rect 7893 28859 7927 28881
rect 7893 28813 7927 28821
rect 7893 28787 7927 28813
rect 7893 28745 7927 28749
rect 7893 28715 7927 28745
rect 7893 28643 7927 28677
rect 8351 29867 8385 29901
rect 8351 29799 8385 29829
rect 8351 29795 8385 29799
rect 8351 29731 8385 29757
rect 8351 29723 8385 29731
rect 8351 29663 8385 29685
rect 8351 29651 8385 29663
rect 8351 29595 8385 29613
rect 8351 29579 8385 29595
rect 8351 29527 8385 29541
rect 8351 29507 8385 29527
rect 8351 29459 8385 29469
rect 8351 29435 8385 29459
rect 8351 29391 8385 29397
rect 8351 29363 8385 29391
rect 8351 29323 8385 29325
rect 8351 29291 8385 29323
rect 8351 29221 8385 29253
rect 8351 29219 8385 29221
rect 8351 29153 8385 29181
rect 8351 29147 8385 29153
rect 8351 29085 8385 29109
rect 8351 29075 8385 29085
rect 8351 29017 8385 29037
rect 8351 29003 8385 29017
rect 8351 28949 8385 28965
rect 8351 28931 8385 28949
rect 8351 28881 8385 28893
rect 8351 28859 8385 28881
rect 8351 28813 8385 28821
rect 8351 28787 8385 28813
rect 8351 28745 8385 28749
rect 8351 28715 8385 28745
rect 8351 28643 8385 28677
rect 8809 29867 8843 29901
rect 8809 29799 8843 29829
rect 8809 29795 8843 29799
rect 8809 29731 8843 29757
rect 8809 29723 8843 29731
rect 8809 29663 8843 29685
rect 8809 29651 8843 29663
rect 8809 29595 8843 29613
rect 8809 29579 8843 29595
rect 8809 29527 8843 29541
rect 8809 29507 8843 29527
rect 8809 29459 8843 29469
rect 8809 29435 8843 29459
rect 8809 29391 8843 29397
rect 8809 29363 8843 29391
rect 8809 29323 8843 29325
rect 8809 29291 8843 29323
rect 8809 29221 8843 29253
rect 8809 29219 8843 29221
rect 8809 29153 8843 29181
rect 8809 29147 8843 29153
rect 8809 29085 8843 29109
rect 8809 29075 8843 29085
rect 8809 29017 8843 29037
rect 8809 29003 8843 29017
rect 8809 28949 8843 28965
rect 8809 28931 8843 28949
rect 8809 28881 8843 28893
rect 8809 28859 8843 28881
rect 8809 28813 8843 28821
rect 8809 28787 8843 28813
rect 8809 28745 8843 28749
rect 8809 28715 8843 28745
rect 8809 28643 8843 28677
rect 9267 29867 9301 29901
rect 9267 29799 9301 29829
rect 9267 29795 9301 29799
rect 9267 29731 9301 29757
rect 9267 29723 9301 29731
rect 9267 29663 9301 29685
rect 9267 29651 9301 29663
rect 9267 29595 9301 29613
rect 9267 29579 9301 29595
rect 9267 29527 9301 29541
rect 9267 29507 9301 29527
rect 9267 29459 9301 29469
rect 9267 29435 9301 29459
rect 9267 29391 9301 29397
rect 9267 29363 9301 29391
rect 9267 29323 9301 29325
rect 9267 29291 9301 29323
rect 9267 29221 9301 29253
rect 9267 29219 9301 29221
rect 9267 29153 9301 29181
rect 9267 29147 9301 29153
rect 9267 29085 9301 29109
rect 9267 29075 9301 29085
rect 9267 29017 9301 29037
rect 9267 29003 9301 29017
rect 9267 28949 9301 28965
rect 9267 28931 9301 28949
rect 9267 28881 9301 28893
rect 9267 28859 9301 28881
rect 9267 28813 9301 28821
rect 9267 28787 9301 28813
rect 9267 28745 9301 28749
rect 9267 28715 9301 28745
rect 9267 28643 9301 28677
rect 9725 29867 9759 29901
rect 9725 29799 9759 29829
rect 9725 29795 9759 29799
rect 9725 29731 9759 29757
rect 9725 29723 9759 29731
rect 9725 29663 9759 29685
rect 9725 29651 9759 29663
rect 9725 29595 9759 29613
rect 9725 29579 9759 29595
rect 9725 29527 9759 29541
rect 9725 29507 9759 29527
rect 9725 29459 9759 29469
rect 9725 29435 9759 29459
rect 9725 29391 9759 29397
rect 9725 29363 9759 29391
rect 9725 29323 9759 29325
rect 9725 29291 9759 29323
rect 9725 29221 9759 29253
rect 9725 29219 9759 29221
rect 9725 29153 9759 29181
rect 9725 29147 9759 29153
rect 9725 29085 9759 29109
rect 9725 29075 9759 29085
rect 9725 29017 9759 29037
rect 9725 29003 9759 29017
rect 9725 28949 9759 28965
rect 9725 28931 9759 28949
rect 9725 28881 9759 28893
rect 9725 28859 9759 28881
rect 9725 28813 9759 28821
rect 9725 28787 9759 28813
rect 9725 28745 9759 28749
rect 9725 28715 9759 28745
rect 9725 28643 9759 28677
rect 10183 29867 10217 29901
rect 10183 29799 10217 29829
rect 10183 29795 10217 29799
rect 10183 29731 10217 29757
rect 10183 29723 10217 29731
rect 10183 29663 10217 29685
rect 10183 29651 10217 29663
rect 10183 29595 10217 29613
rect 10183 29579 10217 29595
rect 10183 29527 10217 29541
rect 10183 29507 10217 29527
rect 10183 29459 10217 29469
rect 10183 29435 10217 29459
rect 10183 29391 10217 29397
rect 10183 29363 10217 29391
rect 10183 29323 10217 29325
rect 10183 29291 10217 29323
rect 10183 29221 10217 29253
rect 10183 29219 10217 29221
rect 10183 29153 10217 29181
rect 10183 29147 10217 29153
rect 10183 29085 10217 29109
rect 10183 29075 10217 29085
rect 10183 29017 10217 29037
rect 10183 29003 10217 29017
rect 10183 28949 10217 28965
rect 10183 28931 10217 28949
rect 10183 28881 10217 28893
rect 10183 28859 10217 28881
rect 10183 28813 10217 28821
rect 10183 28787 10217 28813
rect 10183 28745 10217 28749
rect 10183 28715 10217 28745
rect 10183 28643 10217 28677
rect 10641 29867 10675 29901
rect 10641 29799 10675 29829
rect 10641 29795 10675 29799
rect 10641 29731 10675 29757
rect 10641 29723 10675 29731
rect 10641 29663 10675 29685
rect 10641 29651 10675 29663
rect 10641 29595 10675 29613
rect 10641 29579 10675 29595
rect 10641 29527 10675 29541
rect 10641 29507 10675 29527
rect 10641 29459 10675 29469
rect 10641 29435 10675 29459
rect 10641 29391 10675 29397
rect 10641 29363 10675 29391
rect 10641 29323 10675 29325
rect 10641 29291 10675 29323
rect 10641 29221 10675 29253
rect 10641 29219 10675 29221
rect 10641 29153 10675 29181
rect 10641 29147 10675 29153
rect 10641 29085 10675 29109
rect 10641 29075 10675 29085
rect 10641 29017 10675 29037
rect 10641 29003 10675 29017
rect 10641 28949 10675 28965
rect 10641 28931 10675 28949
rect 10641 28881 10675 28893
rect 10641 28859 10675 28881
rect 10641 28813 10675 28821
rect 10641 28787 10675 28813
rect 10641 28745 10675 28749
rect 10641 28715 10675 28745
rect 10641 28643 10675 28677
rect 11099 29867 11133 29901
rect 11099 29799 11133 29829
rect 11099 29795 11133 29799
rect 11099 29731 11133 29757
rect 11099 29723 11133 29731
rect 11099 29663 11133 29685
rect 11099 29651 11133 29663
rect 11099 29595 11133 29613
rect 11099 29579 11133 29595
rect 11099 29527 11133 29541
rect 11099 29507 11133 29527
rect 11099 29459 11133 29469
rect 11099 29435 11133 29459
rect 11099 29391 11133 29397
rect 11099 29363 11133 29391
rect 11099 29323 11133 29325
rect 11099 29291 11133 29323
rect 11099 29221 11133 29253
rect 11099 29219 11133 29221
rect 11099 29153 11133 29181
rect 11099 29147 11133 29153
rect 11099 29085 11133 29109
rect 11099 29075 11133 29085
rect 11099 29017 11133 29037
rect 11099 29003 11133 29017
rect 11099 28949 11133 28965
rect 11099 28931 11133 28949
rect 11099 28881 11133 28893
rect 11099 28859 11133 28881
rect 11099 28813 11133 28821
rect 11099 28787 11133 28813
rect 11099 28745 11133 28749
rect 11099 28715 11133 28745
rect 11099 28643 11133 28677
rect 11557 29867 11591 29901
rect 11557 29799 11591 29829
rect 11557 29795 11591 29799
rect 11557 29731 11591 29757
rect 11557 29723 11591 29731
rect 11557 29663 11591 29685
rect 11557 29651 11591 29663
rect 11557 29595 11591 29613
rect 11557 29579 11591 29595
rect 11557 29527 11591 29541
rect 11557 29507 11591 29527
rect 11557 29459 11591 29469
rect 11557 29435 11591 29459
rect 11557 29391 11591 29397
rect 11557 29363 11591 29391
rect 11557 29323 11591 29325
rect 11557 29291 11591 29323
rect 11557 29221 11591 29253
rect 11557 29219 11591 29221
rect 11557 29153 11591 29181
rect 11557 29147 11591 29153
rect 11557 29085 11591 29109
rect 11557 29075 11591 29085
rect 11557 29017 11591 29037
rect 11557 29003 11591 29017
rect 11557 28949 11591 28965
rect 11557 28931 11591 28949
rect 11557 28881 11591 28893
rect 11557 28859 11591 28881
rect 11557 28813 11591 28821
rect 11557 28787 11591 28813
rect 11557 28745 11591 28749
rect 11557 28715 11591 28745
rect 11557 28643 11591 28677
rect 12015 29867 12049 29901
rect 12015 29799 12049 29829
rect 12015 29795 12049 29799
rect 12015 29731 12049 29757
rect 12015 29723 12049 29731
rect 12015 29663 12049 29685
rect 12015 29651 12049 29663
rect 12015 29595 12049 29613
rect 12015 29579 12049 29595
rect 12015 29527 12049 29541
rect 12015 29507 12049 29527
rect 12015 29459 12049 29469
rect 12015 29435 12049 29459
rect 12015 29391 12049 29397
rect 12015 29363 12049 29391
rect 12015 29323 12049 29325
rect 12015 29291 12049 29323
rect 12015 29221 12049 29253
rect 12015 29219 12049 29221
rect 12015 29153 12049 29181
rect 12015 29147 12049 29153
rect 12015 29085 12049 29109
rect 12015 29075 12049 29085
rect 12015 29017 12049 29037
rect 12015 29003 12049 29017
rect 12015 28949 12049 28965
rect 12015 28931 12049 28949
rect 12015 28881 12049 28893
rect 12015 28859 12049 28881
rect 12015 28813 12049 28821
rect 12015 28787 12049 28813
rect 12015 28745 12049 28749
rect 12015 28715 12049 28745
rect 12015 28643 12049 28677
rect 12473 29867 12507 29901
rect 12473 29799 12507 29829
rect 12473 29795 12507 29799
rect 12473 29731 12507 29757
rect 12473 29723 12507 29731
rect 12473 29663 12507 29685
rect 12473 29651 12507 29663
rect 12473 29595 12507 29613
rect 12473 29579 12507 29595
rect 12473 29527 12507 29541
rect 12473 29507 12507 29527
rect 12473 29459 12507 29469
rect 12473 29435 12507 29459
rect 12473 29391 12507 29397
rect 12473 29363 12507 29391
rect 12473 29323 12507 29325
rect 12473 29291 12507 29323
rect 12473 29221 12507 29253
rect 12473 29219 12507 29221
rect 12473 29153 12507 29181
rect 12473 29147 12507 29153
rect 12473 29085 12507 29109
rect 12473 29075 12507 29085
rect 12473 29017 12507 29037
rect 12473 29003 12507 29017
rect 12473 28949 12507 28965
rect 12473 28931 12507 28949
rect 12473 28881 12507 28893
rect 12473 28859 12507 28881
rect 12473 28813 12507 28821
rect 12473 28787 12507 28813
rect 12473 28745 12507 28749
rect 12473 28715 12507 28745
rect 12473 28643 12507 28677
rect 12931 29867 12965 29901
rect 12931 29799 12965 29829
rect 12931 29795 12965 29799
rect 12931 29731 12965 29757
rect 12931 29723 12965 29731
rect 12931 29663 12965 29685
rect 12931 29651 12965 29663
rect 12931 29595 12965 29613
rect 12931 29579 12965 29595
rect 12931 29527 12965 29541
rect 12931 29507 12965 29527
rect 12931 29459 12965 29469
rect 12931 29435 12965 29459
rect 12931 29391 12965 29397
rect 12931 29363 12965 29391
rect 12931 29323 12965 29325
rect 12931 29291 12965 29323
rect 12931 29221 12965 29253
rect 12931 29219 12965 29221
rect 12931 29153 12965 29181
rect 12931 29147 12965 29153
rect 12931 29085 12965 29109
rect 12931 29075 12965 29085
rect 12931 29017 12965 29037
rect 12931 29003 12965 29017
rect 12931 28949 12965 28965
rect 12931 28931 12965 28949
rect 12931 28881 12965 28893
rect 12931 28859 12965 28881
rect 12931 28813 12965 28821
rect 12931 28787 12965 28813
rect 12931 28745 12965 28749
rect 12931 28715 12965 28745
rect 12931 28643 12965 28677
rect 13389 29867 13423 29901
rect 13389 29799 13423 29829
rect 13389 29795 13423 29799
rect 13389 29731 13423 29757
rect 13389 29723 13423 29731
rect 13389 29663 13423 29685
rect 13389 29651 13423 29663
rect 13389 29595 13423 29613
rect 13389 29579 13423 29595
rect 13389 29527 13423 29541
rect 13389 29507 13423 29527
rect 13389 29459 13423 29469
rect 13389 29435 13423 29459
rect 13389 29391 13423 29397
rect 13389 29363 13423 29391
rect 13389 29323 13423 29325
rect 13389 29291 13423 29323
rect 13389 29221 13423 29253
rect 13389 29219 13423 29221
rect 13389 29153 13423 29181
rect 13389 29147 13423 29153
rect 13389 29085 13423 29109
rect 13389 29075 13423 29085
rect 13389 29017 13423 29037
rect 13389 29003 13423 29017
rect 13389 28949 13423 28965
rect 13389 28931 13423 28949
rect 13389 28881 13423 28893
rect 13389 28859 13423 28881
rect 13389 28813 13423 28821
rect 13389 28787 13423 28813
rect 13389 28745 13423 28749
rect 13389 28715 13423 28745
rect 13389 28643 13423 28677
rect 13847 29867 13881 29901
rect 13847 29799 13881 29829
rect 13847 29795 13881 29799
rect 13847 29731 13881 29757
rect 13847 29723 13881 29731
rect 13847 29663 13881 29685
rect 13847 29651 13881 29663
rect 13847 29595 13881 29613
rect 13847 29579 13881 29595
rect 13847 29527 13881 29541
rect 13847 29507 13881 29527
rect 13847 29459 13881 29469
rect 13847 29435 13881 29459
rect 13847 29391 13881 29397
rect 13847 29363 13881 29391
rect 13847 29323 13881 29325
rect 13847 29291 13881 29323
rect 13847 29221 13881 29253
rect 13847 29219 13881 29221
rect 13847 29153 13881 29181
rect 13847 29147 13881 29153
rect 13847 29085 13881 29109
rect 13847 29075 13881 29085
rect 13847 29017 13881 29037
rect 13847 29003 13881 29017
rect 13847 28949 13881 28965
rect 13847 28931 13881 28949
rect 13847 28881 13881 28893
rect 13847 28859 13881 28881
rect 13847 28813 13881 28821
rect 13847 28787 13881 28813
rect 13847 28745 13881 28749
rect 13847 28715 13881 28745
rect 13847 28643 13881 28677
rect 14305 29867 14339 29901
rect 14305 29799 14339 29829
rect 14305 29795 14339 29799
rect 14305 29731 14339 29757
rect 14305 29723 14339 29731
rect 14305 29663 14339 29685
rect 14305 29651 14339 29663
rect 14305 29595 14339 29613
rect 14305 29579 14339 29595
rect 14305 29527 14339 29541
rect 14305 29507 14339 29527
rect 14305 29459 14339 29469
rect 14305 29435 14339 29459
rect 14305 29391 14339 29397
rect 14305 29363 14339 29391
rect 14305 29323 14339 29325
rect 14305 29291 14339 29323
rect 14305 29221 14339 29253
rect 14305 29219 14339 29221
rect 14305 29153 14339 29181
rect 14305 29147 14339 29153
rect 14305 29085 14339 29109
rect 14305 29075 14339 29085
rect 14305 29017 14339 29037
rect 14305 29003 14339 29017
rect 14305 28949 14339 28965
rect 14305 28931 14339 28949
rect 14305 28881 14339 28893
rect 14305 28859 14339 28881
rect 14305 28813 14339 28821
rect 14305 28787 14339 28813
rect 14305 28745 14339 28749
rect 14305 28715 14339 28745
rect 14305 28643 14339 28677
rect 14763 29867 14797 29901
rect 14763 29799 14797 29829
rect 14763 29795 14797 29799
rect 14763 29731 14797 29757
rect 14763 29723 14797 29731
rect 14763 29663 14797 29685
rect 14763 29651 14797 29663
rect 14763 29595 14797 29613
rect 14763 29579 14797 29595
rect 14763 29527 14797 29541
rect 14763 29507 14797 29527
rect 14763 29459 14797 29469
rect 14763 29435 14797 29459
rect 14763 29391 14797 29397
rect 14763 29363 14797 29391
rect 14763 29323 14797 29325
rect 14763 29291 14797 29323
rect 14763 29221 14797 29253
rect 14763 29219 14797 29221
rect 14763 29153 14797 29181
rect 14763 29147 14797 29153
rect 14763 29085 14797 29109
rect 14763 29075 14797 29085
rect 14763 29017 14797 29037
rect 14763 29003 14797 29017
rect 14763 28949 14797 28965
rect 14763 28931 14797 28949
rect 14763 28881 14797 28893
rect 14763 28859 14797 28881
rect 14763 28813 14797 28821
rect 14763 28787 14797 28813
rect 14763 28745 14797 28749
rect 14763 28715 14797 28745
rect 14763 28643 14797 28677
rect 15221 29867 15255 29901
rect 15221 29799 15255 29829
rect 15221 29795 15255 29799
rect 15221 29731 15255 29757
rect 15221 29723 15255 29731
rect 15221 29663 15255 29685
rect 15221 29651 15255 29663
rect 15221 29595 15255 29613
rect 15221 29579 15255 29595
rect 15221 29527 15255 29541
rect 15221 29507 15255 29527
rect 15221 29459 15255 29469
rect 15221 29435 15255 29459
rect 15221 29391 15255 29397
rect 15221 29363 15255 29391
rect 15221 29323 15255 29325
rect 15221 29291 15255 29323
rect 15221 29221 15255 29253
rect 15221 29219 15255 29221
rect 15221 29153 15255 29181
rect 15221 29147 15255 29153
rect 15221 29085 15255 29109
rect 15221 29075 15255 29085
rect 15221 29017 15255 29037
rect 15221 29003 15255 29017
rect 15221 28949 15255 28965
rect 15221 28931 15255 28949
rect 15221 28881 15255 28893
rect 15221 28859 15255 28881
rect 15221 28813 15255 28821
rect 15221 28787 15255 28813
rect 15221 28745 15255 28749
rect 15221 28715 15255 28745
rect 15221 28643 15255 28677
rect 15679 29867 15713 29901
rect 15679 29799 15713 29829
rect 15679 29795 15713 29799
rect 15679 29731 15713 29757
rect 15679 29723 15713 29731
rect 15679 29663 15713 29685
rect 15679 29651 15713 29663
rect 15679 29595 15713 29613
rect 15679 29579 15713 29595
rect 15679 29527 15713 29541
rect 15679 29507 15713 29527
rect 15679 29459 15713 29469
rect 15679 29435 15713 29459
rect 15679 29391 15713 29397
rect 15679 29363 15713 29391
rect 15679 29323 15713 29325
rect 15679 29291 15713 29323
rect 15679 29221 15713 29253
rect 15679 29219 15713 29221
rect 15679 29153 15713 29181
rect 15679 29147 15713 29153
rect 15679 29085 15713 29109
rect 15679 29075 15713 29085
rect 15679 29017 15713 29037
rect 15679 29003 15713 29017
rect 15679 28949 15713 28965
rect 15679 28931 15713 28949
rect 15679 28881 15713 28893
rect 15679 28859 15713 28881
rect 15679 28813 15713 28821
rect 15679 28787 15713 28813
rect 15679 28745 15713 28749
rect 15679 28715 15713 28745
rect 15679 28643 15713 28677
rect 16137 29867 16171 29901
rect 16137 29799 16171 29829
rect 16137 29795 16171 29799
rect 16137 29731 16171 29757
rect 16137 29723 16171 29731
rect 16137 29663 16171 29685
rect 16137 29651 16171 29663
rect 16137 29595 16171 29613
rect 16137 29579 16171 29595
rect 16137 29527 16171 29541
rect 16137 29507 16171 29527
rect 16137 29459 16171 29469
rect 16137 29435 16171 29459
rect 16137 29391 16171 29397
rect 16137 29363 16171 29391
rect 16137 29323 16171 29325
rect 16137 29291 16171 29323
rect 16137 29221 16171 29253
rect 16137 29219 16171 29221
rect 16137 29153 16171 29181
rect 16137 29147 16171 29153
rect 16137 29085 16171 29109
rect 16137 29075 16171 29085
rect 16137 29017 16171 29037
rect 16137 29003 16171 29017
rect 16137 28949 16171 28965
rect 16137 28931 16171 28949
rect 16137 28881 16171 28893
rect 16137 28859 16171 28881
rect 16137 28813 16171 28821
rect 16137 28787 16171 28813
rect 16137 28745 16171 28749
rect 16137 28715 16171 28745
rect 16137 28643 16171 28677
rect 16595 29867 16629 29901
rect 16595 29799 16629 29829
rect 16595 29795 16629 29799
rect 16595 29731 16629 29757
rect 16595 29723 16629 29731
rect 16595 29663 16629 29685
rect 16595 29651 16629 29663
rect 16595 29595 16629 29613
rect 16595 29579 16629 29595
rect 16595 29527 16629 29541
rect 16595 29507 16629 29527
rect 16595 29459 16629 29469
rect 16595 29435 16629 29459
rect 16595 29391 16629 29397
rect 16595 29363 16629 29391
rect 16595 29323 16629 29325
rect 16595 29291 16629 29323
rect 16595 29221 16629 29253
rect 16595 29219 16629 29221
rect 16595 29153 16629 29181
rect 16595 29147 16629 29153
rect 16595 29085 16629 29109
rect 16595 29075 16629 29085
rect 16595 29017 16629 29037
rect 16595 29003 16629 29017
rect 16595 28949 16629 28965
rect 16595 28931 16629 28949
rect 16595 28881 16629 28893
rect 16595 28859 16629 28881
rect 16595 28813 16629 28821
rect 16595 28787 16629 28813
rect 16595 28745 16629 28749
rect 16595 28715 16629 28745
rect 16595 28643 16629 28677
rect 17053 29867 17087 29901
rect 17053 29799 17087 29829
rect 17053 29795 17087 29799
rect 17053 29731 17087 29757
rect 17053 29723 17087 29731
rect 17053 29663 17087 29685
rect 17053 29651 17087 29663
rect 17053 29595 17087 29613
rect 17053 29579 17087 29595
rect 17053 29527 17087 29541
rect 17053 29507 17087 29527
rect 17053 29459 17087 29469
rect 17053 29435 17087 29459
rect 17053 29391 17087 29397
rect 17053 29363 17087 29391
rect 17053 29323 17087 29325
rect 17053 29291 17087 29323
rect 17053 29221 17087 29253
rect 17053 29219 17087 29221
rect 17053 29153 17087 29181
rect 17053 29147 17087 29153
rect 17053 29085 17087 29109
rect 17053 29075 17087 29085
rect 17053 29017 17087 29037
rect 17053 29003 17087 29017
rect 17053 28949 17087 28965
rect 17053 28931 17087 28949
rect 17053 28881 17087 28893
rect 17053 28859 17087 28881
rect 17053 28813 17087 28821
rect 17053 28787 17087 28813
rect 17053 28745 17087 28749
rect 17053 28715 17087 28745
rect 17053 28643 17087 28677
rect 17511 29867 17545 29901
rect 17511 29799 17545 29829
rect 17511 29795 17545 29799
rect 17511 29731 17545 29757
rect 17511 29723 17545 29731
rect 17511 29663 17545 29685
rect 17511 29651 17545 29663
rect 17511 29595 17545 29613
rect 17511 29579 17545 29595
rect 17511 29527 17545 29541
rect 17511 29507 17545 29527
rect 17511 29459 17545 29469
rect 17511 29435 17545 29459
rect 17511 29391 17545 29397
rect 17511 29363 17545 29391
rect 17511 29323 17545 29325
rect 17511 29291 17545 29323
rect 17511 29221 17545 29253
rect 17511 29219 17545 29221
rect 17511 29153 17545 29181
rect 17511 29147 17545 29153
rect 17511 29085 17545 29109
rect 17511 29075 17545 29085
rect 17511 29017 17545 29037
rect 17511 29003 17545 29017
rect 17511 28949 17545 28965
rect 17511 28931 17545 28949
rect 17511 28881 17545 28893
rect 17511 28859 17545 28881
rect 17511 28813 17545 28821
rect 17511 28787 17545 28813
rect 17511 28745 17545 28749
rect 17511 28715 17545 28745
rect 17511 28643 17545 28677
rect 17969 29867 18003 29901
rect 17969 29799 18003 29829
rect 17969 29795 18003 29799
rect 17969 29731 18003 29757
rect 17969 29723 18003 29731
rect 17969 29663 18003 29685
rect 17969 29651 18003 29663
rect 17969 29595 18003 29613
rect 17969 29579 18003 29595
rect 17969 29527 18003 29541
rect 17969 29507 18003 29527
rect 17969 29459 18003 29469
rect 17969 29435 18003 29459
rect 17969 29391 18003 29397
rect 17969 29363 18003 29391
rect 17969 29323 18003 29325
rect 17969 29291 18003 29323
rect 17969 29221 18003 29253
rect 17969 29219 18003 29221
rect 17969 29153 18003 29181
rect 17969 29147 18003 29153
rect 17969 29085 18003 29109
rect 17969 29075 18003 29085
rect 17969 29017 18003 29037
rect 17969 29003 18003 29017
rect 17969 28949 18003 28965
rect 17969 28931 18003 28949
rect 17969 28881 18003 28893
rect 17969 28859 18003 28881
rect 17969 28813 18003 28821
rect 17969 28787 18003 28813
rect 17969 28745 18003 28749
rect 17969 28715 18003 28745
rect 17969 28643 18003 28677
rect 18427 29867 18461 29901
rect 18427 29799 18461 29829
rect 18427 29795 18461 29799
rect 18427 29731 18461 29757
rect 18427 29723 18461 29731
rect 18427 29663 18461 29685
rect 18427 29651 18461 29663
rect 18427 29595 18461 29613
rect 18427 29579 18461 29595
rect 18427 29527 18461 29541
rect 18427 29507 18461 29527
rect 18427 29459 18461 29469
rect 18427 29435 18461 29459
rect 18427 29391 18461 29397
rect 18427 29363 18461 29391
rect 18427 29323 18461 29325
rect 18427 29291 18461 29323
rect 18427 29221 18461 29253
rect 18427 29219 18461 29221
rect 18427 29153 18461 29181
rect 18427 29147 18461 29153
rect 18427 29085 18461 29109
rect 18427 29075 18461 29085
rect 18427 29017 18461 29037
rect 18427 29003 18461 29017
rect 18427 28949 18461 28965
rect 18427 28931 18461 28949
rect 18427 28881 18461 28893
rect 18427 28859 18461 28881
rect 18427 28813 18461 28821
rect 18427 28787 18461 28813
rect 18427 28745 18461 28749
rect 18427 28715 18461 28745
rect 18427 28643 18461 28677
rect 18885 29867 18919 29901
rect 18885 29799 18919 29829
rect 18885 29795 18919 29799
rect 18885 29731 18919 29757
rect 18885 29723 18919 29731
rect 18885 29663 18919 29685
rect 18885 29651 18919 29663
rect 18885 29595 18919 29613
rect 18885 29579 18919 29595
rect 18885 29527 18919 29541
rect 18885 29507 18919 29527
rect 18885 29459 18919 29469
rect 18885 29435 18919 29459
rect 18885 29391 18919 29397
rect 18885 29363 18919 29391
rect 18885 29323 18919 29325
rect 18885 29291 18919 29323
rect 18885 29221 18919 29253
rect 18885 29219 18919 29221
rect 18885 29153 18919 29181
rect 18885 29147 18919 29153
rect 18885 29085 18919 29109
rect 18885 29075 18919 29085
rect 18885 29017 18919 29037
rect 18885 29003 18919 29017
rect 18885 28949 18919 28965
rect 18885 28931 18919 28949
rect 18885 28881 18919 28893
rect 18885 28859 18919 28881
rect 18885 28813 18919 28821
rect 18885 28787 18919 28813
rect 18885 28745 18919 28749
rect 18885 28715 18919 28745
rect 18885 28643 18919 28677
rect 19343 29867 19377 29901
rect 19343 29799 19377 29829
rect 19343 29795 19377 29799
rect 19343 29731 19377 29757
rect 19343 29723 19377 29731
rect 19343 29663 19377 29685
rect 19343 29651 19377 29663
rect 19343 29595 19377 29613
rect 19343 29579 19377 29595
rect 19343 29527 19377 29541
rect 19343 29507 19377 29527
rect 19343 29459 19377 29469
rect 19343 29435 19377 29459
rect 19343 29391 19377 29397
rect 19343 29363 19377 29391
rect 19343 29323 19377 29325
rect 19343 29291 19377 29323
rect 19343 29221 19377 29253
rect 19343 29219 19377 29221
rect 19343 29153 19377 29181
rect 19343 29147 19377 29153
rect 19343 29085 19377 29109
rect 19343 29075 19377 29085
rect 19343 29017 19377 29037
rect 19343 29003 19377 29017
rect 19343 28949 19377 28965
rect 19343 28931 19377 28949
rect 19343 28881 19377 28893
rect 19343 28859 19377 28881
rect 19343 28813 19377 28821
rect 19343 28787 19377 28813
rect 19343 28745 19377 28749
rect 19343 28715 19377 28745
rect 19343 28643 19377 28677
rect 19801 29867 19835 29901
rect 19801 29799 19835 29829
rect 19801 29795 19835 29799
rect 19801 29731 19835 29757
rect 19801 29723 19835 29731
rect 19801 29663 19835 29685
rect 19801 29651 19835 29663
rect 19801 29595 19835 29613
rect 19801 29579 19835 29595
rect 19801 29527 19835 29541
rect 19801 29507 19835 29527
rect 19801 29459 19835 29469
rect 19801 29435 19835 29459
rect 19801 29391 19835 29397
rect 19801 29363 19835 29391
rect 19801 29323 19835 29325
rect 19801 29291 19835 29323
rect 19801 29221 19835 29253
rect 19801 29219 19835 29221
rect 19801 29153 19835 29181
rect 19801 29147 19835 29153
rect 19801 29085 19835 29109
rect 19801 29075 19835 29085
rect 19801 29017 19835 29037
rect 19801 29003 19835 29017
rect 19801 28949 19835 28965
rect 19801 28931 19835 28949
rect 19801 28881 19835 28893
rect 19801 28859 19835 28881
rect 19801 28813 19835 28821
rect 19801 28787 19835 28813
rect 19801 28745 19835 28749
rect 19801 28715 19835 28745
rect 19801 28643 19835 28677
rect 20259 29867 20293 29901
rect 20259 29799 20293 29829
rect 20259 29795 20293 29799
rect 20259 29731 20293 29757
rect 20259 29723 20293 29731
rect 20259 29663 20293 29685
rect 20259 29651 20293 29663
rect 20259 29595 20293 29613
rect 20259 29579 20293 29595
rect 20259 29527 20293 29541
rect 20259 29507 20293 29527
rect 20259 29459 20293 29469
rect 20259 29435 20293 29459
rect 20259 29391 20293 29397
rect 20259 29363 20293 29391
rect 20259 29323 20293 29325
rect 20259 29291 20293 29323
rect 20259 29221 20293 29253
rect 20259 29219 20293 29221
rect 20259 29153 20293 29181
rect 20259 29147 20293 29153
rect 20259 29085 20293 29109
rect 20259 29075 20293 29085
rect 20259 29017 20293 29037
rect 20259 29003 20293 29017
rect 20259 28949 20293 28965
rect 20259 28931 20293 28949
rect 20259 28881 20293 28893
rect 20259 28859 20293 28881
rect 20259 28813 20293 28821
rect 20259 28787 20293 28813
rect 20259 28745 20293 28749
rect 20259 28715 20293 28745
rect 20259 28643 20293 28677
rect 20717 29867 20751 29901
rect 20717 29799 20751 29829
rect 20717 29795 20751 29799
rect 20717 29731 20751 29757
rect 20717 29723 20751 29731
rect 20717 29663 20751 29685
rect 20717 29651 20751 29663
rect 20717 29595 20751 29613
rect 20717 29579 20751 29595
rect 20717 29527 20751 29541
rect 20717 29507 20751 29527
rect 20717 29459 20751 29469
rect 20717 29435 20751 29459
rect 20717 29391 20751 29397
rect 20717 29363 20751 29391
rect 20717 29323 20751 29325
rect 20717 29291 20751 29323
rect 20717 29221 20751 29253
rect 20717 29219 20751 29221
rect 20717 29153 20751 29181
rect 20717 29147 20751 29153
rect 20717 29085 20751 29109
rect 20717 29075 20751 29085
rect 20717 29017 20751 29037
rect 20717 29003 20751 29017
rect 20717 28949 20751 28965
rect 20717 28931 20751 28949
rect 20717 28881 20751 28893
rect 20717 28859 20751 28881
rect 20717 28813 20751 28821
rect 20717 28787 20751 28813
rect 20717 28745 20751 28749
rect 20717 28715 20751 28745
rect 20717 28643 20751 28677
rect 21175 29867 21209 29901
rect 21175 29799 21209 29829
rect 21175 29795 21209 29799
rect 21175 29731 21209 29757
rect 21175 29723 21209 29731
rect 21175 29663 21209 29685
rect 21175 29651 21209 29663
rect 21175 29595 21209 29613
rect 21175 29579 21209 29595
rect 21175 29527 21209 29541
rect 21175 29507 21209 29527
rect 21175 29459 21209 29469
rect 21175 29435 21209 29459
rect 21175 29391 21209 29397
rect 21175 29363 21209 29391
rect 21175 29323 21209 29325
rect 21175 29291 21209 29323
rect 21175 29221 21209 29253
rect 21175 29219 21209 29221
rect 21175 29153 21209 29181
rect 21175 29147 21209 29153
rect 21175 29085 21209 29109
rect 21175 29075 21209 29085
rect 21175 29017 21209 29037
rect 21175 29003 21209 29017
rect 21175 28949 21209 28965
rect 21175 28931 21209 28949
rect 21175 28881 21209 28893
rect 21175 28859 21209 28881
rect 21175 28813 21209 28821
rect 21175 28787 21209 28813
rect 21175 28745 21209 28749
rect 21175 28715 21209 28745
rect 21175 28643 21209 28677
rect 21633 29867 21667 29901
rect 21633 29799 21667 29829
rect 21633 29795 21667 29799
rect 21633 29731 21667 29757
rect 21633 29723 21667 29731
rect 21633 29663 21667 29685
rect 21633 29651 21667 29663
rect 21633 29595 21667 29613
rect 21633 29579 21667 29595
rect 21633 29527 21667 29541
rect 21633 29507 21667 29527
rect 21633 29459 21667 29469
rect 21633 29435 21667 29459
rect 21633 29391 21667 29397
rect 21633 29363 21667 29391
rect 21633 29323 21667 29325
rect 21633 29291 21667 29323
rect 21633 29221 21667 29253
rect 21633 29219 21667 29221
rect 21633 29153 21667 29181
rect 21633 29147 21667 29153
rect 21633 29085 21667 29109
rect 21633 29075 21667 29085
rect 21633 29017 21667 29037
rect 21633 29003 21667 29017
rect 21633 28949 21667 28965
rect 21633 28931 21667 28949
rect 21633 28881 21667 28893
rect 21633 28859 21667 28881
rect 21633 28813 21667 28821
rect 21633 28787 21667 28813
rect 21633 28745 21667 28749
rect 21633 28715 21667 28745
rect 21633 28643 21667 28677
rect 22091 29867 22125 29901
rect 22091 29799 22125 29829
rect 22091 29795 22125 29799
rect 22091 29731 22125 29757
rect 22091 29723 22125 29731
rect 22091 29663 22125 29685
rect 22091 29651 22125 29663
rect 22091 29595 22125 29613
rect 22091 29579 22125 29595
rect 22091 29527 22125 29541
rect 22091 29507 22125 29527
rect 22091 29459 22125 29469
rect 22091 29435 22125 29459
rect 22091 29391 22125 29397
rect 22091 29363 22125 29391
rect 22091 29323 22125 29325
rect 22091 29291 22125 29323
rect 22091 29221 22125 29253
rect 22091 29219 22125 29221
rect 22091 29153 22125 29181
rect 22091 29147 22125 29153
rect 22091 29085 22125 29109
rect 22091 29075 22125 29085
rect 22091 29017 22125 29037
rect 22091 29003 22125 29017
rect 22091 28949 22125 28965
rect 22091 28931 22125 28949
rect 22091 28881 22125 28893
rect 22091 28859 22125 28881
rect 22091 28813 22125 28821
rect 22091 28787 22125 28813
rect 22091 28745 22125 28749
rect 22091 28715 22125 28745
rect 22091 28643 22125 28677
rect 22549 29867 22583 29901
rect 22549 29799 22583 29829
rect 22549 29795 22583 29799
rect 22549 29731 22583 29757
rect 22549 29723 22583 29731
rect 22549 29663 22583 29685
rect 22549 29651 22583 29663
rect 22549 29595 22583 29613
rect 22549 29579 22583 29595
rect 22549 29527 22583 29541
rect 22549 29507 22583 29527
rect 22549 29459 22583 29469
rect 22549 29435 22583 29459
rect 22549 29391 22583 29397
rect 22549 29363 22583 29391
rect 22549 29323 22583 29325
rect 22549 29291 22583 29323
rect 22549 29221 22583 29253
rect 22549 29219 22583 29221
rect 22549 29153 22583 29181
rect 22549 29147 22583 29153
rect 22549 29085 22583 29109
rect 22549 29075 22583 29085
rect 22549 29017 22583 29037
rect 22549 29003 22583 29017
rect 22549 28949 22583 28965
rect 22549 28931 22583 28949
rect 22549 28881 22583 28893
rect 22549 28859 22583 28881
rect 22549 28813 22583 28821
rect 22549 28787 22583 28813
rect 22549 28745 22583 28749
rect 22549 28715 22583 28745
rect 22549 28643 22583 28677
rect 23007 29867 23041 29901
rect 23007 29799 23041 29829
rect 23007 29795 23041 29799
rect 23007 29731 23041 29757
rect 23007 29723 23041 29731
rect 23007 29663 23041 29685
rect 23007 29651 23041 29663
rect 23007 29595 23041 29613
rect 23007 29579 23041 29595
rect 23007 29527 23041 29541
rect 23007 29507 23041 29527
rect 23007 29459 23041 29469
rect 23007 29435 23041 29459
rect 23007 29391 23041 29397
rect 23007 29363 23041 29391
rect 23007 29323 23041 29325
rect 23007 29291 23041 29323
rect 23007 29221 23041 29253
rect 23007 29219 23041 29221
rect 23007 29153 23041 29181
rect 23007 29147 23041 29153
rect 23007 29085 23041 29109
rect 23007 29075 23041 29085
rect 23007 29017 23041 29037
rect 23007 29003 23041 29017
rect 23007 28949 23041 28965
rect 23007 28931 23041 28949
rect 23007 28881 23041 28893
rect 23007 28859 23041 28881
rect 23007 28813 23041 28821
rect 23007 28787 23041 28813
rect 23007 28745 23041 28749
rect 23007 28715 23041 28745
rect 23007 28643 23041 28677
rect 23465 29867 23499 29901
rect 23465 29799 23499 29829
rect 23465 29795 23499 29799
rect 23465 29731 23499 29757
rect 23465 29723 23499 29731
rect 23465 29663 23499 29685
rect 23465 29651 23499 29663
rect 23465 29595 23499 29613
rect 23465 29579 23499 29595
rect 23465 29527 23499 29541
rect 23465 29507 23499 29527
rect 23465 29459 23499 29469
rect 23465 29435 23499 29459
rect 23465 29391 23499 29397
rect 23465 29363 23499 29391
rect 23465 29323 23499 29325
rect 23465 29291 23499 29323
rect 23465 29221 23499 29253
rect 23465 29219 23499 29221
rect 23465 29153 23499 29181
rect 23465 29147 23499 29153
rect 23465 29085 23499 29109
rect 23465 29075 23499 29085
rect 23465 29017 23499 29037
rect 23465 29003 23499 29017
rect 23465 28949 23499 28965
rect 23465 28931 23499 28949
rect 23465 28881 23499 28893
rect 23465 28859 23499 28881
rect 23465 28813 23499 28821
rect 23465 28787 23499 28813
rect 23465 28745 23499 28749
rect 23465 28715 23499 28745
rect 23465 28643 23499 28677
rect 23923 29867 23957 29901
rect 23923 29799 23957 29829
rect 23923 29795 23957 29799
rect 23923 29731 23957 29757
rect 23923 29723 23957 29731
rect 23923 29663 23957 29685
rect 23923 29651 23957 29663
rect 23923 29595 23957 29613
rect 23923 29579 23957 29595
rect 23923 29527 23957 29541
rect 23923 29507 23957 29527
rect 23923 29459 23957 29469
rect 23923 29435 23957 29459
rect 23923 29391 23957 29397
rect 23923 29363 23957 29391
rect 23923 29323 23957 29325
rect 23923 29291 23957 29323
rect 23923 29221 23957 29253
rect 23923 29219 23957 29221
rect 23923 29153 23957 29181
rect 23923 29147 23957 29153
rect 23923 29085 23957 29109
rect 23923 29075 23957 29085
rect 23923 29017 23957 29037
rect 23923 29003 23957 29017
rect 23923 28949 23957 28965
rect 23923 28931 23957 28949
rect 23923 28881 23957 28893
rect 23923 28859 23957 28881
rect 23923 28813 23957 28821
rect 23923 28787 23957 28813
rect 23923 28745 23957 28749
rect 23923 28715 23957 28745
rect 23923 28643 23957 28677
rect 24381 29867 24415 29901
rect 24381 29799 24415 29829
rect 24381 29795 24415 29799
rect 24381 29731 24415 29757
rect 24381 29723 24415 29731
rect 24381 29663 24415 29685
rect 24381 29651 24415 29663
rect 24381 29595 24415 29613
rect 24381 29579 24415 29595
rect 24381 29527 24415 29541
rect 24381 29507 24415 29527
rect 24381 29459 24415 29469
rect 24381 29435 24415 29459
rect 24381 29391 24415 29397
rect 24381 29363 24415 29391
rect 24381 29323 24415 29325
rect 24381 29291 24415 29323
rect 24381 29221 24415 29253
rect 24381 29219 24415 29221
rect 24381 29153 24415 29181
rect 24381 29147 24415 29153
rect 24381 29085 24415 29109
rect 24381 29075 24415 29085
rect 24381 29017 24415 29037
rect 24381 29003 24415 29017
rect 24381 28949 24415 28965
rect 24381 28931 24415 28949
rect 24381 28881 24415 28893
rect 24381 28859 24415 28881
rect 24381 28813 24415 28821
rect 24381 28787 24415 28813
rect 24381 28745 24415 28749
rect 24381 28715 24415 28745
rect 24381 28643 24415 28677
rect 24839 29867 24873 29901
rect 24839 29799 24873 29829
rect 24839 29795 24873 29799
rect 24839 29731 24873 29757
rect 24839 29723 24873 29731
rect 24839 29663 24873 29685
rect 24839 29651 24873 29663
rect 24839 29595 24873 29613
rect 24839 29579 24873 29595
rect 24839 29527 24873 29541
rect 24839 29507 24873 29527
rect 24839 29459 24873 29469
rect 24839 29435 24873 29459
rect 24839 29391 24873 29397
rect 24839 29363 24873 29391
rect 24839 29323 24873 29325
rect 24839 29291 24873 29323
rect 24839 29221 24873 29253
rect 24839 29219 24873 29221
rect 24839 29153 24873 29181
rect 24839 29147 24873 29153
rect 24839 29085 24873 29109
rect 24839 29075 24873 29085
rect 24839 29017 24873 29037
rect 24839 29003 24873 29017
rect 24839 28949 24873 28965
rect 24839 28931 24873 28949
rect 24839 28881 24873 28893
rect 24839 28859 24873 28881
rect 24839 28813 24873 28821
rect 24839 28787 24873 28813
rect 24839 28745 24873 28749
rect 24839 28715 24873 28745
rect 24839 28643 24873 28677
rect 25297 29867 25331 29901
rect 25297 29799 25331 29829
rect 25297 29795 25331 29799
rect 25297 29731 25331 29757
rect 25297 29723 25331 29731
rect 25297 29663 25331 29685
rect 25297 29651 25331 29663
rect 25297 29595 25331 29613
rect 25297 29579 25331 29595
rect 25297 29527 25331 29541
rect 25297 29507 25331 29527
rect 25297 29459 25331 29469
rect 25297 29435 25331 29459
rect 25297 29391 25331 29397
rect 25297 29363 25331 29391
rect 25297 29323 25331 29325
rect 25297 29291 25331 29323
rect 25297 29221 25331 29253
rect 25297 29219 25331 29221
rect 25297 29153 25331 29181
rect 25297 29147 25331 29153
rect 25297 29085 25331 29109
rect 25297 29075 25331 29085
rect 25297 29017 25331 29037
rect 25297 29003 25331 29017
rect 25297 28949 25331 28965
rect 25297 28931 25331 28949
rect 25297 28881 25331 28893
rect 25297 28859 25331 28881
rect 25297 28813 25331 28821
rect 25297 28787 25331 28813
rect 25297 28745 25331 28749
rect 25297 28715 25331 28745
rect 25297 28643 25331 28677
rect 25755 29867 25789 29901
rect 25755 29799 25789 29829
rect 25755 29795 25789 29799
rect 25755 29731 25789 29757
rect 25755 29723 25789 29731
rect 25755 29663 25789 29685
rect 25755 29651 25789 29663
rect 25755 29595 25789 29613
rect 25755 29579 25789 29595
rect 25755 29527 25789 29541
rect 25755 29507 25789 29527
rect 25755 29459 25789 29469
rect 25755 29435 25789 29459
rect 25755 29391 25789 29397
rect 25755 29363 25789 29391
rect 25755 29323 25789 29325
rect 25755 29291 25789 29323
rect 25755 29221 25789 29253
rect 25755 29219 25789 29221
rect 25755 29153 25789 29181
rect 25755 29147 25789 29153
rect 25755 29085 25789 29109
rect 25755 29075 25789 29085
rect 25755 29017 25789 29037
rect 25755 29003 25789 29017
rect 25755 28949 25789 28965
rect 25755 28931 25789 28949
rect 25755 28881 25789 28893
rect 25755 28859 25789 28881
rect 25755 28813 25789 28821
rect 25755 28787 25789 28813
rect 25755 28745 25789 28749
rect 25755 28715 25789 28745
rect 25755 28643 25789 28677
rect 26213 29867 26247 29901
rect 26213 29799 26247 29829
rect 26213 29795 26247 29799
rect 26213 29731 26247 29757
rect 26213 29723 26247 29731
rect 26213 29663 26247 29685
rect 26213 29651 26247 29663
rect 26213 29595 26247 29613
rect 26213 29579 26247 29595
rect 26213 29527 26247 29541
rect 26213 29507 26247 29527
rect 26213 29459 26247 29469
rect 26213 29435 26247 29459
rect 26213 29391 26247 29397
rect 26213 29363 26247 29391
rect 26213 29323 26247 29325
rect 26213 29291 26247 29323
rect 26213 29221 26247 29253
rect 26213 29219 26247 29221
rect 26213 29153 26247 29181
rect 26213 29147 26247 29153
rect 26213 29085 26247 29109
rect 26213 29075 26247 29085
rect 26213 29017 26247 29037
rect 26213 29003 26247 29017
rect 26213 28949 26247 28965
rect 26213 28931 26247 28949
rect 26213 28881 26247 28893
rect 26213 28859 26247 28881
rect 26213 28813 26247 28821
rect 26213 28787 26247 28813
rect 26213 28745 26247 28749
rect 26213 28715 26247 28745
rect 26213 28643 26247 28677
rect 26671 29867 26705 29901
rect 26671 29799 26705 29829
rect 26671 29795 26705 29799
rect 26671 29731 26705 29757
rect 26671 29723 26705 29731
rect 26671 29663 26705 29685
rect 26671 29651 26705 29663
rect 26671 29595 26705 29613
rect 26671 29579 26705 29595
rect 26671 29527 26705 29541
rect 26671 29507 26705 29527
rect 26671 29459 26705 29469
rect 26671 29435 26705 29459
rect 26671 29391 26705 29397
rect 26671 29363 26705 29391
rect 26671 29323 26705 29325
rect 26671 29291 26705 29323
rect 26671 29221 26705 29253
rect 26671 29219 26705 29221
rect 26671 29153 26705 29181
rect 26671 29147 26705 29153
rect 26671 29085 26705 29109
rect 26671 29075 26705 29085
rect 26671 29017 26705 29037
rect 26671 29003 26705 29017
rect 26671 28949 26705 28965
rect 26671 28931 26705 28949
rect 26671 28881 26705 28893
rect 26671 28859 26705 28881
rect 26671 28813 26705 28821
rect 26671 28787 26705 28813
rect 26671 28745 26705 28749
rect 26671 28715 26705 28745
rect 26671 28643 26705 28677
rect 27129 29867 27163 29901
rect 27129 29799 27163 29829
rect 27129 29795 27163 29799
rect 27129 29731 27163 29757
rect 27129 29723 27163 29731
rect 27129 29663 27163 29685
rect 27129 29651 27163 29663
rect 27129 29595 27163 29613
rect 27129 29579 27163 29595
rect 27129 29527 27163 29541
rect 27129 29507 27163 29527
rect 27129 29459 27163 29469
rect 27129 29435 27163 29459
rect 27129 29391 27163 29397
rect 27129 29363 27163 29391
rect 27129 29323 27163 29325
rect 27129 29291 27163 29323
rect 27129 29221 27163 29253
rect 27129 29219 27163 29221
rect 27129 29153 27163 29181
rect 27129 29147 27163 29153
rect 27129 29085 27163 29109
rect 27129 29075 27163 29085
rect 27129 29017 27163 29037
rect 27129 29003 27163 29017
rect 27129 28949 27163 28965
rect 27129 28931 27163 28949
rect 27129 28881 27163 28893
rect 27129 28859 27163 28881
rect 27129 28813 27163 28821
rect 27129 28787 27163 28813
rect 27129 28745 27163 28749
rect 27129 28715 27163 28745
rect 27129 28643 27163 28677
rect 27587 29867 27621 29901
rect 27587 29799 27621 29829
rect 27587 29795 27621 29799
rect 27587 29731 27621 29757
rect 27587 29723 27621 29731
rect 27587 29663 27621 29685
rect 27587 29651 27621 29663
rect 27587 29595 27621 29613
rect 27587 29579 27621 29595
rect 27587 29527 27621 29541
rect 27587 29507 27621 29527
rect 27587 29459 27621 29469
rect 27587 29435 27621 29459
rect 27587 29391 27621 29397
rect 27587 29363 27621 29391
rect 27587 29323 27621 29325
rect 27587 29291 27621 29323
rect 27587 29221 27621 29253
rect 27587 29219 27621 29221
rect 27587 29153 27621 29181
rect 27587 29147 27621 29153
rect 27587 29085 27621 29109
rect 27587 29075 27621 29085
rect 27587 29017 27621 29037
rect 27587 29003 27621 29017
rect 27587 28949 27621 28965
rect 27587 28931 27621 28949
rect 27587 28881 27621 28893
rect 27587 28859 27621 28881
rect 27587 28813 27621 28821
rect 27587 28787 27621 28813
rect 27587 28745 27621 28749
rect 27587 28715 27621 28745
rect 27587 28643 27621 28677
rect 28045 29867 28079 29901
rect 28045 29799 28079 29829
rect 28045 29795 28079 29799
rect 28045 29731 28079 29757
rect 28045 29723 28079 29731
rect 28045 29663 28079 29685
rect 28045 29651 28079 29663
rect 28045 29595 28079 29613
rect 28045 29579 28079 29595
rect 28045 29527 28079 29541
rect 28045 29507 28079 29527
rect 28045 29459 28079 29469
rect 28045 29435 28079 29459
rect 28045 29391 28079 29397
rect 28045 29363 28079 29391
rect 28045 29323 28079 29325
rect 28045 29291 28079 29323
rect 28045 29221 28079 29253
rect 28045 29219 28079 29221
rect 28045 29153 28079 29181
rect 28045 29147 28079 29153
rect 28045 29085 28079 29109
rect 28045 29075 28079 29085
rect 28045 29017 28079 29037
rect 28045 29003 28079 29017
rect 28045 28949 28079 28965
rect 28045 28931 28079 28949
rect 28045 28881 28079 28893
rect 28045 28859 28079 28881
rect 28045 28813 28079 28821
rect 28045 28787 28079 28813
rect 28045 28745 28079 28749
rect 28045 28715 28079 28745
rect 28045 28643 28079 28677
rect 28503 29867 28537 29901
rect 28503 29799 28537 29829
rect 28503 29795 28537 29799
rect 28503 29731 28537 29757
rect 28503 29723 28537 29731
rect 28503 29663 28537 29685
rect 28503 29651 28537 29663
rect 28503 29595 28537 29613
rect 28503 29579 28537 29595
rect 28503 29527 28537 29541
rect 28503 29507 28537 29527
rect 28503 29459 28537 29469
rect 28503 29435 28537 29459
rect 28503 29391 28537 29397
rect 28503 29363 28537 29391
rect 28503 29323 28537 29325
rect 28503 29291 28537 29323
rect 28503 29221 28537 29253
rect 28503 29219 28537 29221
rect 28503 29153 28537 29181
rect 28503 29147 28537 29153
rect 28503 29085 28537 29109
rect 28503 29075 28537 29085
rect 28503 29017 28537 29037
rect 28503 29003 28537 29017
rect 28503 28949 28537 28965
rect 28503 28931 28537 28949
rect 28503 28881 28537 28893
rect 28503 28859 28537 28881
rect 28503 28813 28537 28821
rect 28503 28787 28537 28813
rect 28503 28745 28537 28749
rect 28503 28715 28537 28745
rect 28503 28643 28537 28677
rect 28961 29867 28995 29901
rect 28961 29799 28995 29829
rect 28961 29795 28995 29799
rect 28961 29731 28995 29757
rect 28961 29723 28995 29731
rect 28961 29663 28995 29685
rect 28961 29651 28995 29663
rect 28961 29595 28995 29613
rect 28961 29579 28995 29595
rect 28961 29527 28995 29541
rect 28961 29507 28995 29527
rect 28961 29459 28995 29469
rect 28961 29435 28995 29459
rect 28961 29391 28995 29397
rect 28961 29363 28995 29391
rect 28961 29323 28995 29325
rect 28961 29291 28995 29323
rect 28961 29221 28995 29253
rect 28961 29219 28995 29221
rect 28961 29153 28995 29181
rect 28961 29147 28995 29153
rect 28961 29085 28995 29109
rect 28961 29075 28995 29085
rect 28961 29017 28995 29037
rect 28961 29003 28995 29017
rect 28961 28949 28995 28965
rect 28961 28931 28995 28949
rect 28961 28881 28995 28893
rect 28961 28859 28995 28881
rect 28961 28813 28995 28821
rect 28961 28787 28995 28813
rect 28961 28745 28995 28749
rect 28961 28715 28995 28745
rect 28961 28643 28995 28677
rect 29419 29867 29453 29901
rect 29419 29799 29453 29829
rect 29419 29795 29453 29799
rect 29419 29731 29453 29757
rect 29419 29723 29453 29731
rect 29419 29663 29453 29685
rect 29419 29651 29453 29663
rect 29419 29595 29453 29613
rect 29419 29579 29453 29595
rect 29419 29527 29453 29541
rect 29419 29507 29453 29527
rect 29419 29459 29453 29469
rect 29419 29435 29453 29459
rect 29419 29391 29453 29397
rect 29419 29363 29453 29391
rect 29419 29323 29453 29325
rect 29419 29291 29453 29323
rect 29419 29221 29453 29253
rect 29419 29219 29453 29221
rect 29419 29153 29453 29181
rect 29419 29147 29453 29153
rect 29419 29085 29453 29109
rect 29419 29075 29453 29085
rect 29419 29017 29453 29037
rect 29419 29003 29453 29017
rect 29419 28949 29453 28965
rect 29419 28931 29453 28949
rect 29419 28881 29453 28893
rect 29419 28859 29453 28881
rect 29419 28813 29453 28821
rect 29419 28787 29453 28813
rect 29419 28745 29453 28749
rect 29419 28715 29453 28745
rect 29419 28643 29453 28677
rect 29877 29867 29911 29901
rect 29877 29799 29911 29829
rect 29877 29795 29911 29799
rect 29877 29731 29911 29757
rect 29877 29723 29911 29731
rect 29877 29663 29911 29685
rect 29877 29651 29911 29663
rect 29877 29595 29911 29613
rect 29877 29579 29911 29595
rect 29877 29527 29911 29541
rect 29877 29507 29911 29527
rect 29877 29459 29911 29469
rect 29877 29435 29911 29459
rect 29877 29391 29911 29397
rect 29877 29363 29911 29391
rect 29877 29323 29911 29325
rect 29877 29291 29911 29323
rect 29877 29221 29911 29253
rect 29877 29219 29911 29221
rect 29877 29153 29911 29181
rect 29877 29147 29911 29153
rect 29877 29085 29911 29109
rect 29877 29075 29911 29085
rect 29877 29017 29911 29037
rect 29877 29003 29911 29017
rect 29877 28949 29911 28965
rect 29877 28931 29911 28949
rect 29877 28881 29911 28893
rect 29877 28859 29911 28881
rect 29877 28813 29911 28821
rect 29877 28787 29911 28813
rect 29877 28745 29911 28749
rect 29877 28715 29911 28745
rect 29877 28643 29911 28677
rect 30335 29867 30369 29901
rect 30335 29799 30369 29829
rect 30335 29795 30369 29799
rect 30335 29731 30369 29757
rect 30335 29723 30369 29731
rect 30335 29663 30369 29685
rect 30335 29651 30369 29663
rect 30335 29595 30369 29613
rect 30335 29579 30369 29595
rect 30335 29527 30369 29541
rect 30335 29507 30369 29527
rect 30335 29459 30369 29469
rect 30335 29435 30369 29459
rect 30335 29391 30369 29397
rect 30335 29363 30369 29391
rect 30335 29323 30369 29325
rect 30335 29291 30369 29323
rect 30335 29221 30369 29253
rect 30335 29219 30369 29221
rect 30335 29153 30369 29181
rect 30335 29147 30369 29153
rect 30335 29085 30369 29109
rect 30335 29075 30369 29085
rect 30335 29017 30369 29037
rect 30335 29003 30369 29017
rect 30335 28949 30369 28965
rect 30335 28931 30369 28949
rect 30335 28881 30369 28893
rect 30335 28859 30369 28881
rect 30335 28813 30369 28821
rect 30335 28787 30369 28813
rect 30335 28745 30369 28749
rect 30335 28715 30369 28745
rect 30335 28643 30369 28677
rect 30793 29867 30827 29901
rect 30793 29799 30827 29829
rect 30793 29795 30827 29799
rect 30793 29731 30827 29757
rect 30793 29723 30827 29731
rect 30793 29663 30827 29685
rect 30793 29651 30827 29663
rect 30793 29595 30827 29613
rect 30793 29579 30827 29595
rect 30793 29527 30827 29541
rect 30793 29507 30827 29527
rect 30793 29459 30827 29469
rect 30793 29435 30827 29459
rect 30793 29391 30827 29397
rect 30793 29363 30827 29391
rect 30793 29323 30827 29325
rect 30793 29291 30827 29323
rect 30793 29221 30827 29253
rect 30793 29219 30827 29221
rect 30793 29153 30827 29181
rect 30793 29147 30827 29153
rect 30793 29085 30827 29109
rect 30793 29075 30827 29085
rect 30793 29017 30827 29037
rect 30793 29003 30827 29017
rect 30793 28949 30827 28965
rect 30793 28931 30827 28949
rect 30793 28881 30827 28893
rect 30793 28859 30827 28881
rect 30793 28813 30827 28821
rect 30793 28787 30827 28813
rect 30793 28745 30827 28749
rect 30793 28715 30827 28745
rect 30793 28643 30827 28677
rect 31251 29867 31285 29901
rect 31251 29799 31285 29829
rect 31251 29795 31285 29799
rect 31251 29731 31285 29757
rect 31251 29723 31285 29731
rect 31251 29663 31285 29685
rect 31251 29651 31285 29663
rect 31251 29595 31285 29613
rect 31251 29579 31285 29595
rect 31251 29527 31285 29541
rect 31251 29507 31285 29527
rect 31251 29459 31285 29469
rect 31251 29435 31285 29459
rect 31251 29391 31285 29397
rect 31251 29363 31285 29391
rect 31251 29323 31285 29325
rect 31251 29291 31285 29323
rect 31251 29221 31285 29253
rect 31251 29219 31285 29221
rect 31251 29153 31285 29181
rect 31251 29147 31285 29153
rect 31251 29085 31285 29109
rect 31251 29075 31285 29085
rect 31251 29017 31285 29037
rect 31251 29003 31285 29017
rect 31251 28949 31285 28965
rect 31251 28931 31285 28949
rect 31251 28881 31285 28893
rect 31251 28859 31285 28881
rect 31251 28813 31285 28821
rect 31251 28787 31285 28813
rect 31251 28745 31285 28749
rect 31251 28715 31285 28745
rect 31251 28643 31285 28677
rect 31709 29867 31743 29901
rect 31709 29799 31743 29829
rect 31709 29795 31743 29799
rect 31709 29731 31743 29757
rect 31709 29723 31743 29731
rect 31709 29663 31743 29685
rect 31709 29651 31743 29663
rect 31709 29595 31743 29613
rect 31709 29579 31743 29595
rect 31709 29527 31743 29541
rect 31709 29507 31743 29527
rect 31709 29459 31743 29469
rect 31709 29435 31743 29459
rect 31709 29391 31743 29397
rect 31709 29363 31743 29391
rect 31709 29323 31743 29325
rect 31709 29291 31743 29323
rect 31709 29221 31743 29253
rect 31709 29219 31743 29221
rect 31709 29153 31743 29181
rect 31709 29147 31743 29153
rect 31709 29085 31743 29109
rect 31709 29075 31743 29085
rect 31709 29017 31743 29037
rect 31709 29003 31743 29017
rect 31709 28949 31743 28965
rect 31709 28931 31743 28949
rect 31709 28881 31743 28893
rect 31709 28859 31743 28881
rect 31709 28813 31743 28821
rect 31709 28787 31743 28813
rect 31709 28745 31743 28749
rect 31709 28715 31743 28745
rect 31709 28643 31743 28677
rect 32167 29867 32201 29901
rect 32167 29799 32201 29829
rect 32167 29795 32201 29799
rect 32167 29731 32201 29757
rect 32167 29723 32201 29731
rect 32167 29663 32201 29685
rect 32167 29651 32201 29663
rect 32167 29595 32201 29613
rect 32167 29579 32201 29595
rect 32167 29527 32201 29541
rect 32167 29507 32201 29527
rect 32167 29459 32201 29469
rect 32167 29435 32201 29459
rect 32167 29391 32201 29397
rect 32167 29363 32201 29391
rect 32167 29323 32201 29325
rect 32167 29291 32201 29323
rect 32167 29221 32201 29253
rect 32167 29219 32201 29221
rect 32167 29153 32201 29181
rect 32167 29147 32201 29153
rect 32167 29085 32201 29109
rect 32167 29075 32201 29085
rect 32167 29017 32201 29037
rect 32167 29003 32201 29017
rect 32167 28949 32201 28965
rect 32167 28931 32201 28949
rect 32167 28881 32201 28893
rect 32167 28859 32201 28881
rect 32167 28813 32201 28821
rect 32167 28787 32201 28813
rect 32167 28745 32201 28749
rect 32167 28715 32201 28745
rect 32167 28643 32201 28677
rect 32625 29867 32659 29901
rect 32625 29799 32659 29829
rect 32625 29795 32659 29799
rect 32625 29731 32659 29757
rect 32625 29723 32659 29731
rect 32625 29663 32659 29685
rect 32625 29651 32659 29663
rect 32625 29595 32659 29613
rect 32625 29579 32659 29595
rect 32625 29527 32659 29541
rect 32625 29507 32659 29527
rect 32625 29459 32659 29469
rect 32625 29435 32659 29459
rect 32625 29391 32659 29397
rect 32625 29363 32659 29391
rect 32625 29323 32659 29325
rect 32625 29291 32659 29323
rect 32625 29221 32659 29253
rect 32625 29219 32659 29221
rect 32625 29153 32659 29181
rect 32625 29147 32659 29153
rect 32625 29085 32659 29109
rect 32625 29075 32659 29085
rect 32625 29017 32659 29037
rect 32625 29003 32659 29017
rect 32625 28949 32659 28965
rect 32625 28931 32659 28949
rect 32625 28881 32659 28893
rect 32625 28859 32659 28881
rect 32625 28813 32659 28821
rect 32625 28787 32659 28813
rect 32625 28745 32659 28749
rect 32625 28715 32659 28745
rect 32625 28643 32659 28677
rect 33083 29867 33117 29901
rect 33083 29799 33117 29829
rect 33083 29795 33117 29799
rect 33083 29731 33117 29757
rect 33083 29723 33117 29731
rect 33083 29663 33117 29685
rect 33083 29651 33117 29663
rect 33083 29595 33117 29613
rect 33083 29579 33117 29595
rect 33083 29527 33117 29541
rect 33083 29507 33117 29527
rect 33083 29459 33117 29469
rect 33083 29435 33117 29459
rect 33083 29391 33117 29397
rect 33083 29363 33117 29391
rect 33083 29323 33117 29325
rect 33083 29291 33117 29323
rect 33083 29221 33117 29253
rect 33083 29219 33117 29221
rect 33083 29153 33117 29181
rect 33083 29147 33117 29153
rect 33083 29085 33117 29109
rect 33083 29075 33117 29085
rect 33083 29017 33117 29037
rect 33083 29003 33117 29017
rect 33083 28949 33117 28965
rect 33083 28931 33117 28949
rect 33083 28881 33117 28893
rect 33083 28859 33117 28881
rect 33083 28813 33117 28821
rect 33083 28787 33117 28813
rect 33083 28745 33117 28749
rect 33083 28715 33117 28745
rect 33083 28643 33117 28677
rect 33541 29867 33575 29901
rect 33541 29799 33575 29829
rect 33541 29795 33575 29799
rect 33541 29731 33575 29757
rect 33541 29723 33575 29731
rect 33541 29663 33575 29685
rect 33541 29651 33575 29663
rect 33541 29595 33575 29613
rect 33541 29579 33575 29595
rect 33541 29527 33575 29541
rect 33541 29507 33575 29527
rect 33541 29459 33575 29469
rect 33541 29435 33575 29459
rect 33541 29391 33575 29397
rect 33541 29363 33575 29391
rect 33541 29323 33575 29325
rect 33541 29291 33575 29323
rect 33541 29221 33575 29253
rect 33541 29219 33575 29221
rect 33541 29153 33575 29181
rect 33541 29147 33575 29153
rect 33541 29085 33575 29109
rect 33541 29075 33575 29085
rect 33541 29017 33575 29037
rect 33541 29003 33575 29017
rect 33541 28949 33575 28965
rect 33541 28931 33575 28949
rect 33541 28881 33575 28893
rect 33541 28859 33575 28881
rect 33541 28813 33575 28821
rect 33541 28787 33575 28813
rect 33541 28745 33575 28749
rect 33541 28715 33575 28745
rect 33541 28643 33575 28677
rect 34089 29867 34123 29901
rect 34089 29799 34123 29829
rect 34089 29795 34123 29799
rect 34089 29731 34123 29757
rect 34089 29723 34123 29731
rect 34089 29663 34123 29685
rect 34089 29651 34123 29663
rect 34089 29595 34123 29613
rect 34089 29579 34123 29595
rect 34089 29527 34123 29541
rect 34089 29507 34123 29527
rect 34089 29459 34123 29469
rect 34089 29435 34123 29459
rect 34089 29391 34123 29397
rect 34089 29363 34123 29391
rect 34089 29323 34123 29325
rect 34089 29291 34123 29323
rect 34089 29221 34123 29253
rect 34089 29219 34123 29221
rect 34089 29153 34123 29181
rect 34089 29147 34123 29153
rect 34089 29085 34123 29109
rect 34089 29075 34123 29085
rect 34089 29017 34123 29037
rect 34089 29003 34123 29017
rect 34089 28949 34123 28965
rect 34089 28931 34123 28949
rect 34089 28881 34123 28893
rect 34089 28859 34123 28881
rect 34089 28813 34123 28821
rect 34089 28787 34123 28813
rect 34089 28745 34123 28749
rect 34089 28715 34123 28745
rect 34089 28643 34123 28677
rect 34547 29867 34581 29901
rect 34547 29799 34581 29829
rect 34547 29795 34581 29799
rect 34547 29731 34581 29757
rect 34547 29723 34581 29731
rect 34547 29663 34581 29685
rect 34547 29651 34581 29663
rect 34547 29595 34581 29613
rect 34547 29579 34581 29595
rect 34547 29527 34581 29541
rect 34547 29507 34581 29527
rect 34547 29459 34581 29469
rect 34547 29435 34581 29459
rect 34547 29391 34581 29397
rect 34547 29363 34581 29391
rect 34547 29323 34581 29325
rect 34547 29291 34581 29323
rect 34547 29221 34581 29253
rect 34547 29219 34581 29221
rect 34547 29153 34581 29181
rect 34547 29147 34581 29153
rect 34547 29085 34581 29109
rect 34547 29075 34581 29085
rect 34547 29017 34581 29037
rect 34547 29003 34581 29017
rect 34547 28949 34581 28965
rect 34547 28931 34581 28949
rect 34547 28881 34581 28893
rect 34547 28859 34581 28881
rect 34547 28813 34581 28821
rect 34547 28787 34581 28813
rect 34547 28745 34581 28749
rect 34547 28715 34581 28745
rect 34547 28643 34581 28677
rect 35005 29867 35039 29901
rect 35005 29799 35039 29829
rect 35005 29795 35039 29799
rect 35005 29731 35039 29757
rect 35005 29723 35039 29731
rect 35005 29663 35039 29685
rect 35005 29651 35039 29663
rect 35005 29595 35039 29613
rect 35005 29579 35039 29595
rect 35005 29527 35039 29541
rect 35005 29507 35039 29527
rect 35005 29459 35039 29469
rect 35005 29435 35039 29459
rect 35005 29391 35039 29397
rect 35005 29363 35039 29391
rect 35005 29323 35039 29325
rect 35005 29291 35039 29323
rect 35005 29221 35039 29253
rect 35005 29219 35039 29221
rect 35005 29153 35039 29181
rect 35005 29147 35039 29153
rect 35005 29085 35039 29109
rect 35005 29075 35039 29085
rect 35005 29017 35039 29037
rect 35005 29003 35039 29017
rect 35005 28949 35039 28965
rect 35005 28931 35039 28949
rect 35005 28881 35039 28893
rect 35005 28859 35039 28881
rect 35005 28813 35039 28821
rect 35005 28787 35039 28813
rect 35005 28745 35039 28749
rect 35005 28715 35039 28745
rect 35005 28643 35039 28677
rect 35463 29867 35497 29901
rect 35463 29799 35497 29829
rect 35463 29795 35497 29799
rect 35463 29731 35497 29757
rect 35463 29723 35497 29731
rect 35463 29663 35497 29685
rect 35463 29651 35497 29663
rect 35463 29595 35497 29613
rect 35463 29579 35497 29595
rect 35463 29527 35497 29541
rect 35463 29507 35497 29527
rect 35463 29459 35497 29469
rect 35463 29435 35497 29459
rect 35463 29391 35497 29397
rect 35463 29363 35497 29391
rect 35463 29323 35497 29325
rect 35463 29291 35497 29323
rect 35463 29221 35497 29253
rect 35463 29219 35497 29221
rect 35463 29153 35497 29181
rect 35463 29147 35497 29153
rect 35463 29085 35497 29109
rect 35463 29075 35497 29085
rect 35463 29017 35497 29037
rect 35463 29003 35497 29017
rect 35463 28949 35497 28965
rect 35463 28931 35497 28949
rect 35463 28881 35497 28893
rect 35463 28859 35497 28881
rect 35463 28813 35497 28821
rect 35463 28787 35497 28813
rect 35463 28745 35497 28749
rect 35463 28715 35497 28745
rect 35463 28643 35497 28677
rect 35921 29867 35955 29901
rect 35921 29799 35955 29829
rect 35921 29795 35955 29799
rect 35921 29731 35955 29757
rect 35921 29723 35955 29731
rect 35921 29663 35955 29685
rect 35921 29651 35955 29663
rect 35921 29595 35955 29613
rect 35921 29579 35955 29595
rect 35921 29527 35955 29541
rect 35921 29507 35955 29527
rect 35921 29459 35955 29469
rect 35921 29435 35955 29459
rect 35921 29391 35955 29397
rect 35921 29363 35955 29391
rect 35921 29323 35955 29325
rect 35921 29291 35955 29323
rect 35921 29221 35955 29253
rect 35921 29219 35955 29221
rect 35921 29153 35955 29181
rect 35921 29147 35955 29153
rect 35921 29085 35955 29109
rect 35921 29075 35955 29085
rect 35921 29017 35955 29037
rect 35921 29003 35955 29017
rect 35921 28949 35955 28965
rect 35921 28931 35955 28949
rect 35921 28881 35955 28893
rect 35921 28859 35955 28881
rect 35921 28813 35955 28821
rect 35921 28787 35955 28813
rect 35921 28745 35955 28749
rect 35921 28715 35955 28745
rect 35921 28643 35955 28677
rect 36379 29867 36413 29901
rect 36379 29799 36413 29829
rect 36379 29795 36413 29799
rect 36379 29731 36413 29757
rect 36379 29723 36413 29731
rect 36379 29663 36413 29685
rect 36379 29651 36413 29663
rect 36379 29595 36413 29613
rect 36379 29579 36413 29595
rect 36379 29527 36413 29541
rect 36379 29507 36413 29527
rect 36379 29459 36413 29469
rect 36379 29435 36413 29459
rect 36379 29391 36413 29397
rect 36379 29363 36413 29391
rect 36379 29323 36413 29325
rect 36379 29291 36413 29323
rect 36379 29221 36413 29253
rect 36379 29219 36413 29221
rect 36379 29153 36413 29181
rect 36379 29147 36413 29153
rect 36379 29085 36413 29109
rect 36379 29075 36413 29085
rect 36379 29017 36413 29037
rect 36379 29003 36413 29017
rect 36379 28949 36413 28965
rect 36379 28931 36413 28949
rect 36379 28881 36413 28893
rect 36379 28859 36413 28881
rect 36379 28813 36413 28821
rect 36379 28787 36413 28813
rect 36379 28745 36413 28749
rect 36379 28715 36413 28745
rect 36379 28643 36413 28677
rect 36837 29867 36871 29901
rect 36837 29799 36871 29829
rect 36837 29795 36871 29799
rect 36837 29731 36871 29757
rect 36837 29723 36871 29731
rect 36837 29663 36871 29685
rect 36837 29651 36871 29663
rect 36837 29595 36871 29613
rect 36837 29579 36871 29595
rect 36837 29527 36871 29541
rect 36837 29507 36871 29527
rect 36837 29459 36871 29469
rect 36837 29435 36871 29459
rect 36837 29391 36871 29397
rect 36837 29363 36871 29391
rect 37413 29363 37807 29901
rect 39420 29363 39814 29901
rect 40157 29363 40551 29901
rect 42164 29363 42558 29901
rect 36837 29323 36871 29325
rect 36837 29291 36871 29323
rect 36837 29221 36871 29253
rect 36837 29219 36871 29221
rect 36837 29153 36871 29181
rect 36837 29147 36871 29153
rect 36837 29085 36871 29109
rect 36837 29075 36871 29085
rect 36837 29017 36871 29037
rect 36837 29003 36871 29017
rect 36837 28949 36871 28965
rect 36837 28931 36871 28949
rect 36837 28881 36871 28893
rect 36837 28859 36871 28881
rect 36837 28813 36871 28821
rect 36837 28787 36871 28813
rect 36837 28745 36871 28749
rect 36837 28715 36871 28745
rect 36837 28643 36871 28677
rect 12541 28373 12575 28407
rect 14197 28389 14231 28407
rect 23397 28389 23431 28407
rect 14197 28373 14231 28389
rect 23397 28373 23431 28389
rect 34069 28373 34103 28407
rect 37413 28403 37807 28941
rect 39420 28403 39814 28941
rect 40157 28403 40551 28941
rect 42164 28403 42558 28941
rect 6197 28255 6231 28289
rect 6597 28255 6631 28289
rect 6997 28255 7031 28289
rect 7397 28255 7431 28289
rect 7797 28255 7831 28289
rect 8197 28255 8231 28289
rect 8597 28255 8631 28289
rect 8997 28255 9031 28289
rect 9397 28255 9431 28289
rect 9797 28255 9831 28289
rect 10197 28255 10231 28289
rect 10597 28255 10631 28289
rect 10997 28255 11031 28289
rect 11397 28255 11431 28289
rect 11797 28255 11831 28289
rect 12197 28255 12231 28289
rect 12597 28255 12631 28289
rect 12997 28255 13031 28289
rect 13397 28255 13431 28289
rect 13797 28255 13831 28289
rect 14197 28255 14231 28289
rect 14597 28255 14631 28289
rect 14997 28255 15031 28289
rect 15397 28255 15431 28289
rect 15797 28255 15831 28289
rect 16197 28255 16231 28289
rect 16597 28255 16631 28289
rect 16997 28255 17031 28289
rect 17397 28255 17431 28289
rect 17797 28255 17831 28289
rect 18197 28255 18231 28289
rect 18597 28255 18631 28289
rect 18997 28255 19031 28289
rect 19397 28255 19431 28289
rect 19797 28255 19831 28289
rect 20197 28255 20231 28289
rect 20597 28255 20631 28289
rect 20997 28255 21031 28289
rect 21397 28255 21431 28289
rect 21797 28255 21831 28289
rect 22197 28255 22231 28289
rect 22597 28255 22631 28289
rect 22997 28255 23031 28289
rect 23397 28255 23431 28289
rect 23797 28255 23831 28289
rect 24197 28255 24231 28289
rect 24597 28255 24631 28289
rect 24997 28255 25031 28289
rect 25397 28255 25431 28289
rect 25797 28255 25831 28289
rect 26197 28255 26231 28289
rect 26597 28255 26631 28289
rect 26997 28255 27031 28289
rect 27397 28255 27431 28289
rect 27797 28255 27831 28289
rect 28197 28255 28231 28289
rect 28597 28255 28631 28289
rect 28997 28255 29031 28289
rect 29397 28255 29431 28289
rect 29797 28255 29831 28289
rect 30197 28255 30231 28289
rect 30597 28255 30631 28289
rect 30997 28255 31031 28289
rect 31397 28255 31431 28289
rect 31797 28255 31831 28289
rect 32197 28255 32231 28289
rect 32597 28255 32631 28289
rect 32997 28255 33031 28289
rect 33397 28255 33431 28289
rect 34225 28255 34259 28289
rect 34625 28255 34659 28289
rect 35025 28255 35059 28289
rect 35425 28255 35459 28289
rect 35825 28255 35859 28289
rect 36225 28255 36259 28289
rect 36625 28255 36659 28289
rect 37577 28255 37611 28289
rect 37777 28255 37811 28289
rect 37977 28255 38011 28289
rect 38177 28255 38211 28289
rect 38377 28255 38411 28289
rect 38577 28255 38611 28289
rect 38777 28255 38811 28289
rect 38977 28255 39011 28289
rect 39177 28255 39211 28289
rect 39377 28255 39411 28289
rect 39577 28255 39611 28289
rect 40321 28255 40355 28289
rect 40521 28255 40555 28289
rect 40721 28255 40755 28289
rect 40921 28255 40955 28289
rect 41121 28255 41155 28289
rect 41321 28255 41355 28289
rect 41521 28255 41555 28289
rect 41721 28255 41755 28289
rect 41921 28255 41955 28289
rect 42121 28255 42155 28289
rect 42321 28255 42355 28289
rect 6903 26375 6937 26409
rect 7103 26375 7137 26409
rect 7303 26375 7337 26409
rect 7503 26375 7537 26409
rect 7703 26375 7737 26409
rect 7903 26375 7937 26409
rect 8103 26375 8137 26409
rect 8303 26375 8337 26409
rect 8503 26375 8537 26409
rect 8703 26375 8737 26409
rect 8903 26375 8937 26409
rect 9725 26375 9759 26409
rect 10125 26375 10159 26409
rect 10525 26375 10559 26409
rect 10925 26375 10959 26409
rect 11325 26375 11359 26409
rect 11725 26375 11759 26409
rect 12125 26375 12159 26409
rect 12525 26375 12559 26409
rect 12925 26375 12959 26409
rect 13325 26375 13359 26409
rect 13725 26375 13759 26409
rect 14125 26375 14159 26409
rect 14525 26375 14559 26409
rect 14925 26375 14959 26409
rect 15607 26375 15641 26409
rect 16007 26375 16041 26409
rect 16407 26375 16441 26409
rect 16807 26375 16841 26409
rect 17207 26375 17241 26409
rect 17607 26375 17641 26409
rect 18007 26375 18041 26409
rect 18407 26375 18441 26409
rect 18807 26375 18841 26409
rect 19207 26375 19241 26409
rect 19607 26375 19641 26409
rect 20007 26375 20041 26409
rect 20407 26375 20441 26409
rect 20807 26375 20841 26409
rect 21207 26375 21241 26409
rect 21607 26375 21641 26409
rect 22007 26375 22041 26409
rect 22407 26375 22441 26409
rect 23151 26375 23185 26409
rect 23551 26375 23585 26409
rect 23951 26375 23985 26409
rect 24351 26375 24385 26409
rect 24751 26375 24785 26409
rect 25151 26375 25185 26409
rect 25551 26375 25585 26409
rect 25951 26375 25985 26409
rect 26351 26375 26385 26409
rect 26751 26375 26785 26409
rect 28443 26375 28477 26409
rect 28643 26375 28677 26409
rect 28843 26375 28877 26409
rect 29043 26375 29077 26409
rect 29243 26375 29277 26409
rect 29443 26375 29477 26409
rect 29643 26375 29677 26409
rect 29843 26375 29877 26409
rect 30043 26375 30077 26409
rect 30243 26375 30277 26409
rect 30443 26375 30477 26409
rect 30643 26375 30677 26409
rect 30843 26375 30877 26409
rect 31043 26375 31077 26409
rect 31243 26375 31277 26409
rect 31443 26375 31477 26409
rect 31643 26375 31677 26409
rect 31843 26375 31877 26409
rect 32043 26375 32077 26409
rect 32243 26375 32277 26409
rect 32443 26375 32477 26409
rect 32643 26375 32677 26409
rect 32843 26375 32877 26409
rect 33043 26375 33077 26409
rect 33243 26375 33277 26409
rect 33443 26375 33477 26409
rect 33643 26375 33677 26409
rect 33843 26375 33877 26409
rect 34043 26375 34077 26409
rect 34243 26375 34277 26409
rect 34443 26375 34477 26409
rect 34643 26375 34677 26409
rect 34843 26375 34877 26409
rect 35043 26375 35077 26409
rect 35243 26375 35277 26409
rect 35443 26375 35477 26409
rect 35643 26375 35677 26409
rect 35843 26375 35877 26409
rect 36043 26375 36077 26409
rect 36243 26375 36277 26409
rect 36443 26375 36477 26409
rect 36643 26375 36677 26409
rect 36843 26375 36877 26409
rect 37043 26375 37077 26409
rect 37243 26375 37277 26409
rect 37443 26375 37477 26409
rect 37643 26375 37677 26409
rect 37843 26375 37877 26409
rect 38043 26375 38077 26409
rect 38243 26375 38277 26409
rect 38443 26375 38477 26409
rect 38643 26375 38677 26409
rect 38843 26375 38877 26409
rect 39929 26375 39963 26409
rect 40129 26375 40163 26409
rect 40329 26375 40363 26409
rect 40529 26375 40563 26409
rect 40729 26375 40763 26409
rect 40929 26375 40963 26409
rect 41129 26375 41163 26409
rect 41329 26375 41363 26409
rect 41529 26375 41563 26409
rect 41729 26375 41763 26409
rect 41929 26375 41963 26409
rect 6739 25603 7133 26141
rect 8746 25603 9140 26141
rect 6739 24643 7133 25181
rect 8746 24643 9140 25181
rect 9589 26107 9623 26141
rect 9589 26039 9623 26069
rect 9589 26035 9623 26039
rect 9589 25971 9623 25997
rect 9589 25963 9623 25971
rect 9589 25903 9623 25925
rect 9589 25891 9623 25903
rect 9589 25835 9623 25853
rect 9589 25819 9623 25835
rect 9589 25767 9623 25781
rect 9589 25747 9623 25767
rect 9589 25699 9623 25709
rect 9589 25675 9623 25699
rect 9589 25631 9623 25637
rect 9589 25603 9623 25631
rect 9589 25563 9623 25565
rect 9589 25531 9623 25563
rect 9589 25461 9623 25493
rect 9589 25459 9623 25461
rect 9589 25393 9623 25421
rect 9589 25387 9623 25393
rect 9589 25325 9623 25349
rect 9589 25315 9623 25325
rect 9589 25257 9623 25277
rect 9589 25243 9623 25257
rect 9589 25189 9623 25205
rect 9589 25171 9623 25189
rect 9589 25121 9623 25133
rect 9589 25099 9623 25121
rect 9589 25053 9623 25061
rect 9589 25027 9623 25053
rect 9589 24985 9623 24989
rect 9589 24955 9623 24985
rect 9589 24883 9623 24917
rect 10047 26107 10081 26141
rect 10047 26039 10081 26069
rect 10047 26035 10081 26039
rect 10047 25971 10081 25997
rect 10047 25963 10081 25971
rect 10047 25903 10081 25925
rect 10047 25891 10081 25903
rect 10047 25835 10081 25853
rect 10047 25819 10081 25835
rect 10047 25767 10081 25781
rect 10047 25747 10081 25767
rect 10047 25699 10081 25709
rect 10047 25675 10081 25699
rect 10047 25631 10081 25637
rect 10047 25603 10081 25631
rect 10047 25563 10081 25565
rect 10047 25531 10081 25563
rect 10047 25461 10081 25493
rect 10047 25459 10081 25461
rect 10047 25393 10081 25421
rect 10047 25387 10081 25393
rect 10047 25325 10081 25349
rect 10047 25315 10081 25325
rect 10047 25257 10081 25277
rect 10047 25243 10081 25257
rect 10047 25189 10081 25205
rect 10047 25171 10081 25189
rect 10047 25121 10081 25133
rect 10047 25099 10081 25121
rect 10047 25053 10081 25061
rect 10047 25027 10081 25053
rect 10047 24985 10081 24989
rect 10047 24955 10081 24985
rect 10047 24883 10081 24917
rect 10505 26107 10539 26141
rect 10505 26039 10539 26069
rect 10505 26035 10539 26039
rect 10505 25971 10539 25997
rect 10505 25963 10539 25971
rect 10505 25903 10539 25925
rect 10505 25891 10539 25903
rect 10505 25835 10539 25853
rect 10505 25819 10539 25835
rect 10505 25767 10539 25781
rect 10505 25747 10539 25767
rect 10505 25699 10539 25709
rect 10505 25675 10539 25699
rect 10505 25631 10539 25637
rect 10505 25603 10539 25631
rect 10505 25563 10539 25565
rect 10505 25531 10539 25563
rect 10505 25461 10539 25493
rect 10505 25459 10539 25461
rect 10505 25393 10539 25421
rect 10505 25387 10539 25393
rect 10505 25325 10539 25349
rect 10505 25315 10539 25325
rect 10505 25257 10539 25277
rect 10505 25243 10539 25257
rect 10505 25189 10539 25205
rect 10505 25171 10539 25189
rect 10505 25121 10539 25133
rect 10505 25099 10539 25121
rect 10505 25053 10539 25061
rect 10505 25027 10539 25053
rect 10505 24985 10539 24989
rect 10505 24955 10539 24985
rect 10505 24883 10539 24917
rect 10963 26107 10997 26141
rect 10963 26039 10997 26069
rect 10963 26035 10997 26039
rect 10963 25971 10997 25997
rect 10963 25963 10997 25971
rect 10963 25903 10997 25925
rect 10963 25891 10997 25903
rect 10963 25835 10997 25853
rect 10963 25819 10997 25835
rect 10963 25767 10997 25781
rect 10963 25747 10997 25767
rect 10963 25699 10997 25709
rect 10963 25675 10997 25699
rect 10963 25631 10997 25637
rect 10963 25603 10997 25631
rect 10963 25563 10997 25565
rect 10963 25531 10997 25563
rect 10963 25461 10997 25493
rect 10963 25459 10997 25461
rect 10963 25393 10997 25421
rect 10963 25387 10997 25393
rect 10963 25325 10997 25349
rect 10963 25315 10997 25325
rect 10963 25257 10997 25277
rect 10963 25243 10997 25257
rect 10963 25189 10997 25205
rect 10963 25171 10997 25189
rect 10963 25121 10997 25133
rect 10963 25099 10997 25121
rect 10963 25053 10997 25061
rect 10963 25027 10997 25053
rect 10963 24985 10997 24989
rect 10963 24955 10997 24985
rect 10963 24883 10997 24917
rect 11421 26107 11455 26141
rect 11421 26039 11455 26069
rect 11421 26035 11455 26039
rect 11421 25971 11455 25997
rect 11421 25963 11455 25971
rect 11421 25903 11455 25925
rect 11421 25891 11455 25903
rect 11421 25835 11455 25853
rect 11421 25819 11455 25835
rect 11421 25767 11455 25781
rect 11421 25747 11455 25767
rect 11421 25699 11455 25709
rect 11421 25675 11455 25699
rect 11421 25631 11455 25637
rect 11421 25603 11455 25631
rect 11421 25563 11455 25565
rect 11421 25531 11455 25563
rect 11421 25461 11455 25493
rect 11421 25459 11455 25461
rect 11421 25393 11455 25421
rect 11421 25387 11455 25393
rect 11421 25325 11455 25349
rect 11421 25315 11455 25325
rect 11421 25257 11455 25277
rect 11421 25243 11455 25257
rect 11421 25189 11455 25205
rect 11421 25171 11455 25189
rect 11421 25121 11455 25133
rect 11421 25099 11455 25121
rect 11421 25053 11455 25061
rect 11421 25027 11455 25053
rect 11421 24985 11455 24989
rect 11421 24955 11455 24985
rect 11421 24883 11455 24917
rect 11879 26107 11913 26141
rect 11879 26039 11913 26069
rect 11879 26035 11913 26039
rect 11879 25971 11913 25997
rect 11879 25963 11913 25971
rect 11879 25903 11913 25925
rect 11879 25891 11913 25903
rect 11879 25835 11913 25853
rect 11879 25819 11913 25835
rect 11879 25767 11913 25781
rect 11879 25747 11913 25767
rect 11879 25699 11913 25709
rect 11879 25675 11913 25699
rect 11879 25631 11913 25637
rect 11879 25603 11913 25631
rect 11879 25563 11913 25565
rect 11879 25531 11913 25563
rect 11879 25461 11913 25493
rect 11879 25459 11913 25461
rect 11879 25393 11913 25421
rect 11879 25387 11913 25393
rect 11879 25325 11913 25349
rect 11879 25315 11913 25325
rect 11879 25257 11913 25277
rect 11879 25243 11913 25257
rect 11879 25189 11913 25205
rect 11879 25171 11913 25189
rect 11879 25121 11913 25133
rect 11879 25099 11913 25121
rect 11879 25053 11913 25061
rect 11879 25027 11913 25053
rect 11879 24985 11913 24989
rect 11879 24955 11913 24985
rect 11879 24883 11913 24917
rect 12337 26107 12371 26141
rect 12337 26039 12371 26069
rect 12337 26035 12371 26039
rect 12337 25971 12371 25997
rect 12337 25963 12371 25971
rect 12337 25903 12371 25925
rect 12337 25891 12371 25903
rect 12337 25835 12371 25853
rect 12337 25819 12371 25835
rect 12337 25767 12371 25781
rect 12337 25747 12371 25767
rect 12337 25699 12371 25709
rect 12337 25675 12371 25699
rect 12337 25631 12371 25637
rect 12337 25603 12371 25631
rect 12337 25563 12371 25565
rect 12337 25531 12371 25563
rect 12337 25461 12371 25493
rect 12337 25459 12371 25461
rect 12337 25393 12371 25421
rect 12337 25387 12371 25393
rect 12337 25325 12371 25349
rect 12337 25315 12371 25325
rect 12337 25257 12371 25277
rect 12337 25243 12371 25257
rect 12337 25189 12371 25205
rect 12337 25171 12371 25189
rect 12337 25121 12371 25133
rect 12337 25099 12371 25121
rect 12337 25053 12371 25061
rect 12337 25027 12371 25053
rect 12337 24985 12371 24989
rect 12337 24955 12371 24985
rect 12337 24883 12371 24917
rect 12795 26107 12829 26141
rect 12795 26039 12829 26069
rect 12795 26035 12829 26039
rect 12795 25971 12829 25997
rect 12795 25963 12829 25971
rect 12795 25903 12829 25925
rect 12795 25891 12829 25903
rect 12795 25835 12829 25853
rect 12795 25819 12829 25835
rect 12795 25767 12829 25781
rect 12795 25747 12829 25767
rect 12795 25699 12829 25709
rect 12795 25675 12829 25699
rect 12795 25631 12829 25637
rect 12795 25603 12829 25631
rect 12795 25563 12829 25565
rect 12795 25531 12829 25563
rect 12795 25461 12829 25493
rect 12795 25459 12829 25461
rect 12795 25393 12829 25421
rect 12795 25387 12829 25393
rect 12795 25325 12829 25349
rect 12795 25315 12829 25325
rect 12795 25257 12829 25277
rect 12795 25243 12829 25257
rect 12795 25189 12829 25205
rect 12795 25171 12829 25189
rect 12795 25121 12829 25133
rect 12795 25099 12829 25121
rect 12795 25053 12829 25061
rect 12795 25027 12829 25053
rect 12795 24985 12829 24989
rect 12795 24955 12829 24985
rect 12795 24883 12829 24917
rect 13253 26107 13287 26141
rect 13253 26039 13287 26069
rect 13253 26035 13287 26039
rect 13253 25971 13287 25997
rect 13253 25963 13287 25971
rect 13253 25903 13287 25925
rect 13253 25891 13287 25903
rect 13253 25835 13287 25853
rect 13253 25819 13287 25835
rect 13253 25767 13287 25781
rect 13253 25747 13287 25767
rect 13253 25699 13287 25709
rect 13253 25675 13287 25699
rect 13253 25631 13287 25637
rect 13253 25603 13287 25631
rect 13253 25563 13287 25565
rect 13253 25531 13287 25563
rect 13253 25461 13287 25493
rect 13253 25459 13287 25461
rect 13253 25393 13287 25421
rect 13253 25387 13287 25393
rect 13253 25325 13287 25349
rect 13253 25315 13287 25325
rect 13253 25257 13287 25277
rect 13253 25243 13287 25257
rect 13253 25189 13287 25205
rect 13253 25171 13287 25189
rect 13253 25121 13287 25133
rect 13253 25099 13287 25121
rect 13253 25053 13287 25061
rect 13253 25027 13287 25053
rect 13253 24985 13287 24989
rect 13253 24955 13287 24985
rect 13253 24883 13287 24917
rect 13711 26107 13745 26141
rect 13711 26039 13745 26069
rect 13711 26035 13745 26039
rect 13711 25971 13745 25997
rect 13711 25963 13745 25971
rect 13711 25903 13745 25925
rect 13711 25891 13745 25903
rect 13711 25835 13745 25853
rect 13711 25819 13745 25835
rect 13711 25767 13745 25781
rect 13711 25747 13745 25767
rect 13711 25699 13745 25709
rect 13711 25675 13745 25699
rect 13711 25631 13745 25637
rect 13711 25603 13745 25631
rect 13711 25563 13745 25565
rect 13711 25531 13745 25563
rect 13711 25461 13745 25493
rect 13711 25459 13745 25461
rect 13711 25393 13745 25421
rect 13711 25387 13745 25393
rect 13711 25325 13745 25349
rect 13711 25315 13745 25325
rect 13711 25257 13745 25277
rect 13711 25243 13745 25257
rect 13711 25189 13745 25205
rect 13711 25171 13745 25189
rect 13711 25121 13745 25133
rect 13711 25099 13745 25121
rect 13711 25053 13745 25061
rect 13711 25027 13745 25053
rect 13711 24985 13745 24989
rect 13711 24955 13745 24985
rect 13711 24883 13745 24917
rect 14169 26107 14203 26141
rect 14169 26039 14203 26069
rect 14169 26035 14203 26039
rect 14169 25971 14203 25997
rect 14169 25963 14203 25971
rect 14169 25903 14203 25925
rect 14169 25891 14203 25903
rect 14169 25835 14203 25853
rect 14169 25819 14203 25835
rect 14169 25767 14203 25781
rect 14169 25747 14203 25767
rect 14169 25699 14203 25709
rect 14169 25675 14203 25699
rect 14169 25631 14203 25637
rect 14169 25603 14203 25631
rect 14169 25563 14203 25565
rect 14169 25531 14203 25563
rect 14169 25461 14203 25493
rect 14169 25459 14203 25461
rect 14169 25393 14203 25421
rect 14169 25387 14203 25393
rect 14169 25325 14203 25349
rect 14169 25315 14203 25325
rect 14169 25257 14203 25277
rect 14169 25243 14203 25257
rect 14169 25189 14203 25205
rect 14169 25171 14203 25189
rect 14169 25121 14203 25133
rect 14169 25099 14203 25121
rect 14169 25053 14203 25061
rect 14169 25027 14203 25053
rect 14169 24985 14203 24989
rect 14169 24955 14203 24985
rect 14169 24883 14203 24917
rect 14627 26107 14661 26141
rect 14627 26039 14661 26069
rect 14627 26035 14661 26039
rect 14627 25971 14661 25997
rect 14627 25963 14661 25971
rect 14627 25903 14661 25925
rect 14627 25891 14661 25903
rect 14627 25835 14661 25853
rect 14627 25819 14661 25835
rect 14627 25767 14661 25781
rect 14627 25747 14661 25767
rect 14627 25699 14661 25709
rect 14627 25675 14661 25699
rect 14627 25631 14661 25637
rect 14627 25603 14661 25631
rect 14627 25563 14661 25565
rect 14627 25531 14661 25563
rect 14627 25461 14661 25493
rect 14627 25459 14661 25461
rect 14627 25393 14661 25421
rect 14627 25387 14661 25393
rect 14627 25325 14661 25349
rect 14627 25315 14661 25325
rect 14627 25257 14661 25277
rect 14627 25243 14661 25257
rect 14627 25189 14661 25205
rect 14627 25171 14661 25189
rect 14627 25121 14661 25133
rect 14627 25099 14661 25121
rect 14627 25053 14661 25061
rect 14627 25027 14661 25053
rect 14627 24985 14661 24989
rect 14627 24955 14661 24985
rect 14627 24883 14661 24917
rect 15085 26107 15119 26141
rect 15085 26039 15119 26069
rect 15085 26035 15119 26039
rect 15085 25971 15119 25997
rect 15085 25963 15119 25971
rect 15085 25903 15119 25925
rect 26157 26197 26191 26231
rect 28306 26042 28340 26076
rect 28396 26061 28430 26076
rect 28486 26061 28520 26076
rect 28576 26061 28610 26076
rect 28666 26061 28700 26076
rect 28756 26061 28790 26076
rect 28846 26061 28880 26076
rect 28936 26061 28970 26076
rect 29026 26061 29060 26076
rect 29116 26061 29150 26076
rect 29206 26061 29240 26076
rect 29296 26061 29330 26076
rect 29386 26061 29420 26076
rect 28396 26042 28416 26061
rect 28416 26042 28430 26061
rect 28486 26042 28506 26061
rect 28506 26042 28520 26061
rect 28576 26042 28596 26061
rect 28596 26042 28610 26061
rect 28666 26042 28686 26061
rect 28686 26042 28700 26061
rect 28756 26042 28776 26061
rect 28776 26042 28790 26061
rect 28846 26042 28866 26061
rect 28866 26042 28880 26061
rect 28936 26042 28956 26061
rect 28956 26042 28970 26061
rect 29026 26042 29046 26061
rect 29046 26042 29060 26061
rect 29116 26042 29136 26061
rect 29136 26042 29150 26061
rect 29206 26042 29226 26061
rect 29226 26042 29240 26061
rect 29296 26042 29316 26061
rect 29316 26042 29330 26061
rect 29386 26042 29406 26061
rect 29406 26042 29420 26061
rect 29476 26042 29510 26076
rect 29646 26042 29680 26076
rect 29736 26061 29770 26076
rect 29826 26061 29860 26076
rect 29916 26061 29950 26076
rect 30006 26061 30040 26076
rect 30096 26061 30130 26076
rect 30186 26061 30220 26076
rect 30276 26061 30310 26076
rect 30366 26061 30400 26076
rect 30456 26061 30490 26076
rect 30546 26061 30580 26076
rect 30636 26061 30670 26076
rect 30726 26061 30760 26076
rect 29736 26042 29756 26061
rect 29756 26042 29770 26061
rect 29826 26042 29846 26061
rect 29846 26042 29860 26061
rect 29916 26042 29936 26061
rect 29936 26042 29950 26061
rect 30006 26042 30026 26061
rect 30026 26042 30040 26061
rect 30096 26042 30116 26061
rect 30116 26042 30130 26061
rect 30186 26042 30206 26061
rect 30206 26042 30220 26061
rect 30276 26042 30296 26061
rect 30296 26042 30310 26061
rect 30366 26042 30386 26061
rect 30386 26042 30400 26061
rect 30456 26042 30476 26061
rect 30476 26042 30490 26061
rect 30546 26042 30566 26061
rect 30566 26042 30580 26061
rect 30636 26042 30656 26061
rect 30656 26042 30670 26061
rect 30726 26042 30746 26061
rect 30746 26042 30760 26061
rect 30816 26042 30850 26076
rect 30986 26042 31020 26076
rect 31076 26061 31110 26076
rect 31166 26061 31200 26076
rect 31256 26061 31290 26076
rect 31346 26061 31380 26076
rect 31436 26061 31470 26076
rect 31526 26061 31560 26076
rect 31616 26061 31650 26076
rect 31706 26061 31740 26076
rect 31796 26061 31830 26076
rect 31886 26061 31920 26076
rect 31976 26061 32010 26076
rect 32066 26061 32100 26076
rect 31076 26042 31096 26061
rect 31096 26042 31110 26061
rect 31166 26042 31186 26061
rect 31186 26042 31200 26061
rect 31256 26042 31276 26061
rect 31276 26042 31290 26061
rect 31346 26042 31366 26061
rect 31366 26042 31380 26061
rect 31436 26042 31456 26061
rect 31456 26042 31470 26061
rect 31526 26042 31546 26061
rect 31546 26042 31560 26061
rect 31616 26042 31636 26061
rect 31636 26042 31650 26061
rect 31706 26042 31726 26061
rect 31726 26042 31740 26061
rect 31796 26042 31816 26061
rect 31816 26042 31830 26061
rect 31886 26042 31906 26061
rect 31906 26042 31920 26061
rect 31976 26042 31996 26061
rect 31996 26042 32010 26061
rect 32066 26042 32086 26061
rect 32086 26042 32100 26061
rect 32156 26042 32190 26076
rect 32326 26042 32360 26076
rect 32416 26061 32450 26076
rect 32506 26061 32540 26076
rect 32596 26061 32630 26076
rect 32686 26061 32720 26076
rect 32776 26061 32810 26076
rect 32866 26061 32900 26076
rect 32956 26061 32990 26076
rect 33046 26061 33080 26076
rect 33136 26061 33170 26076
rect 33226 26061 33260 26076
rect 33316 26061 33350 26076
rect 33406 26061 33440 26076
rect 32416 26042 32436 26061
rect 32436 26042 32450 26061
rect 32506 26042 32526 26061
rect 32526 26042 32540 26061
rect 32596 26042 32616 26061
rect 32616 26042 32630 26061
rect 32686 26042 32706 26061
rect 32706 26042 32720 26061
rect 32776 26042 32796 26061
rect 32796 26042 32810 26061
rect 32866 26042 32886 26061
rect 32886 26042 32900 26061
rect 32956 26042 32976 26061
rect 32976 26042 32990 26061
rect 33046 26042 33066 26061
rect 33066 26042 33080 26061
rect 33136 26042 33156 26061
rect 33156 26042 33170 26061
rect 33226 26042 33246 26061
rect 33246 26042 33260 26061
rect 33316 26042 33336 26061
rect 33336 26042 33350 26061
rect 33406 26042 33426 26061
rect 33426 26042 33440 26061
rect 33496 26042 33530 26076
rect 33666 26042 33700 26076
rect 33756 26061 33790 26076
rect 33846 26061 33880 26076
rect 33936 26061 33970 26076
rect 34026 26061 34060 26076
rect 34116 26061 34150 26076
rect 34206 26061 34240 26076
rect 34296 26061 34330 26076
rect 34386 26061 34420 26076
rect 34476 26061 34510 26076
rect 34566 26061 34600 26076
rect 34656 26061 34690 26076
rect 34746 26061 34780 26076
rect 33756 26042 33776 26061
rect 33776 26042 33790 26061
rect 33846 26042 33866 26061
rect 33866 26042 33880 26061
rect 33936 26042 33956 26061
rect 33956 26042 33970 26061
rect 34026 26042 34046 26061
rect 34046 26042 34060 26061
rect 34116 26042 34136 26061
rect 34136 26042 34150 26061
rect 34206 26042 34226 26061
rect 34226 26042 34240 26061
rect 34296 26042 34316 26061
rect 34316 26042 34330 26061
rect 34386 26042 34406 26061
rect 34406 26042 34420 26061
rect 34476 26042 34496 26061
rect 34496 26042 34510 26061
rect 34566 26042 34586 26061
rect 34586 26042 34600 26061
rect 34656 26042 34676 26061
rect 34676 26042 34690 26061
rect 34746 26042 34766 26061
rect 34766 26042 34780 26061
rect 34836 26042 34870 26076
rect 35006 26042 35040 26076
rect 35096 26061 35130 26076
rect 35186 26061 35220 26076
rect 35276 26061 35310 26076
rect 35366 26061 35400 26076
rect 35456 26061 35490 26076
rect 35546 26061 35580 26076
rect 35636 26061 35670 26076
rect 35726 26061 35760 26076
rect 35816 26061 35850 26076
rect 35906 26061 35940 26076
rect 35996 26061 36030 26076
rect 36086 26061 36120 26076
rect 35096 26042 35116 26061
rect 35116 26042 35130 26061
rect 35186 26042 35206 26061
rect 35206 26042 35220 26061
rect 35276 26042 35296 26061
rect 35296 26042 35310 26061
rect 35366 26042 35386 26061
rect 35386 26042 35400 26061
rect 35456 26042 35476 26061
rect 35476 26042 35490 26061
rect 35546 26042 35566 26061
rect 35566 26042 35580 26061
rect 35636 26042 35656 26061
rect 35656 26042 35670 26061
rect 35726 26042 35746 26061
rect 35746 26042 35760 26061
rect 35816 26042 35836 26061
rect 35836 26042 35850 26061
rect 35906 26042 35926 26061
rect 35926 26042 35940 26061
rect 35996 26042 36016 26061
rect 36016 26042 36030 26061
rect 36086 26042 36106 26061
rect 36106 26042 36120 26061
rect 36176 26042 36210 26076
rect 36346 26042 36380 26076
rect 36436 26061 36470 26076
rect 36526 26061 36560 26076
rect 36616 26061 36650 26076
rect 36706 26061 36740 26076
rect 36796 26061 36830 26076
rect 36886 26061 36920 26076
rect 36976 26061 37010 26076
rect 37066 26061 37100 26076
rect 37156 26061 37190 26076
rect 37246 26061 37280 26076
rect 37336 26061 37370 26076
rect 37426 26061 37460 26076
rect 36436 26042 36456 26061
rect 36456 26042 36470 26061
rect 36526 26042 36546 26061
rect 36546 26042 36560 26061
rect 36616 26042 36636 26061
rect 36636 26042 36650 26061
rect 36706 26042 36726 26061
rect 36726 26042 36740 26061
rect 36796 26042 36816 26061
rect 36816 26042 36830 26061
rect 36886 26042 36906 26061
rect 36906 26042 36920 26061
rect 36976 26042 36996 26061
rect 36996 26042 37010 26061
rect 37066 26042 37086 26061
rect 37086 26042 37100 26061
rect 37156 26042 37176 26061
rect 37176 26042 37190 26061
rect 37246 26042 37266 26061
rect 37266 26042 37280 26061
rect 37336 26042 37356 26061
rect 37356 26042 37370 26061
rect 37426 26042 37446 26061
rect 37446 26042 37460 26061
rect 37516 26042 37550 26076
rect 37686 26042 37720 26076
rect 37776 26061 37810 26076
rect 37866 26061 37900 26076
rect 37956 26061 37990 26076
rect 38046 26061 38080 26076
rect 38136 26061 38170 26076
rect 38226 26061 38260 26076
rect 38316 26061 38350 26076
rect 38406 26061 38440 26076
rect 38496 26061 38530 26076
rect 38586 26061 38620 26076
rect 38676 26061 38710 26076
rect 38766 26061 38800 26076
rect 37776 26042 37796 26061
rect 37796 26042 37810 26061
rect 37866 26042 37886 26061
rect 37886 26042 37900 26061
rect 37956 26042 37976 26061
rect 37976 26042 37990 26061
rect 38046 26042 38066 26061
rect 38066 26042 38080 26061
rect 38136 26042 38156 26061
rect 38156 26042 38170 26061
rect 38226 26042 38246 26061
rect 38246 26042 38260 26061
rect 38316 26042 38336 26061
rect 38336 26042 38350 26061
rect 38406 26042 38426 26061
rect 38426 26042 38440 26061
rect 38496 26042 38516 26061
rect 38516 26042 38530 26061
rect 38586 26042 38606 26061
rect 38606 26042 38620 26061
rect 38676 26042 38696 26061
rect 38696 26042 38710 26061
rect 38766 26042 38786 26061
rect 38786 26042 38800 26061
rect 38856 26042 38890 26076
rect 15085 25891 15119 25903
rect 15085 25835 15119 25853
rect 15085 25819 15119 25835
rect 15085 25767 15119 25781
rect 15085 25747 15119 25767
rect 15085 25699 15119 25709
rect 15085 25675 15119 25699
rect 15085 25631 15119 25637
rect 15085 25603 15119 25631
rect 15085 25563 15119 25565
rect 15085 25531 15119 25563
rect 15085 25461 15119 25493
rect 15085 25459 15119 25461
rect 15085 25393 15119 25421
rect 15085 25387 15119 25393
rect 15085 25325 15119 25349
rect 15085 25315 15119 25325
rect 15085 25257 15119 25277
rect 15085 25243 15119 25257
rect 15085 25189 15119 25205
rect 15085 25171 15119 25189
rect 22980 25869 23014 25889
rect 22980 25855 23014 25869
rect 22980 25801 23014 25817
rect 22980 25783 23014 25801
rect 22980 25733 23014 25745
rect 22980 25711 23014 25733
rect 22980 25665 23014 25673
rect 22980 25639 23014 25665
rect 22980 25597 23014 25601
rect 22980 25567 23014 25597
rect 22980 25495 23014 25529
rect 22980 25427 23014 25457
rect 22980 25423 23014 25427
rect 22980 25359 23014 25385
rect 22980 25351 23014 25359
rect 22980 25291 23014 25313
rect 22980 25279 23014 25291
rect 22980 25223 23014 25241
rect 22980 25207 23014 25223
rect 15085 25121 15119 25133
rect 15085 25099 15119 25121
rect 15085 25053 15119 25061
rect 15085 25027 15119 25053
rect 22980 25155 23014 25169
rect 22980 25135 23014 25155
rect 23438 25869 23472 25889
rect 23438 25855 23472 25869
rect 23438 25801 23472 25817
rect 23438 25783 23472 25801
rect 23438 25733 23472 25745
rect 23438 25711 23472 25733
rect 23438 25665 23472 25673
rect 23438 25639 23472 25665
rect 23438 25597 23472 25601
rect 23438 25567 23472 25597
rect 23438 25495 23472 25529
rect 23438 25427 23472 25457
rect 23438 25423 23472 25427
rect 23438 25359 23472 25385
rect 23438 25351 23472 25359
rect 23438 25291 23472 25313
rect 23438 25279 23472 25291
rect 23438 25223 23472 25241
rect 23438 25207 23472 25223
rect 23438 25155 23472 25169
rect 23896 25869 23930 25889
rect 23896 25855 23930 25869
rect 23896 25801 23930 25817
rect 23896 25783 23930 25801
rect 23896 25733 23930 25745
rect 23896 25711 23930 25733
rect 23896 25665 23930 25673
rect 23896 25639 23930 25665
rect 23896 25597 23930 25601
rect 23896 25567 23930 25597
rect 23896 25495 23930 25529
rect 23896 25427 23930 25457
rect 23896 25423 23930 25427
rect 23896 25359 23930 25385
rect 23896 25351 23930 25359
rect 23896 25291 23930 25313
rect 23896 25279 23930 25291
rect 23896 25223 23930 25241
rect 23896 25207 23930 25223
rect 23438 25135 23472 25155
rect 23896 25155 23930 25169
rect 23896 25135 23930 25155
rect 24354 25869 24388 25889
rect 24354 25855 24388 25869
rect 24354 25801 24388 25817
rect 24354 25783 24388 25801
rect 24354 25733 24388 25745
rect 24354 25711 24388 25733
rect 24354 25665 24388 25673
rect 24354 25639 24388 25665
rect 24354 25597 24388 25601
rect 24354 25567 24388 25597
rect 24354 25495 24388 25529
rect 24354 25427 24388 25457
rect 24354 25423 24388 25427
rect 24354 25359 24388 25385
rect 24354 25351 24388 25359
rect 24354 25291 24388 25313
rect 24354 25279 24388 25291
rect 24354 25223 24388 25241
rect 24354 25207 24388 25223
rect 24354 25155 24388 25169
rect 24812 25869 24846 25889
rect 24812 25855 24846 25869
rect 24812 25801 24846 25817
rect 24812 25783 24846 25801
rect 24812 25733 24846 25745
rect 24812 25711 24846 25733
rect 24812 25665 24846 25673
rect 24812 25639 24846 25665
rect 24812 25597 24846 25601
rect 24812 25567 24846 25597
rect 24812 25495 24846 25529
rect 24812 25427 24846 25457
rect 24812 25423 24846 25427
rect 24812 25359 24846 25385
rect 24812 25351 24846 25359
rect 24812 25291 24846 25313
rect 24812 25279 24846 25291
rect 24812 25223 24846 25241
rect 24812 25207 24846 25223
rect 24354 25135 24388 25155
rect 24812 25155 24846 25169
rect 24812 25135 24846 25155
rect 25270 25869 25304 25889
rect 25270 25855 25304 25869
rect 25270 25801 25304 25817
rect 25270 25783 25304 25801
rect 25270 25733 25304 25745
rect 25270 25711 25304 25733
rect 25270 25665 25304 25673
rect 25270 25639 25304 25665
rect 25270 25597 25304 25601
rect 25270 25567 25304 25597
rect 25270 25495 25304 25529
rect 25270 25427 25304 25457
rect 25270 25423 25304 25427
rect 25270 25359 25304 25385
rect 25270 25351 25304 25359
rect 25270 25291 25304 25313
rect 25270 25279 25304 25291
rect 25270 25223 25304 25241
rect 25270 25207 25304 25223
rect 25270 25155 25304 25169
rect 25728 25869 25762 25889
rect 25728 25855 25762 25869
rect 25728 25801 25762 25817
rect 25728 25783 25762 25801
rect 25728 25733 25762 25745
rect 25728 25711 25762 25733
rect 25728 25665 25762 25673
rect 25728 25639 25762 25665
rect 25728 25597 25762 25601
rect 25728 25567 25762 25597
rect 25728 25495 25762 25529
rect 25728 25427 25762 25457
rect 25728 25423 25762 25427
rect 25728 25359 25762 25385
rect 25728 25351 25762 25359
rect 25728 25291 25762 25313
rect 25728 25279 25762 25291
rect 25728 25223 25762 25241
rect 25728 25207 25762 25223
rect 25270 25135 25304 25155
rect 25728 25155 25762 25169
rect 25728 25135 25762 25155
rect 26186 25869 26220 25889
rect 26186 25855 26220 25869
rect 26186 25801 26220 25817
rect 26186 25783 26220 25801
rect 26186 25733 26220 25745
rect 26186 25711 26220 25733
rect 26186 25665 26220 25673
rect 26186 25639 26220 25665
rect 26186 25597 26220 25601
rect 26186 25567 26220 25597
rect 26186 25495 26220 25529
rect 26186 25427 26220 25457
rect 26186 25423 26220 25427
rect 26186 25359 26220 25385
rect 26186 25351 26220 25359
rect 26186 25291 26220 25313
rect 26186 25279 26220 25291
rect 26186 25223 26220 25241
rect 26186 25207 26220 25223
rect 26186 25155 26220 25169
rect 26644 25869 26678 25889
rect 26644 25855 26678 25869
rect 26644 25801 26678 25817
rect 26644 25783 26678 25801
rect 26644 25733 26678 25745
rect 26644 25711 26678 25733
rect 26644 25665 26678 25673
rect 26644 25639 26678 25665
rect 26644 25597 26678 25601
rect 26644 25567 26678 25597
rect 26644 25495 26678 25529
rect 26644 25427 26678 25457
rect 26644 25423 26678 25427
rect 26644 25359 26678 25385
rect 26644 25351 26678 25359
rect 26644 25291 26678 25313
rect 26644 25279 26678 25291
rect 26644 25223 26678 25241
rect 26644 25207 26678 25223
rect 26186 25135 26220 25155
rect 26644 25155 26678 25169
rect 26644 25135 26678 25155
rect 27102 25869 27136 25889
rect 27102 25855 27136 25869
rect 27102 25801 27136 25817
rect 27102 25783 27136 25801
rect 27102 25733 27136 25745
rect 27102 25711 27136 25733
rect 27102 25665 27136 25673
rect 27102 25639 27136 25665
rect 27102 25597 27136 25601
rect 27102 25567 27136 25597
rect 27102 25495 27136 25529
rect 27102 25427 27136 25457
rect 27102 25423 27136 25427
rect 27102 25359 27136 25385
rect 27102 25351 27136 25359
rect 27102 25291 27136 25313
rect 27102 25279 27136 25291
rect 27102 25223 27136 25241
rect 27102 25207 27136 25223
rect 27102 25155 27136 25169
rect 27102 25135 27136 25155
rect 15085 24985 15119 24989
rect 15085 24955 15119 24985
rect 23397 24973 23431 25007
rect 15085 24883 15119 24917
rect 28470 25882 28504 25916
rect 28560 25914 28594 25916
rect 28650 25914 28684 25916
rect 28740 25914 28774 25916
rect 28830 25914 28864 25916
rect 28920 25914 28954 25916
rect 29010 25914 29044 25916
rect 29100 25914 29134 25916
rect 29190 25914 29224 25916
rect 29280 25914 29314 25916
rect 28560 25882 28580 25914
rect 28580 25882 28594 25914
rect 28650 25882 28670 25914
rect 28670 25882 28684 25914
rect 28740 25882 28760 25914
rect 28760 25882 28774 25914
rect 28830 25882 28850 25914
rect 28850 25882 28864 25914
rect 28920 25882 28940 25914
rect 28940 25882 28954 25914
rect 29010 25882 29030 25914
rect 29030 25882 29044 25914
rect 29100 25882 29120 25914
rect 29120 25882 29134 25914
rect 29190 25882 29210 25914
rect 29210 25882 29224 25914
rect 29280 25882 29300 25914
rect 29300 25882 29314 25914
rect 29370 25882 29404 25916
rect 28656 25706 28678 25712
rect 28678 25706 28690 25712
rect 28756 25706 28768 25712
rect 28768 25706 28790 25712
rect 28856 25706 28858 25712
rect 28858 25706 28890 25712
rect 28656 25678 28690 25706
rect 28756 25678 28790 25706
rect 28856 25678 28890 25706
rect 28956 25678 28990 25712
rect 29056 25678 29090 25712
rect 29156 25706 29184 25712
rect 29184 25706 29190 25712
rect 29156 25678 29190 25706
rect 28656 25578 28690 25612
rect 28756 25578 28790 25612
rect 28856 25578 28890 25612
rect 28956 25578 28990 25612
rect 29056 25578 29090 25612
rect 29156 25578 29190 25612
rect 28656 25478 28690 25512
rect 28756 25478 28790 25512
rect 28856 25478 28890 25512
rect 28956 25478 28990 25512
rect 29056 25478 29090 25512
rect 29156 25478 29190 25512
rect 28656 25380 28690 25412
rect 28756 25380 28790 25412
rect 28856 25380 28890 25412
rect 28656 25378 28678 25380
rect 28678 25378 28690 25380
rect 28756 25378 28768 25380
rect 28768 25378 28790 25380
rect 28856 25378 28858 25380
rect 28858 25378 28890 25380
rect 28956 25378 28990 25412
rect 29056 25378 29090 25412
rect 29156 25380 29190 25412
rect 29156 25378 29184 25380
rect 29184 25378 29190 25380
rect 28656 25290 28690 25312
rect 28756 25290 28790 25312
rect 28856 25290 28890 25312
rect 28656 25278 28678 25290
rect 28678 25278 28690 25290
rect 28756 25278 28768 25290
rect 28768 25278 28790 25290
rect 28856 25278 28858 25290
rect 28858 25278 28890 25290
rect 28956 25278 28990 25312
rect 29056 25278 29090 25312
rect 29156 25290 29190 25312
rect 29156 25278 29184 25290
rect 29184 25278 29190 25290
rect 28656 25200 28690 25212
rect 28756 25200 28790 25212
rect 28856 25200 28890 25212
rect 28656 25178 28678 25200
rect 28678 25178 28690 25200
rect 28756 25178 28768 25200
rect 28768 25178 28790 25200
rect 28856 25178 28858 25200
rect 28858 25178 28890 25200
rect 28956 25178 28990 25212
rect 29056 25178 29090 25212
rect 29156 25200 29190 25212
rect 29156 25178 29184 25200
rect 29184 25178 29190 25200
rect 29810 25882 29844 25916
rect 29900 25914 29934 25916
rect 29990 25914 30024 25916
rect 30080 25914 30114 25916
rect 30170 25914 30204 25916
rect 30260 25914 30294 25916
rect 30350 25914 30384 25916
rect 30440 25914 30474 25916
rect 30530 25914 30564 25916
rect 30620 25914 30654 25916
rect 29900 25882 29920 25914
rect 29920 25882 29934 25914
rect 29990 25882 30010 25914
rect 30010 25882 30024 25914
rect 30080 25882 30100 25914
rect 30100 25882 30114 25914
rect 30170 25882 30190 25914
rect 30190 25882 30204 25914
rect 30260 25882 30280 25914
rect 30280 25882 30294 25914
rect 30350 25882 30370 25914
rect 30370 25882 30384 25914
rect 30440 25882 30460 25914
rect 30460 25882 30474 25914
rect 30530 25882 30550 25914
rect 30550 25882 30564 25914
rect 30620 25882 30640 25914
rect 30640 25882 30654 25914
rect 30710 25882 30744 25916
rect 29996 25706 30018 25712
rect 30018 25706 30030 25712
rect 30096 25706 30108 25712
rect 30108 25706 30130 25712
rect 30196 25706 30198 25712
rect 30198 25706 30230 25712
rect 29996 25678 30030 25706
rect 30096 25678 30130 25706
rect 30196 25678 30230 25706
rect 30296 25678 30330 25712
rect 30396 25678 30430 25712
rect 30496 25706 30524 25712
rect 30524 25706 30530 25712
rect 30496 25678 30530 25706
rect 29996 25578 30030 25612
rect 30096 25578 30130 25612
rect 30196 25578 30230 25612
rect 30296 25578 30330 25612
rect 30396 25578 30430 25612
rect 30496 25578 30530 25612
rect 29996 25478 30030 25512
rect 30096 25478 30130 25512
rect 30196 25478 30230 25512
rect 30296 25478 30330 25512
rect 30396 25478 30430 25512
rect 30496 25478 30530 25512
rect 29996 25380 30030 25412
rect 30096 25380 30130 25412
rect 30196 25380 30230 25412
rect 29996 25378 30018 25380
rect 30018 25378 30030 25380
rect 30096 25378 30108 25380
rect 30108 25378 30130 25380
rect 30196 25378 30198 25380
rect 30198 25378 30230 25380
rect 30296 25378 30330 25412
rect 30396 25378 30430 25412
rect 30496 25380 30530 25412
rect 30496 25378 30524 25380
rect 30524 25378 30530 25380
rect 29996 25290 30030 25312
rect 30096 25290 30130 25312
rect 30196 25290 30230 25312
rect 29996 25278 30018 25290
rect 30018 25278 30030 25290
rect 30096 25278 30108 25290
rect 30108 25278 30130 25290
rect 30196 25278 30198 25290
rect 30198 25278 30230 25290
rect 30296 25278 30330 25312
rect 30396 25278 30430 25312
rect 30496 25290 30530 25312
rect 30496 25278 30524 25290
rect 30524 25278 30530 25290
rect 29996 25200 30030 25212
rect 30096 25200 30130 25212
rect 30196 25200 30230 25212
rect 29996 25178 30018 25200
rect 30018 25178 30030 25200
rect 30096 25178 30108 25200
rect 30108 25178 30130 25200
rect 30196 25178 30198 25200
rect 30198 25178 30230 25200
rect 30296 25178 30330 25212
rect 30396 25178 30430 25212
rect 30496 25200 30530 25212
rect 30496 25178 30524 25200
rect 30524 25178 30530 25200
rect 31150 25882 31184 25916
rect 31240 25914 31274 25916
rect 31330 25914 31364 25916
rect 31420 25914 31454 25916
rect 31510 25914 31544 25916
rect 31600 25914 31634 25916
rect 31690 25914 31724 25916
rect 31780 25914 31814 25916
rect 31870 25914 31904 25916
rect 31960 25914 31994 25916
rect 31240 25882 31260 25914
rect 31260 25882 31274 25914
rect 31330 25882 31350 25914
rect 31350 25882 31364 25914
rect 31420 25882 31440 25914
rect 31440 25882 31454 25914
rect 31510 25882 31530 25914
rect 31530 25882 31544 25914
rect 31600 25882 31620 25914
rect 31620 25882 31634 25914
rect 31690 25882 31710 25914
rect 31710 25882 31724 25914
rect 31780 25882 31800 25914
rect 31800 25882 31814 25914
rect 31870 25882 31890 25914
rect 31890 25882 31904 25914
rect 31960 25882 31980 25914
rect 31980 25882 31994 25914
rect 32050 25882 32084 25916
rect 31336 25706 31358 25712
rect 31358 25706 31370 25712
rect 31436 25706 31448 25712
rect 31448 25706 31470 25712
rect 31536 25706 31538 25712
rect 31538 25706 31570 25712
rect 31336 25678 31370 25706
rect 31436 25678 31470 25706
rect 31536 25678 31570 25706
rect 31636 25678 31670 25712
rect 31736 25678 31770 25712
rect 31836 25706 31864 25712
rect 31864 25706 31870 25712
rect 31836 25678 31870 25706
rect 31336 25578 31370 25612
rect 31436 25578 31470 25612
rect 31536 25578 31570 25612
rect 31636 25578 31670 25612
rect 31736 25578 31770 25612
rect 31836 25578 31870 25612
rect 31336 25478 31370 25512
rect 31436 25478 31470 25512
rect 31536 25478 31570 25512
rect 31636 25478 31670 25512
rect 31736 25478 31770 25512
rect 31836 25478 31870 25512
rect 31336 25380 31370 25412
rect 31436 25380 31470 25412
rect 31536 25380 31570 25412
rect 31336 25378 31358 25380
rect 31358 25378 31370 25380
rect 31436 25378 31448 25380
rect 31448 25378 31470 25380
rect 31536 25378 31538 25380
rect 31538 25378 31570 25380
rect 31636 25378 31670 25412
rect 31736 25378 31770 25412
rect 31836 25380 31870 25412
rect 31836 25378 31864 25380
rect 31864 25378 31870 25380
rect 31336 25290 31370 25312
rect 31436 25290 31470 25312
rect 31536 25290 31570 25312
rect 31336 25278 31358 25290
rect 31358 25278 31370 25290
rect 31436 25278 31448 25290
rect 31448 25278 31470 25290
rect 31536 25278 31538 25290
rect 31538 25278 31570 25290
rect 31636 25278 31670 25312
rect 31736 25278 31770 25312
rect 31836 25290 31870 25312
rect 31836 25278 31864 25290
rect 31864 25278 31870 25290
rect 31336 25200 31370 25212
rect 31436 25200 31470 25212
rect 31536 25200 31570 25212
rect 31336 25178 31358 25200
rect 31358 25178 31370 25200
rect 31436 25178 31448 25200
rect 31448 25178 31470 25200
rect 31536 25178 31538 25200
rect 31538 25178 31570 25200
rect 31636 25178 31670 25212
rect 31736 25178 31770 25212
rect 31836 25200 31870 25212
rect 31836 25178 31864 25200
rect 31864 25178 31870 25200
rect 32490 25882 32524 25916
rect 32580 25914 32614 25916
rect 32670 25914 32704 25916
rect 32760 25914 32794 25916
rect 32850 25914 32884 25916
rect 32940 25914 32974 25916
rect 33030 25914 33064 25916
rect 33120 25914 33154 25916
rect 33210 25914 33244 25916
rect 33300 25914 33334 25916
rect 32580 25882 32600 25914
rect 32600 25882 32614 25914
rect 32670 25882 32690 25914
rect 32690 25882 32704 25914
rect 32760 25882 32780 25914
rect 32780 25882 32794 25914
rect 32850 25882 32870 25914
rect 32870 25882 32884 25914
rect 32940 25882 32960 25914
rect 32960 25882 32974 25914
rect 33030 25882 33050 25914
rect 33050 25882 33064 25914
rect 33120 25882 33140 25914
rect 33140 25882 33154 25914
rect 33210 25882 33230 25914
rect 33230 25882 33244 25914
rect 33300 25882 33320 25914
rect 33320 25882 33334 25914
rect 33390 25882 33424 25916
rect 32676 25706 32698 25712
rect 32698 25706 32710 25712
rect 32776 25706 32788 25712
rect 32788 25706 32810 25712
rect 32876 25706 32878 25712
rect 32878 25706 32910 25712
rect 32676 25678 32710 25706
rect 32776 25678 32810 25706
rect 32876 25678 32910 25706
rect 32976 25678 33010 25712
rect 33076 25678 33110 25712
rect 33176 25706 33204 25712
rect 33204 25706 33210 25712
rect 33176 25678 33210 25706
rect 32676 25578 32710 25612
rect 32776 25578 32810 25612
rect 32876 25578 32910 25612
rect 32976 25578 33010 25612
rect 33076 25578 33110 25612
rect 33176 25578 33210 25612
rect 32676 25478 32710 25512
rect 32776 25478 32810 25512
rect 32876 25478 32910 25512
rect 32976 25478 33010 25512
rect 33076 25478 33110 25512
rect 33176 25478 33210 25512
rect 32676 25380 32710 25412
rect 32776 25380 32810 25412
rect 32876 25380 32910 25412
rect 32676 25378 32698 25380
rect 32698 25378 32710 25380
rect 32776 25378 32788 25380
rect 32788 25378 32810 25380
rect 32876 25378 32878 25380
rect 32878 25378 32910 25380
rect 32976 25378 33010 25412
rect 33076 25378 33110 25412
rect 33176 25380 33210 25412
rect 33176 25378 33204 25380
rect 33204 25378 33210 25380
rect 32676 25290 32710 25312
rect 32776 25290 32810 25312
rect 32876 25290 32910 25312
rect 32676 25278 32698 25290
rect 32698 25278 32710 25290
rect 32776 25278 32788 25290
rect 32788 25278 32810 25290
rect 32876 25278 32878 25290
rect 32878 25278 32910 25290
rect 32976 25278 33010 25312
rect 33076 25278 33110 25312
rect 33176 25290 33210 25312
rect 33176 25278 33204 25290
rect 33204 25278 33210 25290
rect 32676 25200 32710 25212
rect 32776 25200 32810 25212
rect 32876 25200 32910 25212
rect 32676 25178 32698 25200
rect 32698 25178 32710 25200
rect 32776 25178 32788 25200
rect 32788 25178 32810 25200
rect 32876 25178 32878 25200
rect 32878 25178 32910 25200
rect 32976 25178 33010 25212
rect 33076 25178 33110 25212
rect 33176 25200 33210 25212
rect 33176 25178 33204 25200
rect 33204 25178 33210 25200
rect 33830 25882 33864 25916
rect 33920 25914 33954 25916
rect 34010 25914 34044 25916
rect 34100 25914 34134 25916
rect 34190 25914 34224 25916
rect 34280 25914 34314 25916
rect 34370 25914 34404 25916
rect 34460 25914 34494 25916
rect 34550 25914 34584 25916
rect 34640 25914 34674 25916
rect 33920 25882 33940 25914
rect 33940 25882 33954 25914
rect 34010 25882 34030 25914
rect 34030 25882 34044 25914
rect 34100 25882 34120 25914
rect 34120 25882 34134 25914
rect 34190 25882 34210 25914
rect 34210 25882 34224 25914
rect 34280 25882 34300 25914
rect 34300 25882 34314 25914
rect 34370 25882 34390 25914
rect 34390 25882 34404 25914
rect 34460 25882 34480 25914
rect 34480 25882 34494 25914
rect 34550 25882 34570 25914
rect 34570 25882 34584 25914
rect 34640 25882 34660 25914
rect 34660 25882 34674 25914
rect 34730 25882 34764 25916
rect 34016 25706 34038 25712
rect 34038 25706 34050 25712
rect 34116 25706 34128 25712
rect 34128 25706 34150 25712
rect 34216 25706 34218 25712
rect 34218 25706 34250 25712
rect 34016 25678 34050 25706
rect 34116 25678 34150 25706
rect 34216 25678 34250 25706
rect 34316 25678 34350 25712
rect 34416 25678 34450 25712
rect 34516 25706 34544 25712
rect 34544 25706 34550 25712
rect 34516 25678 34550 25706
rect 34016 25578 34050 25612
rect 34116 25578 34150 25612
rect 34216 25578 34250 25612
rect 34316 25578 34350 25612
rect 34416 25578 34450 25612
rect 34516 25578 34550 25612
rect 34016 25478 34050 25512
rect 34116 25478 34150 25512
rect 34216 25478 34250 25512
rect 34316 25478 34350 25512
rect 34416 25478 34450 25512
rect 34516 25478 34550 25512
rect 34016 25380 34050 25412
rect 34116 25380 34150 25412
rect 34216 25380 34250 25412
rect 34016 25378 34038 25380
rect 34038 25378 34050 25380
rect 34116 25378 34128 25380
rect 34128 25378 34150 25380
rect 34216 25378 34218 25380
rect 34218 25378 34250 25380
rect 34316 25378 34350 25412
rect 34416 25378 34450 25412
rect 34516 25380 34550 25412
rect 34516 25378 34544 25380
rect 34544 25378 34550 25380
rect 34016 25290 34050 25312
rect 34116 25290 34150 25312
rect 34216 25290 34250 25312
rect 34016 25278 34038 25290
rect 34038 25278 34050 25290
rect 34116 25278 34128 25290
rect 34128 25278 34150 25290
rect 34216 25278 34218 25290
rect 34218 25278 34250 25290
rect 34316 25278 34350 25312
rect 34416 25278 34450 25312
rect 34516 25290 34550 25312
rect 34516 25278 34544 25290
rect 34544 25278 34550 25290
rect 34016 25200 34050 25212
rect 34116 25200 34150 25212
rect 34216 25200 34250 25212
rect 34016 25178 34038 25200
rect 34038 25178 34050 25200
rect 34116 25178 34128 25200
rect 34128 25178 34150 25200
rect 34216 25178 34218 25200
rect 34218 25178 34250 25200
rect 34316 25178 34350 25212
rect 34416 25178 34450 25212
rect 34516 25200 34550 25212
rect 34516 25178 34544 25200
rect 34544 25178 34550 25200
rect 35170 25882 35204 25916
rect 35260 25914 35294 25916
rect 35350 25914 35384 25916
rect 35440 25914 35474 25916
rect 35530 25914 35564 25916
rect 35620 25914 35654 25916
rect 35710 25914 35744 25916
rect 35800 25914 35834 25916
rect 35890 25914 35924 25916
rect 35980 25914 36014 25916
rect 35260 25882 35280 25914
rect 35280 25882 35294 25914
rect 35350 25882 35370 25914
rect 35370 25882 35384 25914
rect 35440 25882 35460 25914
rect 35460 25882 35474 25914
rect 35530 25882 35550 25914
rect 35550 25882 35564 25914
rect 35620 25882 35640 25914
rect 35640 25882 35654 25914
rect 35710 25882 35730 25914
rect 35730 25882 35744 25914
rect 35800 25882 35820 25914
rect 35820 25882 35834 25914
rect 35890 25882 35910 25914
rect 35910 25882 35924 25914
rect 35980 25882 36000 25914
rect 36000 25882 36014 25914
rect 36070 25882 36104 25916
rect 35356 25706 35378 25712
rect 35378 25706 35390 25712
rect 35456 25706 35468 25712
rect 35468 25706 35490 25712
rect 35556 25706 35558 25712
rect 35558 25706 35590 25712
rect 35356 25678 35390 25706
rect 35456 25678 35490 25706
rect 35556 25678 35590 25706
rect 35656 25678 35690 25712
rect 35756 25678 35790 25712
rect 35856 25706 35884 25712
rect 35884 25706 35890 25712
rect 35856 25678 35890 25706
rect 35356 25578 35390 25612
rect 35456 25578 35490 25612
rect 35556 25578 35590 25612
rect 35656 25578 35690 25612
rect 35756 25578 35790 25612
rect 35856 25578 35890 25612
rect 35356 25478 35390 25512
rect 35456 25478 35490 25512
rect 35556 25478 35590 25512
rect 35656 25478 35690 25512
rect 35756 25478 35790 25512
rect 35856 25478 35890 25512
rect 35356 25380 35390 25412
rect 35456 25380 35490 25412
rect 35556 25380 35590 25412
rect 35356 25378 35378 25380
rect 35378 25378 35390 25380
rect 35456 25378 35468 25380
rect 35468 25378 35490 25380
rect 35556 25378 35558 25380
rect 35558 25378 35590 25380
rect 35656 25378 35690 25412
rect 35756 25378 35790 25412
rect 35856 25380 35890 25412
rect 35856 25378 35884 25380
rect 35884 25378 35890 25380
rect 35356 25290 35390 25312
rect 35456 25290 35490 25312
rect 35556 25290 35590 25312
rect 35356 25278 35378 25290
rect 35378 25278 35390 25290
rect 35456 25278 35468 25290
rect 35468 25278 35490 25290
rect 35556 25278 35558 25290
rect 35558 25278 35590 25290
rect 35656 25278 35690 25312
rect 35756 25278 35790 25312
rect 35856 25290 35890 25312
rect 35856 25278 35884 25290
rect 35884 25278 35890 25290
rect 35356 25200 35390 25212
rect 35456 25200 35490 25212
rect 35556 25200 35590 25212
rect 35356 25178 35378 25200
rect 35378 25178 35390 25200
rect 35456 25178 35468 25200
rect 35468 25178 35490 25200
rect 35556 25178 35558 25200
rect 35558 25178 35590 25200
rect 35656 25178 35690 25212
rect 35756 25178 35790 25212
rect 35856 25200 35890 25212
rect 35856 25178 35884 25200
rect 35884 25178 35890 25200
rect 36510 25882 36544 25916
rect 36600 25914 36634 25916
rect 36690 25914 36724 25916
rect 36780 25914 36814 25916
rect 36870 25914 36904 25916
rect 36960 25914 36994 25916
rect 37050 25914 37084 25916
rect 37140 25914 37174 25916
rect 37230 25914 37264 25916
rect 37320 25914 37354 25916
rect 36600 25882 36620 25914
rect 36620 25882 36634 25914
rect 36690 25882 36710 25914
rect 36710 25882 36724 25914
rect 36780 25882 36800 25914
rect 36800 25882 36814 25914
rect 36870 25882 36890 25914
rect 36890 25882 36904 25914
rect 36960 25882 36980 25914
rect 36980 25882 36994 25914
rect 37050 25882 37070 25914
rect 37070 25882 37084 25914
rect 37140 25882 37160 25914
rect 37160 25882 37174 25914
rect 37230 25882 37250 25914
rect 37250 25882 37264 25914
rect 37320 25882 37340 25914
rect 37340 25882 37354 25914
rect 37410 25882 37444 25916
rect 36696 25706 36718 25712
rect 36718 25706 36730 25712
rect 36796 25706 36808 25712
rect 36808 25706 36830 25712
rect 36896 25706 36898 25712
rect 36898 25706 36930 25712
rect 36696 25678 36730 25706
rect 36796 25678 36830 25706
rect 36896 25678 36930 25706
rect 36996 25678 37030 25712
rect 37096 25678 37130 25712
rect 37196 25706 37224 25712
rect 37224 25706 37230 25712
rect 37196 25678 37230 25706
rect 36696 25578 36730 25612
rect 36796 25578 36830 25612
rect 36896 25578 36930 25612
rect 36996 25578 37030 25612
rect 37096 25578 37130 25612
rect 37196 25578 37230 25612
rect 36696 25478 36730 25512
rect 36796 25478 36830 25512
rect 36896 25478 36930 25512
rect 36996 25478 37030 25512
rect 37096 25478 37130 25512
rect 37196 25478 37230 25512
rect 36696 25380 36730 25412
rect 36796 25380 36830 25412
rect 36896 25380 36930 25412
rect 36696 25378 36718 25380
rect 36718 25378 36730 25380
rect 36796 25378 36808 25380
rect 36808 25378 36830 25380
rect 36896 25378 36898 25380
rect 36898 25378 36930 25380
rect 36996 25378 37030 25412
rect 37096 25378 37130 25412
rect 37196 25380 37230 25412
rect 37196 25378 37224 25380
rect 37224 25378 37230 25380
rect 36696 25290 36730 25312
rect 36796 25290 36830 25312
rect 36896 25290 36930 25312
rect 36696 25278 36718 25290
rect 36718 25278 36730 25290
rect 36796 25278 36808 25290
rect 36808 25278 36830 25290
rect 36896 25278 36898 25290
rect 36898 25278 36930 25290
rect 36996 25278 37030 25312
rect 37096 25278 37130 25312
rect 37196 25290 37230 25312
rect 37196 25278 37224 25290
rect 37224 25278 37230 25290
rect 36696 25200 36730 25212
rect 36796 25200 36830 25212
rect 36896 25200 36930 25212
rect 36696 25178 36718 25200
rect 36718 25178 36730 25200
rect 36796 25178 36808 25200
rect 36808 25178 36830 25200
rect 36896 25178 36898 25200
rect 36898 25178 36930 25200
rect 36996 25178 37030 25212
rect 37096 25178 37130 25212
rect 37196 25200 37230 25212
rect 37196 25178 37224 25200
rect 37224 25178 37230 25200
rect 37850 25882 37884 25916
rect 37940 25914 37974 25916
rect 38030 25914 38064 25916
rect 38120 25914 38154 25916
rect 38210 25914 38244 25916
rect 38300 25914 38334 25916
rect 38390 25914 38424 25916
rect 38480 25914 38514 25916
rect 38570 25914 38604 25916
rect 38660 25914 38694 25916
rect 37940 25882 37960 25914
rect 37960 25882 37974 25914
rect 38030 25882 38050 25914
rect 38050 25882 38064 25914
rect 38120 25882 38140 25914
rect 38140 25882 38154 25914
rect 38210 25882 38230 25914
rect 38230 25882 38244 25914
rect 38300 25882 38320 25914
rect 38320 25882 38334 25914
rect 38390 25882 38410 25914
rect 38410 25882 38424 25914
rect 38480 25882 38500 25914
rect 38500 25882 38514 25914
rect 38570 25882 38590 25914
rect 38590 25882 38604 25914
rect 38660 25882 38680 25914
rect 38680 25882 38694 25914
rect 38750 25882 38784 25916
rect 38036 25706 38058 25712
rect 38058 25706 38070 25712
rect 38136 25706 38148 25712
rect 38148 25706 38170 25712
rect 38236 25706 38238 25712
rect 38238 25706 38270 25712
rect 38036 25678 38070 25706
rect 38136 25678 38170 25706
rect 38236 25678 38270 25706
rect 38336 25678 38370 25712
rect 38436 25678 38470 25712
rect 38536 25706 38564 25712
rect 38564 25706 38570 25712
rect 38536 25678 38570 25706
rect 38036 25578 38070 25612
rect 38136 25578 38170 25612
rect 38236 25578 38270 25612
rect 38336 25578 38370 25612
rect 38436 25578 38470 25612
rect 38536 25578 38570 25612
rect 38036 25478 38070 25512
rect 38136 25478 38170 25512
rect 38236 25478 38270 25512
rect 38336 25478 38370 25512
rect 38436 25478 38470 25512
rect 38536 25478 38570 25512
rect 38036 25380 38070 25412
rect 38136 25380 38170 25412
rect 38236 25380 38270 25412
rect 38036 25378 38058 25380
rect 38058 25378 38070 25380
rect 38136 25378 38148 25380
rect 38148 25378 38170 25380
rect 38236 25378 38238 25380
rect 38238 25378 38270 25380
rect 38336 25378 38370 25412
rect 38436 25378 38470 25412
rect 38536 25380 38570 25412
rect 38536 25378 38564 25380
rect 38564 25378 38570 25380
rect 38036 25290 38070 25312
rect 38136 25290 38170 25312
rect 38236 25290 38270 25312
rect 38036 25278 38058 25290
rect 38058 25278 38070 25290
rect 38136 25278 38148 25290
rect 38148 25278 38170 25290
rect 38236 25278 38238 25290
rect 38238 25278 38270 25290
rect 38336 25278 38370 25312
rect 38436 25278 38470 25312
rect 38536 25290 38570 25312
rect 38536 25278 38564 25290
rect 38564 25278 38570 25290
rect 38036 25200 38070 25212
rect 38136 25200 38170 25212
rect 38236 25200 38270 25212
rect 38036 25178 38058 25200
rect 38058 25178 38070 25200
rect 38136 25178 38148 25200
rect 38148 25178 38170 25200
rect 38236 25178 38238 25200
rect 38238 25178 38270 25200
rect 38336 25178 38370 25212
rect 38436 25178 38470 25212
rect 38536 25200 38570 25212
rect 38536 25178 38564 25200
rect 38564 25178 38570 25200
rect 39765 25603 40159 26141
rect 41772 25603 42166 26141
rect 23305 24837 23339 24871
rect 9689 24633 9723 24667
rect 12541 24663 12575 24667
rect 12541 24633 12559 24663
rect 12559 24633 12575 24663
rect 39765 24643 40159 25181
rect 41772 24643 42166 25181
rect 6903 24495 6937 24529
rect 7103 24495 7137 24529
rect 7303 24495 7337 24529
rect 7503 24495 7537 24529
rect 7703 24495 7737 24529
rect 7903 24495 7937 24529
rect 8103 24495 8137 24529
rect 8303 24495 8337 24529
rect 8503 24495 8537 24529
rect 8703 24495 8737 24529
rect 8903 24495 8937 24529
rect 9725 24495 9759 24529
rect 10125 24495 10159 24529
rect 10525 24495 10559 24529
rect 10925 24495 10959 24529
rect 11325 24495 11359 24529
rect 11725 24495 11759 24529
rect 12125 24495 12159 24529
rect 12525 24495 12559 24529
rect 12925 24495 12959 24529
rect 13325 24495 13359 24529
rect 13725 24495 13759 24529
rect 14125 24495 14159 24529
rect 14525 24495 14559 24529
rect 14925 24495 14959 24529
rect 15607 24495 15641 24529
rect 16007 24495 16041 24529
rect 16407 24495 16441 24529
rect 16807 24495 16841 24529
rect 17207 24495 17241 24529
rect 17607 24495 17641 24529
rect 18007 24495 18041 24529
rect 18407 24495 18441 24529
rect 18807 24495 18841 24529
rect 19207 24495 19241 24529
rect 19607 24495 19641 24529
rect 20007 24495 20041 24529
rect 20407 24495 20441 24529
rect 20807 24495 20841 24529
rect 21207 24495 21241 24529
rect 21607 24495 21641 24529
rect 22007 24495 22041 24529
rect 22407 24495 22441 24529
rect 23151 24495 23185 24529
rect 23551 24495 23585 24529
rect 23951 24495 23985 24529
rect 24351 24495 24385 24529
rect 24751 24495 24785 24529
rect 25151 24495 25185 24529
rect 25551 24495 25585 24529
rect 25951 24495 25985 24529
rect 26351 24495 26385 24529
rect 26751 24495 26785 24529
rect 28443 24495 28477 24529
rect 28643 24495 28677 24529
rect 28843 24495 28877 24529
rect 29043 24495 29077 24529
rect 29243 24495 29277 24529
rect 29443 24495 29477 24529
rect 29643 24495 29677 24529
rect 29843 24495 29877 24529
rect 30043 24495 30077 24529
rect 30243 24495 30277 24529
rect 30443 24495 30477 24529
rect 30643 24495 30677 24529
rect 30843 24495 30877 24529
rect 31043 24495 31077 24529
rect 31243 24495 31277 24529
rect 31443 24495 31477 24529
rect 31643 24495 31677 24529
rect 31843 24495 31877 24529
rect 32043 24495 32077 24529
rect 32243 24495 32277 24529
rect 32443 24495 32477 24529
rect 32643 24495 32677 24529
rect 32843 24495 32877 24529
rect 33043 24495 33077 24529
rect 33243 24495 33277 24529
rect 33443 24495 33477 24529
rect 33643 24495 33677 24529
rect 33843 24495 33877 24529
rect 34043 24495 34077 24529
rect 34243 24495 34277 24529
rect 34443 24495 34477 24529
rect 34643 24495 34677 24529
rect 34843 24495 34877 24529
rect 35043 24495 35077 24529
rect 35243 24495 35277 24529
rect 35443 24495 35477 24529
rect 35643 24495 35677 24529
rect 35843 24495 35877 24529
rect 36043 24495 36077 24529
rect 36243 24495 36277 24529
rect 36443 24495 36477 24529
rect 36643 24495 36677 24529
rect 36843 24495 36877 24529
rect 37043 24495 37077 24529
rect 37243 24495 37277 24529
rect 37443 24495 37477 24529
rect 37643 24495 37677 24529
rect 37843 24495 37877 24529
rect 38043 24495 38077 24529
rect 38243 24495 38277 24529
rect 38443 24495 38477 24529
rect 38643 24495 38677 24529
rect 38843 24495 38877 24529
rect 39929 24495 39963 24529
rect 40129 24495 40163 24529
rect 40329 24495 40363 24529
rect 40529 24495 40563 24529
rect 40729 24495 40763 24529
rect 40929 24495 40963 24529
rect 41129 24495 41163 24529
rect 41329 24495 41363 24529
rect 41529 24495 41563 24529
rect 41729 24495 41763 24529
rect 41929 24495 41963 24529
rect 7863 22615 7897 22649
rect 8263 22615 8297 22649
rect 8663 22615 8697 22649
rect 9063 22615 9097 22649
rect 9463 22615 9497 22649
rect 9863 22615 9897 22649
rect 10263 22615 10297 22649
rect 10663 22615 10697 22649
rect 11063 22615 11097 22649
rect 11463 22615 11497 22649
rect 11863 22615 11897 22649
rect 12263 22615 12297 22649
rect 12663 22615 12697 22649
rect 13063 22615 13097 22649
rect 13745 22615 13779 22649
rect 14145 22615 14179 22649
rect 14545 22615 14579 22649
rect 14945 22615 14979 22649
rect 15345 22615 15379 22649
rect 15745 22615 15779 22649
rect 16145 22615 16179 22649
rect 16545 22615 16579 22649
rect 16945 22615 16979 22649
rect 17345 22615 17379 22649
rect 17745 22615 17779 22649
rect 18145 22615 18179 22649
rect 18545 22615 18579 22649
rect 18945 22615 18979 22649
rect 19345 22615 19379 22649
rect 19745 22615 19779 22649
rect 20145 22615 20179 22649
rect 20545 22615 20579 22649
rect 21191 22615 21225 22649
rect 21391 22615 21425 22649
rect 21591 22615 21625 22649
rect 21791 22615 21825 22649
rect 21991 22615 22025 22649
rect 22191 22615 22225 22649
rect 23151 22615 23185 22649
rect 23551 22615 23585 22649
rect 23951 22615 23985 22649
rect 24351 22615 24385 22649
rect 24751 22615 24785 22649
rect 25151 22615 25185 22649
rect 25551 22615 25585 22649
rect 25951 22615 25985 22649
rect 26351 22615 26385 22649
rect 26751 22615 26785 22649
rect 28443 22615 28477 22649
rect 28643 22615 28677 22649
rect 28843 22615 28877 22649
rect 29043 22615 29077 22649
rect 29243 22615 29277 22649
rect 29443 22615 29477 22649
rect 29643 22615 29677 22649
rect 29843 22615 29877 22649
rect 30043 22615 30077 22649
rect 30243 22615 30277 22649
rect 30443 22615 30477 22649
rect 30643 22615 30677 22649
rect 30843 22615 30877 22649
rect 31043 22615 31077 22649
rect 31243 22615 31277 22649
rect 31443 22615 31477 22649
rect 31643 22615 31677 22649
rect 31843 22615 31877 22649
rect 32043 22615 32077 22649
rect 32243 22615 32277 22649
rect 32443 22615 32477 22649
rect 32643 22615 32677 22649
rect 32843 22615 32877 22649
rect 33043 22615 33077 22649
rect 33243 22615 33277 22649
rect 33443 22615 33477 22649
rect 33643 22615 33677 22649
rect 33843 22615 33877 22649
rect 34043 22615 34077 22649
rect 34243 22615 34277 22649
rect 34443 22615 34477 22649
rect 34643 22615 34677 22649
rect 34843 22615 34877 22649
rect 35043 22615 35077 22649
rect 35243 22615 35277 22649
rect 35443 22615 35477 22649
rect 35643 22615 35677 22649
rect 35843 22615 35877 22649
rect 36043 22615 36077 22649
rect 36243 22615 36277 22649
rect 36443 22615 36477 22649
rect 36643 22615 36677 22649
rect 36843 22615 36877 22649
rect 37043 22615 37077 22649
rect 37243 22615 37277 22649
rect 37443 22615 37477 22649
rect 37643 22615 37677 22649
rect 37843 22615 37877 22649
rect 38043 22615 38077 22649
rect 38243 22615 38277 22649
rect 38443 22615 38477 22649
rect 38643 22615 38677 22649
rect 38843 22615 38877 22649
rect 39929 22615 39963 22649
rect 40129 22615 40163 22649
rect 40329 22615 40363 22649
rect 40529 22615 40563 22649
rect 40729 22615 40763 22649
rect 40929 22615 40963 22649
rect 41129 22615 41163 22649
rect 41329 22615 41363 22649
rect 41529 22615 41563 22649
rect 41729 22615 41763 22649
rect 41929 22615 41963 22649
rect 8309 22457 8343 22491
rect 26433 22457 26467 22491
rect 7727 22347 7761 22381
rect 7727 22279 7761 22309
rect 7727 22275 7761 22279
rect 7727 22211 7761 22237
rect 7727 22203 7761 22211
rect 7727 22143 7761 22165
rect 7727 22131 7761 22143
rect 7727 22075 7761 22093
rect 7727 22059 7761 22075
rect 7727 22007 7761 22021
rect 7727 21987 7761 22007
rect 7727 21939 7761 21949
rect 7727 21915 7761 21939
rect 7727 21871 7761 21877
rect 7727 21843 7761 21871
rect 7727 21803 7761 21805
rect 7727 21771 7761 21803
rect 7727 21701 7761 21733
rect 7727 21699 7761 21701
rect 7727 21633 7761 21661
rect 7727 21627 7761 21633
rect 7727 21565 7761 21589
rect 7727 21555 7761 21565
rect 7727 21497 7761 21517
rect 7727 21483 7761 21497
rect 7727 21429 7761 21445
rect 7727 21411 7761 21429
rect 7727 21361 7761 21373
rect 7727 21339 7761 21361
rect 7727 21293 7761 21301
rect 7727 21267 7761 21293
rect 7727 21225 7761 21229
rect 7727 21195 7761 21225
rect 7727 21123 7761 21157
rect 8185 22347 8219 22381
rect 8185 22279 8219 22309
rect 8185 22275 8219 22279
rect 8185 22211 8219 22237
rect 8185 22203 8219 22211
rect 8185 22143 8219 22165
rect 8185 22131 8219 22143
rect 8185 22075 8219 22093
rect 8185 22059 8219 22075
rect 8185 22007 8219 22021
rect 8185 21987 8219 22007
rect 8185 21939 8219 21949
rect 8185 21915 8219 21939
rect 8185 21871 8219 21877
rect 8185 21843 8219 21871
rect 8185 21803 8219 21805
rect 8185 21771 8219 21803
rect 8185 21701 8219 21733
rect 8185 21699 8219 21701
rect 8185 21633 8219 21661
rect 8185 21627 8219 21633
rect 8185 21565 8219 21589
rect 8185 21555 8219 21565
rect 8185 21497 8219 21517
rect 8185 21483 8219 21497
rect 8185 21429 8219 21445
rect 8185 21411 8219 21429
rect 8185 21361 8219 21373
rect 8185 21339 8219 21361
rect 8185 21293 8219 21301
rect 8185 21267 8219 21293
rect 8185 21225 8219 21229
rect 8185 21195 8219 21225
rect 8185 21123 8219 21157
rect 8643 22347 8677 22381
rect 8643 22279 8677 22309
rect 8643 22275 8677 22279
rect 8643 22211 8677 22237
rect 8643 22203 8677 22211
rect 8643 22143 8677 22165
rect 8643 22131 8677 22143
rect 8643 22075 8677 22093
rect 8643 22059 8677 22075
rect 8643 22007 8677 22021
rect 8643 21987 8677 22007
rect 8643 21939 8677 21949
rect 8643 21915 8677 21939
rect 8643 21871 8677 21877
rect 8643 21843 8677 21871
rect 8643 21803 8677 21805
rect 8643 21771 8677 21803
rect 8643 21701 8677 21733
rect 8643 21699 8677 21701
rect 8643 21633 8677 21661
rect 8643 21627 8677 21633
rect 8643 21565 8677 21589
rect 8643 21555 8677 21565
rect 8643 21497 8677 21517
rect 8643 21483 8677 21497
rect 8643 21429 8677 21445
rect 8643 21411 8677 21429
rect 8643 21361 8677 21373
rect 8643 21339 8677 21361
rect 8643 21293 8677 21301
rect 8643 21267 8677 21293
rect 8643 21225 8677 21229
rect 8643 21195 8677 21225
rect 8643 21123 8677 21157
rect 9101 22347 9135 22381
rect 9101 22279 9135 22309
rect 9101 22275 9135 22279
rect 9101 22211 9135 22237
rect 9101 22203 9135 22211
rect 9101 22143 9135 22165
rect 9101 22131 9135 22143
rect 9101 22075 9135 22093
rect 9101 22059 9135 22075
rect 9101 22007 9135 22021
rect 9101 21987 9135 22007
rect 9101 21939 9135 21949
rect 9101 21915 9135 21939
rect 9101 21871 9135 21877
rect 9101 21843 9135 21871
rect 9101 21803 9135 21805
rect 9101 21771 9135 21803
rect 9101 21701 9135 21733
rect 9101 21699 9135 21701
rect 9101 21633 9135 21661
rect 9101 21627 9135 21633
rect 9101 21565 9135 21589
rect 9101 21555 9135 21565
rect 9101 21497 9135 21517
rect 9101 21483 9135 21497
rect 9101 21429 9135 21445
rect 9101 21411 9135 21429
rect 9101 21361 9135 21373
rect 9101 21339 9135 21361
rect 9101 21293 9135 21301
rect 9101 21267 9135 21293
rect 9101 21225 9135 21229
rect 9101 21195 9135 21225
rect 9101 21123 9135 21157
rect 9559 22347 9593 22381
rect 9559 22279 9593 22309
rect 9559 22275 9593 22279
rect 9559 22211 9593 22237
rect 9559 22203 9593 22211
rect 9559 22143 9593 22165
rect 9559 22131 9593 22143
rect 9559 22075 9593 22093
rect 9559 22059 9593 22075
rect 9559 22007 9593 22021
rect 9559 21987 9593 22007
rect 9559 21939 9593 21949
rect 9559 21915 9593 21939
rect 9559 21871 9593 21877
rect 9559 21843 9593 21871
rect 9559 21803 9593 21805
rect 9559 21771 9593 21803
rect 9559 21701 9593 21733
rect 9559 21699 9593 21701
rect 9559 21633 9593 21661
rect 9559 21627 9593 21633
rect 9559 21565 9593 21589
rect 9559 21555 9593 21565
rect 9559 21497 9593 21517
rect 9559 21483 9593 21497
rect 9559 21429 9593 21445
rect 9559 21411 9593 21429
rect 9559 21361 9593 21373
rect 9559 21339 9593 21361
rect 9559 21293 9593 21301
rect 9559 21267 9593 21293
rect 9559 21225 9593 21229
rect 9559 21195 9593 21225
rect 9559 21123 9593 21157
rect 10017 22347 10051 22381
rect 10017 22279 10051 22309
rect 10017 22275 10051 22279
rect 10017 22211 10051 22237
rect 10017 22203 10051 22211
rect 10017 22143 10051 22165
rect 10017 22131 10051 22143
rect 10017 22075 10051 22093
rect 10017 22059 10051 22075
rect 10017 22007 10051 22021
rect 10017 21987 10051 22007
rect 10017 21939 10051 21949
rect 10017 21915 10051 21939
rect 10017 21871 10051 21877
rect 10017 21843 10051 21871
rect 10017 21803 10051 21805
rect 10017 21771 10051 21803
rect 10017 21701 10051 21733
rect 10017 21699 10051 21701
rect 10017 21633 10051 21661
rect 10017 21627 10051 21633
rect 10017 21565 10051 21589
rect 10017 21555 10051 21565
rect 10017 21497 10051 21517
rect 10017 21483 10051 21497
rect 10017 21429 10051 21445
rect 10017 21411 10051 21429
rect 10017 21361 10051 21373
rect 10017 21339 10051 21361
rect 10017 21293 10051 21301
rect 10017 21267 10051 21293
rect 10017 21225 10051 21229
rect 10017 21195 10051 21225
rect 10017 21123 10051 21157
rect 10475 22347 10509 22381
rect 10475 22279 10509 22309
rect 10475 22275 10509 22279
rect 10475 22211 10509 22237
rect 10475 22203 10509 22211
rect 10475 22143 10509 22165
rect 10475 22131 10509 22143
rect 10475 22075 10509 22093
rect 10475 22059 10509 22075
rect 10475 22007 10509 22021
rect 10475 21987 10509 22007
rect 10475 21939 10509 21949
rect 10475 21915 10509 21939
rect 10475 21871 10509 21877
rect 10475 21843 10509 21871
rect 10475 21803 10509 21805
rect 10475 21771 10509 21803
rect 10475 21701 10509 21733
rect 10475 21699 10509 21701
rect 10475 21633 10509 21661
rect 10475 21627 10509 21633
rect 10475 21565 10509 21589
rect 10475 21555 10509 21565
rect 10475 21497 10509 21517
rect 10475 21483 10509 21497
rect 10475 21429 10509 21445
rect 10475 21411 10509 21429
rect 10475 21361 10509 21373
rect 10475 21339 10509 21361
rect 10475 21293 10509 21301
rect 10475 21267 10509 21293
rect 10475 21225 10509 21229
rect 10475 21195 10509 21225
rect 10475 21123 10509 21157
rect 10933 22347 10967 22381
rect 10933 22279 10967 22309
rect 10933 22275 10967 22279
rect 10933 22211 10967 22237
rect 10933 22203 10967 22211
rect 10933 22143 10967 22165
rect 10933 22131 10967 22143
rect 10933 22075 10967 22093
rect 10933 22059 10967 22075
rect 10933 22007 10967 22021
rect 10933 21987 10967 22007
rect 10933 21939 10967 21949
rect 10933 21915 10967 21939
rect 10933 21871 10967 21877
rect 10933 21843 10967 21871
rect 10933 21803 10967 21805
rect 10933 21771 10967 21803
rect 10933 21701 10967 21733
rect 10933 21699 10967 21701
rect 10933 21633 10967 21661
rect 10933 21627 10967 21633
rect 10933 21565 10967 21589
rect 10933 21555 10967 21565
rect 10933 21497 10967 21517
rect 10933 21483 10967 21497
rect 10933 21429 10967 21445
rect 10933 21411 10967 21429
rect 10933 21361 10967 21373
rect 10933 21339 10967 21361
rect 10933 21293 10967 21301
rect 10933 21267 10967 21293
rect 10933 21225 10967 21229
rect 10933 21195 10967 21225
rect 10933 21123 10967 21157
rect 11391 22347 11425 22381
rect 11391 22279 11425 22309
rect 11391 22275 11425 22279
rect 11391 22211 11425 22237
rect 11391 22203 11425 22211
rect 11391 22143 11425 22165
rect 11391 22131 11425 22143
rect 11391 22075 11425 22093
rect 11391 22059 11425 22075
rect 11391 22007 11425 22021
rect 11391 21987 11425 22007
rect 11391 21939 11425 21949
rect 11391 21915 11425 21939
rect 11391 21871 11425 21877
rect 11391 21843 11425 21871
rect 11391 21803 11425 21805
rect 11391 21771 11425 21803
rect 11391 21701 11425 21733
rect 11391 21699 11425 21701
rect 11391 21633 11425 21661
rect 11391 21627 11425 21633
rect 11391 21565 11425 21589
rect 11391 21555 11425 21565
rect 11391 21497 11425 21517
rect 11391 21483 11425 21497
rect 11391 21429 11425 21445
rect 11391 21411 11425 21429
rect 11391 21361 11425 21373
rect 11391 21339 11425 21361
rect 11391 21293 11425 21301
rect 11391 21267 11425 21293
rect 11391 21225 11425 21229
rect 11391 21195 11425 21225
rect 11391 21123 11425 21157
rect 11849 22347 11883 22381
rect 11849 22279 11883 22309
rect 11849 22275 11883 22279
rect 11849 22211 11883 22237
rect 11849 22203 11883 22211
rect 11849 22143 11883 22165
rect 11849 22131 11883 22143
rect 11849 22075 11883 22093
rect 11849 22059 11883 22075
rect 11849 22007 11883 22021
rect 11849 21987 11883 22007
rect 11849 21939 11883 21949
rect 11849 21915 11883 21939
rect 11849 21871 11883 21877
rect 11849 21843 11883 21871
rect 11849 21803 11883 21805
rect 11849 21771 11883 21803
rect 11849 21701 11883 21733
rect 11849 21699 11883 21701
rect 11849 21633 11883 21661
rect 11849 21627 11883 21633
rect 11849 21565 11883 21589
rect 11849 21555 11883 21565
rect 11849 21497 11883 21517
rect 11849 21483 11883 21497
rect 11849 21429 11883 21445
rect 11849 21411 11883 21429
rect 11849 21361 11883 21373
rect 11849 21339 11883 21361
rect 11849 21293 11883 21301
rect 11849 21267 11883 21293
rect 11849 21225 11883 21229
rect 11849 21195 11883 21225
rect 11849 21123 11883 21157
rect 12307 22347 12341 22381
rect 12307 22279 12341 22309
rect 12307 22275 12341 22279
rect 12307 22211 12341 22237
rect 12307 22203 12341 22211
rect 12307 22143 12341 22165
rect 12307 22131 12341 22143
rect 12307 22075 12341 22093
rect 12307 22059 12341 22075
rect 12307 22007 12341 22021
rect 12307 21987 12341 22007
rect 12307 21939 12341 21949
rect 12307 21915 12341 21939
rect 12307 21871 12341 21877
rect 12307 21843 12341 21871
rect 12307 21803 12341 21805
rect 12307 21771 12341 21803
rect 12307 21701 12341 21733
rect 12307 21699 12341 21701
rect 12307 21633 12341 21661
rect 12307 21627 12341 21633
rect 12307 21565 12341 21589
rect 12307 21555 12341 21565
rect 12307 21497 12341 21517
rect 12307 21483 12341 21497
rect 12307 21429 12341 21445
rect 12307 21411 12341 21429
rect 12307 21361 12341 21373
rect 12307 21339 12341 21361
rect 12307 21293 12341 21301
rect 12307 21267 12341 21293
rect 12307 21225 12341 21229
rect 12307 21195 12341 21225
rect 12307 21123 12341 21157
rect 12765 22347 12799 22381
rect 12765 22279 12799 22309
rect 12765 22275 12799 22279
rect 12765 22211 12799 22237
rect 12765 22203 12799 22211
rect 12765 22143 12799 22165
rect 12765 22131 12799 22143
rect 12765 22075 12799 22093
rect 12765 22059 12799 22075
rect 12765 22007 12799 22021
rect 12765 21987 12799 22007
rect 12765 21939 12799 21949
rect 12765 21915 12799 21939
rect 12765 21871 12799 21877
rect 12765 21843 12799 21871
rect 12765 21803 12799 21805
rect 12765 21771 12799 21803
rect 12765 21701 12799 21733
rect 12765 21699 12799 21701
rect 12765 21633 12799 21661
rect 12765 21627 12799 21633
rect 12765 21565 12799 21589
rect 12765 21555 12799 21565
rect 12765 21497 12799 21517
rect 12765 21483 12799 21497
rect 12765 21429 12799 21445
rect 12765 21411 12799 21429
rect 12765 21361 12799 21373
rect 12765 21339 12799 21361
rect 12765 21293 12799 21301
rect 12765 21267 12799 21293
rect 12765 21225 12799 21229
rect 12765 21195 12799 21225
rect 12765 21123 12799 21157
rect 13223 22347 13257 22381
rect 13223 22279 13257 22309
rect 13223 22275 13257 22279
rect 13223 22211 13257 22237
rect 13223 22203 13257 22211
rect 13223 22143 13257 22165
rect 13223 22131 13257 22143
rect 13223 22075 13257 22093
rect 13223 22059 13257 22075
rect 13223 22007 13257 22021
rect 13223 21987 13257 22007
rect 13223 21939 13257 21949
rect 13223 21915 13257 21939
rect 13223 21871 13257 21877
rect 13223 21843 13257 21871
rect 13223 21803 13257 21805
rect 13223 21771 13257 21803
rect 13223 21701 13257 21733
rect 13223 21699 13257 21701
rect 13223 21633 13257 21661
rect 13223 21627 13257 21633
rect 13223 21565 13257 21589
rect 13223 21555 13257 21565
rect 13223 21497 13257 21517
rect 13223 21483 13257 21497
rect 13223 21429 13257 21445
rect 13223 21411 13257 21429
rect 13223 21361 13257 21373
rect 13223 21339 13257 21361
rect 13223 21293 13257 21301
rect 13223 21267 13257 21293
rect 13223 21225 13257 21229
rect 13223 21195 13257 21225
rect 13223 21123 13257 21157
rect 21404 21946 21426 21952
rect 21426 21946 21438 21952
rect 21504 21946 21516 21952
rect 21516 21946 21538 21952
rect 21604 21946 21606 21952
rect 21606 21946 21638 21952
rect 21404 21918 21438 21946
rect 21504 21918 21538 21946
rect 21604 21918 21638 21946
rect 21704 21918 21738 21952
rect 21804 21918 21838 21952
rect 21904 21946 21932 21952
rect 21932 21946 21938 21952
rect 21904 21918 21938 21946
rect 21404 21818 21438 21852
rect 21504 21818 21538 21852
rect 21604 21818 21638 21852
rect 21704 21818 21738 21852
rect 21804 21818 21838 21852
rect 21904 21818 21938 21852
rect 21404 21718 21438 21752
rect 21504 21718 21538 21752
rect 21604 21718 21638 21752
rect 21704 21718 21738 21752
rect 21804 21718 21838 21752
rect 21904 21718 21938 21752
rect 21404 21620 21438 21652
rect 21504 21620 21538 21652
rect 21604 21620 21638 21652
rect 21404 21618 21426 21620
rect 21426 21618 21438 21620
rect 21504 21618 21516 21620
rect 21516 21618 21538 21620
rect 21604 21618 21606 21620
rect 21606 21618 21638 21620
rect 21704 21618 21738 21652
rect 21804 21618 21838 21652
rect 21904 21620 21938 21652
rect 21904 21618 21932 21620
rect 21932 21618 21938 21620
rect 21404 21530 21438 21552
rect 21504 21530 21538 21552
rect 21604 21530 21638 21552
rect 21404 21518 21426 21530
rect 21426 21518 21438 21530
rect 21504 21518 21516 21530
rect 21516 21518 21538 21530
rect 21604 21518 21606 21530
rect 21606 21518 21638 21530
rect 21704 21518 21738 21552
rect 21804 21518 21838 21552
rect 21904 21530 21938 21552
rect 21904 21518 21932 21530
rect 21932 21518 21938 21530
rect 21404 21440 21438 21452
rect 21504 21440 21538 21452
rect 21604 21440 21638 21452
rect 21404 21418 21426 21440
rect 21426 21418 21438 21440
rect 21504 21418 21516 21440
rect 21516 21418 21538 21440
rect 21604 21418 21606 21440
rect 21606 21418 21638 21440
rect 21704 21418 21738 21452
rect 21804 21418 21838 21452
rect 21904 21440 21938 21452
rect 21904 21418 21932 21440
rect 21932 21418 21938 21440
rect 21189 21233 21223 21267
rect 28306 22282 28340 22316
rect 28396 22301 28430 22316
rect 28486 22301 28520 22316
rect 28576 22301 28610 22316
rect 28666 22301 28700 22316
rect 28756 22301 28790 22316
rect 28846 22301 28880 22316
rect 28936 22301 28970 22316
rect 29026 22301 29060 22316
rect 29116 22301 29150 22316
rect 29206 22301 29240 22316
rect 29296 22301 29330 22316
rect 29386 22301 29420 22316
rect 28396 22282 28416 22301
rect 28416 22282 28430 22301
rect 28486 22282 28506 22301
rect 28506 22282 28520 22301
rect 28576 22282 28596 22301
rect 28596 22282 28610 22301
rect 28666 22282 28686 22301
rect 28686 22282 28700 22301
rect 28756 22282 28776 22301
rect 28776 22282 28790 22301
rect 28846 22282 28866 22301
rect 28866 22282 28880 22301
rect 28936 22282 28956 22301
rect 28956 22282 28970 22301
rect 29026 22282 29046 22301
rect 29046 22282 29060 22301
rect 29116 22282 29136 22301
rect 29136 22282 29150 22301
rect 29206 22282 29226 22301
rect 29226 22282 29240 22301
rect 29296 22282 29316 22301
rect 29316 22282 29330 22301
rect 29386 22282 29406 22301
rect 29406 22282 29420 22301
rect 29476 22282 29510 22316
rect 29646 22282 29680 22316
rect 29736 22301 29770 22316
rect 29826 22301 29860 22316
rect 29916 22301 29950 22316
rect 30006 22301 30040 22316
rect 30096 22301 30130 22316
rect 30186 22301 30220 22316
rect 30276 22301 30310 22316
rect 30366 22301 30400 22316
rect 30456 22301 30490 22316
rect 30546 22301 30580 22316
rect 30636 22301 30670 22316
rect 30726 22301 30760 22316
rect 29736 22282 29756 22301
rect 29756 22282 29770 22301
rect 29826 22282 29846 22301
rect 29846 22282 29860 22301
rect 29916 22282 29936 22301
rect 29936 22282 29950 22301
rect 30006 22282 30026 22301
rect 30026 22282 30040 22301
rect 30096 22282 30116 22301
rect 30116 22282 30130 22301
rect 30186 22282 30206 22301
rect 30206 22282 30220 22301
rect 30276 22282 30296 22301
rect 30296 22282 30310 22301
rect 30366 22282 30386 22301
rect 30386 22282 30400 22301
rect 30456 22282 30476 22301
rect 30476 22282 30490 22301
rect 30546 22282 30566 22301
rect 30566 22282 30580 22301
rect 30636 22282 30656 22301
rect 30656 22282 30670 22301
rect 30726 22282 30746 22301
rect 30746 22282 30760 22301
rect 30816 22282 30850 22316
rect 30986 22282 31020 22316
rect 31076 22301 31110 22316
rect 31166 22301 31200 22316
rect 31256 22301 31290 22316
rect 31346 22301 31380 22316
rect 31436 22301 31470 22316
rect 31526 22301 31560 22316
rect 31616 22301 31650 22316
rect 31706 22301 31740 22316
rect 31796 22301 31830 22316
rect 31886 22301 31920 22316
rect 31976 22301 32010 22316
rect 32066 22301 32100 22316
rect 31076 22282 31096 22301
rect 31096 22282 31110 22301
rect 31166 22282 31186 22301
rect 31186 22282 31200 22301
rect 31256 22282 31276 22301
rect 31276 22282 31290 22301
rect 31346 22282 31366 22301
rect 31366 22282 31380 22301
rect 31436 22282 31456 22301
rect 31456 22282 31470 22301
rect 31526 22282 31546 22301
rect 31546 22282 31560 22301
rect 31616 22282 31636 22301
rect 31636 22282 31650 22301
rect 31706 22282 31726 22301
rect 31726 22282 31740 22301
rect 31796 22282 31816 22301
rect 31816 22282 31830 22301
rect 31886 22282 31906 22301
rect 31906 22282 31920 22301
rect 31976 22282 31996 22301
rect 31996 22282 32010 22301
rect 32066 22282 32086 22301
rect 32086 22282 32100 22301
rect 32156 22282 32190 22316
rect 32326 22282 32360 22316
rect 32416 22301 32450 22316
rect 32506 22301 32540 22316
rect 32596 22301 32630 22316
rect 32686 22301 32720 22316
rect 32776 22301 32810 22316
rect 32866 22301 32900 22316
rect 32956 22301 32990 22316
rect 33046 22301 33080 22316
rect 33136 22301 33170 22316
rect 33226 22301 33260 22316
rect 33316 22301 33350 22316
rect 33406 22301 33440 22316
rect 32416 22282 32436 22301
rect 32436 22282 32450 22301
rect 32506 22282 32526 22301
rect 32526 22282 32540 22301
rect 32596 22282 32616 22301
rect 32616 22282 32630 22301
rect 32686 22282 32706 22301
rect 32706 22282 32720 22301
rect 32776 22282 32796 22301
rect 32796 22282 32810 22301
rect 32866 22282 32886 22301
rect 32886 22282 32900 22301
rect 32956 22282 32976 22301
rect 32976 22282 32990 22301
rect 33046 22282 33066 22301
rect 33066 22282 33080 22301
rect 33136 22282 33156 22301
rect 33156 22282 33170 22301
rect 33226 22282 33246 22301
rect 33246 22282 33260 22301
rect 33316 22282 33336 22301
rect 33336 22282 33350 22301
rect 33406 22282 33426 22301
rect 33426 22282 33440 22301
rect 33496 22282 33530 22316
rect 33666 22282 33700 22316
rect 33756 22301 33790 22316
rect 33846 22301 33880 22316
rect 33936 22301 33970 22316
rect 34026 22301 34060 22316
rect 34116 22301 34150 22316
rect 34206 22301 34240 22316
rect 34296 22301 34330 22316
rect 34386 22301 34420 22316
rect 34476 22301 34510 22316
rect 34566 22301 34600 22316
rect 34656 22301 34690 22316
rect 34746 22301 34780 22316
rect 33756 22282 33776 22301
rect 33776 22282 33790 22301
rect 33846 22282 33866 22301
rect 33866 22282 33880 22301
rect 33936 22282 33956 22301
rect 33956 22282 33970 22301
rect 34026 22282 34046 22301
rect 34046 22282 34060 22301
rect 34116 22282 34136 22301
rect 34136 22282 34150 22301
rect 34206 22282 34226 22301
rect 34226 22282 34240 22301
rect 34296 22282 34316 22301
rect 34316 22282 34330 22301
rect 34386 22282 34406 22301
rect 34406 22282 34420 22301
rect 34476 22282 34496 22301
rect 34496 22282 34510 22301
rect 34566 22282 34586 22301
rect 34586 22282 34600 22301
rect 34656 22282 34676 22301
rect 34676 22282 34690 22301
rect 34746 22282 34766 22301
rect 34766 22282 34780 22301
rect 34836 22282 34870 22316
rect 35006 22282 35040 22316
rect 35096 22301 35130 22316
rect 35186 22301 35220 22316
rect 35276 22301 35310 22316
rect 35366 22301 35400 22316
rect 35456 22301 35490 22316
rect 35546 22301 35580 22316
rect 35636 22301 35670 22316
rect 35726 22301 35760 22316
rect 35816 22301 35850 22316
rect 35906 22301 35940 22316
rect 35996 22301 36030 22316
rect 36086 22301 36120 22316
rect 35096 22282 35116 22301
rect 35116 22282 35130 22301
rect 35186 22282 35206 22301
rect 35206 22282 35220 22301
rect 35276 22282 35296 22301
rect 35296 22282 35310 22301
rect 35366 22282 35386 22301
rect 35386 22282 35400 22301
rect 35456 22282 35476 22301
rect 35476 22282 35490 22301
rect 35546 22282 35566 22301
rect 35566 22282 35580 22301
rect 35636 22282 35656 22301
rect 35656 22282 35670 22301
rect 35726 22282 35746 22301
rect 35746 22282 35760 22301
rect 35816 22282 35836 22301
rect 35836 22282 35850 22301
rect 35906 22282 35926 22301
rect 35926 22282 35940 22301
rect 35996 22282 36016 22301
rect 36016 22282 36030 22301
rect 36086 22282 36106 22301
rect 36106 22282 36120 22301
rect 36176 22282 36210 22316
rect 36346 22282 36380 22316
rect 36436 22301 36470 22316
rect 36526 22301 36560 22316
rect 36616 22301 36650 22316
rect 36706 22301 36740 22316
rect 36796 22301 36830 22316
rect 36886 22301 36920 22316
rect 36976 22301 37010 22316
rect 37066 22301 37100 22316
rect 37156 22301 37190 22316
rect 37246 22301 37280 22316
rect 37336 22301 37370 22316
rect 37426 22301 37460 22316
rect 36436 22282 36456 22301
rect 36456 22282 36470 22301
rect 36526 22282 36546 22301
rect 36546 22282 36560 22301
rect 36616 22282 36636 22301
rect 36636 22282 36650 22301
rect 36706 22282 36726 22301
rect 36726 22282 36740 22301
rect 36796 22282 36816 22301
rect 36816 22282 36830 22301
rect 36886 22282 36906 22301
rect 36906 22282 36920 22301
rect 36976 22282 36996 22301
rect 36996 22282 37010 22301
rect 37066 22282 37086 22301
rect 37086 22282 37100 22301
rect 37156 22282 37176 22301
rect 37176 22282 37190 22301
rect 37246 22282 37266 22301
rect 37266 22282 37280 22301
rect 37336 22282 37356 22301
rect 37356 22282 37370 22301
rect 37426 22282 37446 22301
rect 37446 22282 37460 22301
rect 37516 22282 37550 22316
rect 37686 22282 37720 22316
rect 37776 22301 37810 22316
rect 37866 22301 37900 22316
rect 37956 22301 37990 22316
rect 38046 22301 38080 22316
rect 38136 22301 38170 22316
rect 38226 22301 38260 22316
rect 38316 22301 38350 22316
rect 38406 22301 38440 22316
rect 38496 22301 38530 22316
rect 38586 22301 38620 22316
rect 38676 22301 38710 22316
rect 38766 22301 38800 22316
rect 37776 22282 37796 22301
rect 37796 22282 37810 22301
rect 37866 22282 37886 22301
rect 37886 22282 37900 22301
rect 37956 22282 37976 22301
rect 37976 22282 37990 22301
rect 38046 22282 38066 22301
rect 38066 22282 38080 22301
rect 38136 22282 38156 22301
rect 38156 22282 38170 22301
rect 38226 22282 38246 22301
rect 38246 22282 38260 22301
rect 38316 22282 38336 22301
rect 38336 22282 38350 22301
rect 38406 22282 38426 22301
rect 38426 22282 38440 22301
rect 38496 22282 38516 22301
rect 38516 22282 38530 22301
rect 38586 22282 38606 22301
rect 38606 22282 38620 22301
rect 38676 22282 38696 22301
rect 38696 22282 38710 22301
rect 38766 22282 38786 22301
rect 38786 22282 38800 22301
rect 38856 22282 38890 22316
rect 22980 22109 23014 22129
rect 22980 22095 23014 22109
rect 22980 22041 23014 22057
rect 22980 22023 23014 22041
rect 22980 21973 23014 21985
rect 22980 21951 23014 21973
rect 22980 21905 23014 21913
rect 22980 21879 23014 21905
rect 22980 21837 23014 21841
rect 22980 21807 23014 21837
rect 22980 21735 23014 21769
rect 22980 21667 23014 21697
rect 22980 21663 23014 21667
rect 22980 21599 23014 21625
rect 22980 21591 23014 21599
rect 22980 21531 23014 21553
rect 22980 21519 23014 21531
rect 22980 21463 23014 21481
rect 22980 21447 23014 21463
rect 22980 21395 23014 21409
rect 22980 21375 23014 21395
rect 23438 22109 23472 22129
rect 23438 22095 23472 22109
rect 23438 22041 23472 22057
rect 23438 22023 23472 22041
rect 23438 21973 23472 21985
rect 23438 21951 23472 21973
rect 23438 21905 23472 21913
rect 23438 21879 23472 21905
rect 23438 21837 23472 21841
rect 23438 21807 23472 21837
rect 23438 21735 23472 21769
rect 23438 21667 23472 21697
rect 23438 21663 23472 21667
rect 23438 21599 23472 21625
rect 23438 21591 23472 21599
rect 23438 21531 23472 21553
rect 23438 21519 23472 21531
rect 23438 21463 23472 21481
rect 23438 21447 23472 21463
rect 23438 21395 23472 21409
rect 23896 22109 23930 22129
rect 23896 22095 23930 22109
rect 23896 22041 23930 22057
rect 23896 22023 23930 22041
rect 23896 21973 23930 21985
rect 23896 21951 23930 21973
rect 23896 21905 23930 21913
rect 23896 21879 23930 21905
rect 23896 21837 23930 21841
rect 23896 21807 23930 21837
rect 23896 21735 23930 21769
rect 23896 21667 23930 21697
rect 23896 21663 23930 21667
rect 23896 21599 23930 21625
rect 23896 21591 23930 21599
rect 23896 21531 23930 21553
rect 23896 21519 23930 21531
rect 23896 21463 23930 21481
rect 23896 21447 23930 21463
rect 23438 21375 23472 21395
rect 23896 21395 23930 21409
rect 23896 21375 23930 21395
rect 24354 22109 24388 22129
rect 24354 22095 24388 22109
rect 24354 22041 24388 22057
rect 24354 22023 24388 22041
rect 24354 21973 24388 21985
rect 24354 21951 24388 21973
rect 24354 21905 24388 21913
rect 24354 21879 24388 21905
rect 24354 21837 24388 21841
rect 24354 21807 24388 21837
rect 24354 21735 24388 21769
rect 24354 21667 24388 21697
rect 24354 21663 24388 21667
rect 24354 21599 24388 21625
rect 24354 21591 24388 21599
rect 24354 21531 24388 21553
rect 24354 21519 24388 21531
rect 24354 21463 24388 21481
rect 24354 21447 24388 21463
rect 24354 21395 24388 21409
rect 24812 22109 24846 22129
rect 24812 22095 24846 22109
rect 24812 22041 24846 22057
rect 24812 22023 24846 22041
rect 24812 21973 24846 21985
rect 24812 21951 24846 21973
rect 24812 21905 24846 21913
rect 24812 21879 24846 21905
rect 24812 21837 24846 21841
rect 24812 21807 24846 21837
rect 24812 21735 24846 21769
rect 24812 21667 24846 21697
rect 24812 21663 24846 21667
rect 24812 21599 24846 21625
rect 24812 21591 24846 21599
rect 24812 21531 24846 21553
rect 24812 21519 24846 21531
rect 24812 21463 24846 21481
rect 24812 21447 24846 21463
rect 24354 21375 24388 21395
rect 24812 21395 24846 21409
rect 24812 21375 24846 21395
rect 25270 22109 25304 22129
rect 25270 22095 25304 22109
rect 25270 22041 25304 22057
rect 25270 22023 25304 22041
rect 25270 21973 25304 21985
rect 25270 21951 25304 21973
rect 25270 21905 25304 21913
rect 25270 21879 25304 21905
rect 25270 21837 25304 21841
rect 25270 21807 25304 21837
rect 25270 21735 25304 21769
rect 25270 21667 25304 21697
rect 25270 21663 25304 21667
rect 25270 21599 25304 21625
rect 25270 21591 25304 21599
rect 25270 21531 25304 21553
rect 25270 21519 25304 21531
rect 25270 21463 25304 21481
rect 25270 21447 25304 21463
rect 25270 21395 25304 21409
rect 25728 22109 25762 22129
rect 25728 22095 25762 22109
rect 25728 22041 25762 22057
rect 25728 22023 25762 22041
rect 25728 21973 25762 21985
rect 25728 21951 25762 21973
rect 25728 21905 25762 21913
rect 25728 21879 25762 21905
rect 25728 21837 25762 21841
rect 25728 21807 25762 21837
rect 25728 21735 25762 21769
rect 25728 21667 25762 21697
rect 25728 21663 25762 21667
rect 25728 21599 25762 21625
rect 25728 21591 25762 21599
rect 25728 21531 25762 21553
rect 25728 21519 25762 21531
rect 25728 21463 25762 21481
rect 25728 21447 25762 21463
rect 25270 21375 25304 21395
rect 25728 21395 25762 21409
rect 25728 21375 25762 21395
rect 26186 22109 26220 22129
rect 26186 22095 26220 22109
rect 26186 22041 26220 22057
rect 26186 22023 26220 22041
rect 26186 21973 26220 21985
rect 26186 21951 26220 21973
rect 26186 21905 26220 21913
rect 26186 21879 26220 21905
rect 26186 21837 26220 21841
rect 26186 21807 26220 21837
rect 26186 21735 26220 21769
rect 26186 21667 26220 21697
rect 26186 21663 26220 21667
rect 26186 21599 26220 21625
rect 26186 21591 26220 21599
rect 26186 21531 26220 21553
rect 26186 21519 26220 21531
rect 26186 21463 26220 21481
rect 26186 21447 26220 21463
rect 26186 21395 26220 21409
rect 26644 22109 26678 22129
rect 26644 22095 26678 22109
rect 26644 22041 26678 22057
rect 26644 22023 26678 22041
rect 26644 21973 26678 21985
rect 26644 21951 26678 21973
rect 26644 21905 26678 21913
rect 26644 21879 26678 21905
rect 26644 21837 26678 21841
rect 26644 21807 26678 21837
rect 26644 21735 26678 21769
rect 26644 21667 26678 21697
rect 26644 21663 26678 21667
rect 26644 21599 26678 21625
rect 26644 21591 26678 21599
rect 26644 21531 26678 21553
rect 26644 21519 26678 21531
rect 26644 21463 26678 21481
rect 26644 21447 26678 21463
rect 26186 21375 26220 21395
rect 26644 21395 26678 21409
rect 26644 21375 26678 21395
rect 27102 22109 27136 22129
rect 27102 22095 27136 22109
rect 27102 22041 27136 22057
rect 27102 22023 27136 22041
rect 27102 21973 27136 21985
rect 27102 21951 27136 21973
rect 27102 21905 27136 21913
rect 27102 21879 27136 21905
rect 27102 21837 27136 21841
rect 27102 21807 27136 21837
rect 27102 21735 27136 21769
rect 27102 21667 27136 21697
rect 27102 21663 27136 21667
rect 27102 21599 27136 21625
rect 27102 21591 27136 21599
rect 27102 21531 27136 21553
rect 27102 21519 27136 21531
rect 27102 21463 27136 21481
rect 27102 21447 27136 21463
rect 27102 21395 27136 21409
rect 27102 21375 27136 21395
rect 26525 21233 26559 21267
rect 28470 22122 28504 22156
rect 28560 22154 28594 22156
rect 28650 22154 28684 22156
rect 28740 22154 28774 22156
rect 28830 22154 28864 22156
rect 28920 22154 28954 22156
rect 29010 22154 29044 22156
rect 29100 22154 29134 22156
rect 29190 22154 29224 22156
rect 29280 22154 29314 22156
rect 28560 22122 28580 22154
rect 28580 22122 28594 22154
rect 28650 22122 28670 22154
rect 28670 22122 28684 22154
rect 28740 22122 28760 22154
rect 28760 22122 28774 22154
rect 28830 22122 28850 22154
rect 28850 22122 28864 22154
rect 28920 22122 28940 22154
rect 28940 22122 28954 22154
rect 29010 22122 29030 22154
rect 29030 22122 29044 22154
rect 29100 22122 29120 22154
rect 29120 22122 29134 22154
rect 29190 22122 29210 22154
rect 29210 22122 29224 22154
rect 29280 22122 29300 22154
rect 29300 22122 29314 22154
rect 29370 22122 29404 22156
rect 28656 21946 28678 21952
rect 28678 21946 28690 21952
rect 28756 21946 28768 21952
rect 28768 21946 28790 21952
rect 28856 21946 28858 21952
rect 28858 21946 28890 21952
rect 28656 21918 28690 21946
rect 28756 21918 28790 21946
rect 28856 21918 28890 21946
rect 28956 21918 28990 21952
rect 29056 21918 29090 21952
rect 29156 21946 29184 21952
rect 29184 21946 29190 21952
rect 29156 21918 29190 21946
rect 28656 21818 28690 21852
rect 28756 21818 28790 21852
rect 28856 21818 28890 21852
rect 28956 21818 28990 21852
rect 29056 21818 29090 21852
rect 29156 21818 29190 21852
rect 28656 21718 28690 21752
rect 28756 21718 28790 21752
rect 28856 21718 28890 21752
rect 28956 21718 28990 21752
rect 29056 21718 29090 21752
rect 29156 21718 29190 21752
rect 28656 21620 28690 21652
rect 28756 21620 28790 21652
rect 28856 21620 28890 21652
rect 28656 21618 28678 21620
rect 28678 21618 28690 21620
rect 28756 21618 28768 21620
rect 28768 21618 28790 21620
rect 28856 21618 28858 21620
rect 28858 21618 28890 21620
rect 28956 21618 28990 21652
rect 29056 21618 29090 21652
rect 29156 21620 29190 21652
rect 29156 21618 29184 21620
rect 29184 21618 29190 21620
rect 28656 21530 28690 21552
rect 28756 21530 28790 21552
rect 28856 21530 28890 21552
rect 28656 21518 28678 21530
rect 28678 21518 28690 21530
rect 28756 21518 28768 21530
rect 28768 21518 28790 21530
rect 28856 21518 28858 21530
rect 28858 21518 28890 21530
rect 28956 21518 28990 21552
rect 29056 21518 29090 21552
rect 29156 21530 29190 21552
rect 29156 21518 29184 21530
rect 29184 21518 29190 21530
rect 28656 21440 28690 21452
rect 28756 21440 28790 21452
rect 28856 21440 28890 21452
rect 28656 21418 28678 21440
rect 28678 21418 28690 21440
rect 28756 21418 28768 21440
rect 28768 21418 28790 21440
rect 28856 21418 28858 21440
rect 28858 21418 28890 21440
rect 28956 21418 28990 21452
rect 29056 21418 29090 21452
rect 29156 21440 29190 21452
rect 29156 21418 29184 21440
rect 29184 21418 29190 21440
rect 29810 22122 29844 22156
rect 29900 22154 29934 22156
rect 29990 22154 30024 22156
rect 30080 22154 30114 22156
rect 30170 22154 30204 22156
rect 30260 22154 30294 22156
rect 30350 22154 30384 22156
rect 30440 22154 30474 22156
rect 30530 22154 30564 22156
rect 30620 22154 30654 22156
rect 29900 22122 29920 22154
rect 29920 22122 29934 22154
rect 29990 22122 30010 22154
rect 30010 22122 30024 22154
rect 30080 22122 30100 22154
rect 30100 22122 30114 22154
rect 30170 22122 30190 22154
rect 30190 22122 30204 22154
rect 30260 22122 30280 22154
rect 30280 22122 30294 22154
rect 30350 22122 30370 22154
rect 30370 22122 30384 22154
rect 30440 22122 30460 22154
rect 30460 22122 30474 22154
rect 30530 22122 30550 22154
rect 30550 22122 30564 22154
rect 30620 22122 30640 22154
rect 30640 22122 30654 22154
rect 30710 22122 30744 22156
rect 29996 21946 30018 21952
rect 30018 21946 30030 21952
rect 30096 21946 30108 21952
rect 30108 21946 30130 21952
rect 30196 21946 30198 21952
rect 30198 21946 30230 21952
rect 29996 21918 30030 21946
rect 30096 21918 30130 21946
rect 30196 21918 30230 21946
rect 30296 21918 30330 21952
rect 30396 21918 30430 21952
rect 30496 21946 30524 21952
rect 30524 21946 30530 21952
rect 30496 21918 30530 21946
rect 29996 21818 30030 21852
rect 30096 21818 30130 21852
rect 30196 21818 30230 21852
rect 30296 21818 30330 21852
rect 30396 21818 30430 21852
rect 30496 21818 30530 21852
rect 29996 21718 30030 21752
rect 30096 21718 30130 21752
rect 30196 21718 30230 21752
rect 30296 21718 30330 21752
rect 30396 21718 30430 21752
rect 30496 21718 30530 21752
rect 29996 21620 30030 21652
rect 30096 21620 30130 21652
rect 30196 21620 30230 21652
rect 29996 21618 30018 21620
rect 30018 21618 30030 21620
rect 30096 21618 30108 21620
rect 30108 21618 30130 21620
rect 30196 21618 30198 21620
rect 30198 21618 30230 21620
rect 30296 21618 30330 21652
rect 30396 21618 30430 21652
rect 30496 21620 30530 21652
rect 30496 21618 30524 21620
rect 30524 21618 30530 21620
rect 29996 21530 30030 21552
rect 30096 21530 30130 21552
rect 30196 21530 30230 21552
rect 29996 21518 30018 21530
rect 30018 21518 30030 21530
rect 30096 21518 30108 21530
rect 30108 21518 30130 21530
rect 30196 21518 30198 21530
rect 30198 21518 30230 21530
rect 30296 21518 30330 21552
rect 30396 21518 30430 21552
rect 30496 21530 30530 21552
rect 30496 21518 30524 21530
rect 30524 21518 30530 21530
rect 29996 21440 30030 21452
rect 30096 21440 30130 21452
rect 30196 21440 30230 21452
rect 29996 21418 30018 21440
rect 30018 21418 30030 21440
rect 30096 21418 30108 21440
rect 30108 21418 30130 21440
rect 30196 21418 30198 21440
rect 30198 21418 30230 21440
rect 30296 21418 30330 21452
rect 30396 21418 30430 21452
rect 30496 21440 30530 21452
rect 30496 21418 30524 21440
rect 30524 21418 30530 21440
rect 31150 22122 31184 22156
rect 31240 22154 31274 22156
rect 31330 22154 31364 22156
rect 31420 22154 31454 22156
rect 31510 22154 31544 22156
rect 31600 22154 31634 22156
rect 31690 22154 31724 22156
rect 31780 22154 31814 22156
rect 31870 22154 31904 22156
rect 31960 22154 31994 22156
rect 31240 22122 31260 22154
rect 31260 22122 31274 22154
rect 31330 22122 31350 22154
rect 31350 22122 31364 22154
rect 31420 22122 31440 22154
rect 31440 22122 31454 22154
rect 31510 22122 31530 22154
rect 31530 22122 31544 22154
rect 31600 22122 31620 22154
rect 31620 22122 31634 22154
rect 31690 22122 31710 22154
rect 31710 22122 31724 22154
rect 31780 22122 31800 22154
rect 31800 22122 31814 22154
rect 31870 22122 31890 22154
rect 31890 22122 31904 22154
rect 31960 22122 31980 22154
rect 31980 22122 31994 22154
rect 32050 22122 32084 22156
rect 31336 21946 31358 21952
rect 31358 21946 31370 21952
rect 31436 21946 31448 21952
rect 31448 21946 31470 21952
rect 31536 21946 31538 21952
rect 31538 21946 31570 21952
rect 31336 21918 31370 21946
rect 31436 21918 31470 21946
rect 31536 21918 31570 21946
rect 31636 21918 31670 21952
rect 31736 21918 31770 21952
rect 31836 21946 31864 21952
rect 31864 21946 31870 21952
rect 31836 21918 31870 21946
rect 31336 21818 31370 21852
rect 31436 21818 31470 21852
rect 31536 21818 31570 21852
rect 31636 21818 31670 21852
rect 31736 21818 31770 21852
rect 31836 21818 31870 21852
rect 31336 21718 31370 21752
rect 31436 21718 31470 21752
rect 31536 21718 31570 21752
rect 31636 21718 31670 21752
rect 31736 21718 31770 21752
rect 31836 21718 31870 21752
rect 31336 21620 31370 21652
rect 31436 21620 31470 21652
rect 31536 21620 31570 21652
rect 31336 21618 31358 21620
rect 31358 21618 31370 21620
rect 31436 21618 31448 21620
rect 31448 21618 31470 21620
rect 31536 21618 31538 21620
rect 31538 21618 31570 21620
rect 31636 21618 31670 21652
rect 31736 21618 31770 21652
rect 31836 21620 31870 21652
rect 31836 21618 31864 21620
rect 31864 21618 31870 21620
rect 31336 21530 31370 21552
rect 31436 21530 31470 21552
rect 31536 21530 31570 21552
rect 31336 21518 31358 21530
rect 31358 21518 31370 21530
rect 31436 21518 31448 21530
rect 31448 21518 31470 21530
rect 31536 21518 31538 21530
rect 31538 21518 31570 21530
rect 31636 21518 31670 21552
rect 31736 21518 31770 21552
rect 31836 21530 31870 21552
rect 31836 21518 31864 21530
rect 31864 21518 31870 21530
rect 31336 21440 31370 21452
rect 31436 21440 31470 21452
rect 31536 21440 31570 21452
rect 31336 21418 31358 21440
rect 31358 21418 31370 21440
rect 31436 21418 31448 21440
rect 31448 21418 31470 21440
rect 31536 21418 31538 21440
rect 31538 21418 31570 21440
rect 31636 21418 31670 21452
rect 31736 21418 31770 21452
rect 31836 21440 31870 21452
rect 31836 21418 31864 21440
rect 31864 21418 31870 21440
rect 32490 22122 32524 22156
rect 32580 22154 32614 22156
rect 32670 22154 32704 22156
rect 32760 22154 32794 22156
rect 32850 22154 32884 22156
rect 32940 22154 32974 22156
rect 33030 22154 33064 22156
rect 33120 22154 33154 22156
rect 33210 22154 33244 22156
rect 33300 22154 33334 22156
rect 32580 22122 32600 22154
rect 32600 22122 32614 22154
rect 32670 22122 32690 22154
rect 32690 22122 32704 22154
rect 32760 22122 32780 22154
rect 32780 22122 32794 22154
rect 32850 22122 32870 22154
rect 32870 22122 32884 22154
rect 32940 22122 32960 22154
rect 32960 22122 32974 22154
rect 33030 22122 33050 22154
rect 33050 22122 33064 22154
rect 33120 22122 33140 22154
rect 33140 22122 33154 22154
rect 33210 22122 33230 22154
rect 33230 22122 33244 22154
rect 33300 22122 33320 22154
rect 33320 22122 33334 22154
rect 33390 22122 33424 22156
rect 32676 21946 32698 21952
rect 32698 21946 32710 21952
rect 32776 21946 32788 21952
rect 32788 21946 32810 21952
rect 32876 21946 32878 21952
rect 32878 21946 32910 21952
rect 32676 21918 32710 21946
rect 32776 21918 32810 21946
rect 32876 21918 32910 21946
rect 32976 21918 33010 21952
rect 33076 21918 33110 21952
rect 33176 21946 33204 21952
rect 33204 21946 33210 21952
rect 33176 21918 33210 21946
rect 32676 21818 32710 21852
rect 32776 21818 32810 21852
rect 32876 21818 32910 21852
rect 32976 21818 33010 21852
rect 33076 21818 33110 21852
rect 33176 21818 33210 21852
rect 32676 21718 32710 21752
rect 32776 21718 32810 21752
rect 32876 21718 32910 21752
rect 32976 21718 33010 21752
rect 33076 21718 33110 21752
rect 33176 21718 33210 21752
rect 32676 21620 32710 21652
rect 32776 21620 32810 21652
rect 32876 21620 32910 21652
rect 32676 21618 32698 21620
rect 32698 21618 32710 21620
rect 32776 21618 32788 21620
rect 32788 21618 32810 21620
rect 32876 21618 32878 21620
rect 32878 21618 32910 21620
rect 32976 21618 33010 21652
rect 33076 21618 33110 21652
rect 33176 21620 33210 21652
rect 33176 21618 33204 21620
rect 33204 21618 33210 21620
rect 32676 21530 32710 21552
rect 32776 21530 32810 21552
rect 32876 21530 32910 21552
rect 32676 21518 32698 21530
rect 32698 21518 32710 21530
rect 32776 21518 32788 21530
rect 32788 21518 32810 21530
rect 32876 21518 32878 21530
rect 32878 21518 32910 21530
rect 32976 21518 33010 21552
rect 33076 21518 33110 21552
rect 33176 21530 33210 21552
rect 33176 21518 33204 21530
rect 33204 21518 33210 21530
rect 32676 21440 32710 21452
rect 32776 21440 32810 21452
rect 32876 21440 32910 21452
rect 32676 21418 32698 21440
rect 32698 21418 32710 21440
rect 32776 21418 32788 21440
rect 32788 21418 32810 21440
rect 32876 21418 32878 21440
rect 32878 21418 32910 21440
rect 32976 21418 33010 21452
rect 33076 21418 33110 21452
rect 33176 21440 33210 21452
rect 33176 21418 33204 21440
rect 33204 21418 33210 21440
rect 33830 22122 33864 22156
rect 33920 22154 33954 22156
rect 34010 22154 34044 22156
rect 34100 22154 34134 22156
rect 34190 22154 34224 22156
rect 34280 22154 34314 22156
rect 34370 22154 34404 22156
rect 34460 22154 34494 22156
rect 34550 22154 34584 22156
rect 34640 22154 34674 22156
rect 33920 22122 33940 22154
rect 33940 22122 33954 22154
rect 34010 22122 34030 22154
rect 34030 22122 34044 22154
rect 34100 22122 34120 22154
rect 34120 22122 34134 22154
rect 34190 22122 34210 22154
rect 34210 22122 34224 22154
rect 34280 22122 34300 22154
rect 34300 22122 34314 22154
rect 34370 22122 34390 22154
rect 34390 22122 34404 22154
rect 34460 22122 34480 22154
rect 34480 22122 34494 22154
rect 34550 22122 34570 22154
rect 34570 22122 34584 22154
rect 34640 22122 34660 22154
rect 34660 22122 34674 22154
rect 34730 22122 34764 22156
rect 34016 21946 34038 21952
rect 34038 21946 34050 21952
rect 34116 21946 34128 21952
rect 34128 21946 34150 21952
rect 34216 21946 34218 21952
rect 34218 21946 34250 21952
rect 34016 21918 34050 21946
rect 34116 21918 34150 21946
rect 34216 21918 34250 21946
rect 34316 21918 34350 21952
rect 34416 21918 34450 21952
rect 34516 21946 34544 21952
rect 34544 21946 34550 21952
rect 34516 21918 34550 21946
rect 34016 21818 34050 21852
rect 34116 21818 34150 21852
rect 34216 21818 34250 21852
rect 34316 21818 34350 21852
rect 34416 21818 34450 21852
rect 34516 21818 34550 21852
rect 34016 21718 34050 21752
rect 34116 21718 34150 21752
rect 34216 21718 34250 21752
rect 34316 21718 34350 21752
rect 34416 21718 34450 21752
rect 34516 21718 34550 21752
rect 34016 21620 34050 21652
rect 34116 21620 34150 21652
rect 34216 21620 34250 21652
rect 34016 21618 34038 21620
rect 34038 21618 34050 21620
rect 34116 21618 34128 21620
rect 34128 21618 34150 21620
rect 34216 21618 34218 21620
rect 34218 21618 34250 21620
rect 34316 21618 34350 21652
rect 34416 21618 34450 21652
rect 34516 21620 34550 21652
rect 34516 21618 34544 21620
rect 34544 21618 34550 21620
rect 34016 21530 34050 21552
rect 34116 21530 34150 21552
rect 34216 21530 34250 21552
rect 34016 21518 34038 21530
rect 34038 21518 34050 21530
rect 34116 21518 34128 21530
rect 34128 21518 34150 21530
rect 34216 21518 34218 21530
rect 34218 21518 34250 21530
rect 34316 21518 34350 21552
rect 34416 21518 34450 21552
rect 34516 21530 34550 21552
rect 34516 21518 34544 21530
rect 34544 21518 34550 21530
rect 34016 21440 34050 21452
rect 34116 21440 34150 21452
rect 34216 21440 34250 21452
rect 34016 21418 34038 21440
rect 34038 21418 34050 21440
rect 34116 21418 34128 21440
rect 34128 21418 34150 21440
rect 34216 21418 34218 21440
rect 34218 21418 34250 21440
rect 34316 21418 34350 21452
rect 34416 21418 34450 21452
rect 34516 21440 34550 21452
rect 34516 21418 34544 21440
rect 34544 21418 34550 21440
rect 35170 22122 35204 22156
rect 35260 22154 35294 22156
rect 35350 22154 35384 22156
rect 35440 22154 35474 22156
rect 35530 22154 35564 22156
rect 35620 22154 35654 22156
rect 35710 22154 35744 22156
rect 35800 22154 35834 22156
rect 35890 22154 35924 22156
rect 35980 22154 36014 22156
rect 35260 22122 35280 22154
rect 35280 22122 35294 22154
rect 35350 22122 35370 22154
rect 35370 22122 35384 22154
rect 35440 22122 35460 22154
rect 35460 22122 35474 22154
rect 35530 22122 35550 22154
rect 35550 22122 35564 22154
rect 35620 22122 35640 22154
rect 35640 22122 35654 22154
rect 35710 22122 35730 22154
rect 35730 22122 35744 22154
rect 35800 22122 35820 22154
rect 35820 22122 35834 22154
rect 35890 22122 35910 22154
rect 35910 22122 35924 22154
rect 35980 22122 36000 22154
rect 36000 22122 36014 22154
rect 36070 22122 36104 22156
rect 35356 21946 35378 21952
rect 35378 21946 35390 21952
rect 35456 21946 35468 21952
rect 35468 21946 35490 21952
rect 35556 21946 35558 21952
rect 35558 21946 35590 21952
rect 35356 21918 35390 21946
rect 35456 21918 35490 21946
rect 35556 21918 35590 21946
rect 35656 21918 35690 21952
rect 35756 21918 35790 21952
rect 35856 21946 35884 21952
rect 35884 21946 35890 21952
rect 35856 21918 35890 21946
rect 35356 21818 35390 21852
rect 35456 21818 35490 21852
rect 35556 21818 35590 21852
rect 35656 21818 35690 21852
rect 35756 21818 35790 21852
rect 35856 21818 35890 21852
rect 35356 21718 35390 21752
rect 35456 21718 35490 21752
rect 35556 21718 35590 21752
rect 35656 21718 35690 21752
rect 35756 21718 35790 21752
rect 35856 21718 35890 21752
rect 35356 21620 35390 21652
rect 35456 21620 35490 21652
rect 35556 21620 35590 21652
rect 35356 21618 35378 21620
rect 35378 21618 35390 21620
rect 35456 21618 35468 21620
rect 35468 21618 35490 21620
rect 35556 21618 35558 21620
rect 35558 21618 35590 21620
rect 35656 21618 35690 21652
rect 35756 21618 35790 21652
rect 35856 21620 35890 21652
rect 35856 21618 35884 21620
rect 35884 21618 35890 21620
rect 35356 21530 35390 21552
rect 35456 21530 35490 21552
rect 35556 21530 35590 21552
rect 35356 21518 35378 21530
rect 35378 21518 35390 21530
rect 35456 21518 35468 21530
rect 35468 21518 35490 21530
rect 35556 21518 35558 21530
rect 35558 21518 35590 21530
rect 35656 21518 35690 21552
rect 35756 21518 35790 21552
rect 35856 21530 35890 21552
rect 35856 21518 35884 21530
rect 35884 21518 35890 21530
rect 35356 21440 35390 21452
rect 35456 21440 35490 21452
rect 35556 21440 35590 21452
rect 35356 21418 35378 21440
rect 35378 21418 35390 21440
rect 35456 21418 35468 21440
rect 35468 21418 35490 21440
rect 35556 21418 35558 21440
rect 35558 21418 35590 21440
rect 35656 21418 35690 21452
rect 35756 21418 35790 21452
rect 35856 21440 35890 21452
rect 35856 21418 35884 21440
rect 35884 21418 35890 21440
rect 36510 22122 36544 22156
rect 36600 22154 36634 22156
rect 36690 22154 36724 22156
rect 36780 22154 36814 22156
rect 36870 22154 36904 22156
rect 36960 22154 36994 22156
rect 37050 22154 37084 22156
rect 37140 22154 37174 22156
rect 37230 22154 37264 22156
rect 37320 22154 37354 22156
rect 36600 22122 36620 22154
rect 36620 22122 36634 22154
rect 36690 22122 36710 22154
rect 36710 22122 36724 22154
rect 36780 22122 36800 22154
rect 36800 22122 36814 22154
rect 36870 22122 36890 22154
rect 36890 22122 36904 22154
rect 36960 22122 36980 22154
rect 36980 22122 36994 22154
rect 37050 22122 37070 22154
rect 37070 22122 37084 22154
rect 37140 22122 37160 22154
rect 37160 22122 37174 22154
rect 37230 22122 37250 22154
rect 37250 22122 37264 22154
rect 37320 22122 37340 22154
rect 37340 22122 37354 22154
rect 37410 22122 37444 22156
rect 36696 21946 36718 21952
rect 36718 21946 36730 21952
rect 36796 21946 36808 21952
rect 36808 21946 36830 21952
rect 36896 21946 36898 21952
rect 36898 21946 36930 21952
rect 36696 21918 36730 21946
rect 36796 21918 36830 21946
rect 36896 21918 36930 21946
rect 36996 21918 37030 21952
rect 37096 21918 37130 21952
rect 37196 21946 37224 21952
rect 37224 21946 37230 21952
rect 37196 21918 37230 21946
rect 36696 21818 36730 21852
rect 36796 21818 36830 21852
rect 36896 21818 36930 21852
rect 36996 21818 37030 21852
rect 37096 21818 37130 21852
rect 37196 21818 37230 21852
rect 36696 21718 36730 21752
rect 36796 21718 36830 21752
rect 36896 21718 36930 21752
rect 36996 21718 37030 21752
rect 37096 21718 37130 21752
rect 37196 21718 37230 21752
rect 36696 21620 36730 21652
rect 36796 21620 36830 21652
rect 36896 21620 36930 21652
rect 36696 21618 36718 21620
rect 36718 21618 36730 21620
rect 36796 21618 36808 21620
rect 36808 21618 36830 21620
rect 36896 21618 36898 21620
rect 36898 21618 36930 21620
rect 36996 21618 37030 21652
rect 37096 21618 37130 21652
rect 37196 21620 37230 21652
rect 37196 21618 37224 21620
rect 37224 21618 37230 21620
rect 36696 21530 36730 21552
rect 36796 21530 36830 21552
rect 36896 21530 36930 21552
rect 36696 21518 36718 21530
rect 36718 21518 36730 21530
rect 36796 21518 36808 21530
rect 36808 21518 36830 21530
rect 36896 21518 36898 21530
rect 36898 21518 36930 21530
rect 36996 21518 37030 21552
rect 37096 21518 37130 21552
rect 37196 21530 37230 21552
rect 37196 21518 37224 21530
rect 37224 21518 37230 21530
rect 36696 21440 36730 21452
rect 36796 21440 36830 21452
rect 36896 21440 36930 21452
rect 36696 21418 36718 21440
rect 36718 21418 36730 21440
rect 36796 21418 36808 21440
rect 36808 21418 36830 21440
rect 36896 21418 36898 21440
rect 36898 21418 36930 21440
rect 36996 21418 37030 21452
rect 37096 21418 37130 21452
rect 37196 21440 37230 21452
rect 37196 21418 37224 21440
rect 37224 21418 37230 21440
rect 37850 22122 37884 22156
rect 37940 22154 37974 22156
rect 38030 22154 38064 22156
rect 38120 22154 38154 22156
rect 38210 22154 38244 22156
rect 38300 22154 38334 22156
rect 38390 22154 38424 22156
rect 38480 22154 38514 22156
rect 38570 22154 38604 22156
rect 38660 22154 38694 22156
rect 37940 22122 37960 22154
rect 37960 22122 37974 22154
rect 38030 22122 38050 22154
rect 38050 22122 38064 22154
rect 38120 22122 38140 22154
rect 38140 22122 38154 22154
rect 38210 22122 38230 22154
rect 38230 22122 38244 22154
rect 38300 22122 38320 22154
rect 38320 22122 38334 22154
rect 38390 22122 38410 22154
rect 38410 22122 38424 22154
rect 38480 22122 38500 22154
rect 38500 22122 38514 22154
rect 38570 22122 38590 22154
rect 38590 22122 38604 22154
rect 38660 22122 38680 22154
rect 38680 22122 38694 22154
rect 38750 22122 38784 22156
rect 38036 21946 38058 21952
rect 38058 21946 38070 21952
rect 38136 21946 38148 21952
rect 38148 21946 38170 21952
rect 38236 21946 38238 21952
rect 38238 21946 38270 21952
rect 38036 21918 38070 21946
rect 38136 21918 38170 21946
rect 38236 21918 38270 21946
rect 38336 21918 38370 21952
rect 38436 21918 38470 21952
rect 38536 21946 38564 21952
rect 38564 21946 38570 21952
rect 38536 21918 38570 21946
rect 38036 21818 38070 21852
rect 38136 21818 38170 21852
rect 38236 21818 38270 21852
rect 38336 21818 38370 21852
rect 38436 21818 38470 21852
rect 38536 21818 38570 21852
rect 38036 21718 38070 21752
rect 38136 21718 38170 21752
rect 38236 21718 38270 21752
rect 38336 21718 38370 21752
rect 38436 21718 38470 21752
rect 38536 21718 38570 21752
rect 38036 21620 38070 21652
rect 38136 21620 38170 21652
rect 38236 21620 38270 21652
rect 38036 21618 38058 21620
rect 38058 21618 38070 21620
rect 38136 21618 38148 21620
rect 38148 21618 38170 21620
rect 38236 21618 38238 21620
rect 38238 21618 38270 21620
rect 38336 21618 38370 21652
rect 38436 21618 38470 21652
rect 38536 21620 38570 21652
rect 38536 21618 38564 21620
rect 38564 21618 38570 21620
rect 38036 21530 38070 21552
rect 38136 21530 38170 21552
rect 38236 21530 38270 21552
rect 38036 21518 38058 21530
rect 38058 21518 38070 21530
rect 38136 21518 38148 21530
rect 38148 21518 38170 21530
rect 38236 21518 38238 21530
rect 38238 21518 38270 21530
rect 38336 21518 38370 21552
rect 38436 21518 38470 21552
rect 38536 21530 38570 21552
rect 38536 21518 38564 21530
rect 38564 21518 38570 21530
rect 38036 21440 38070 21452
rect 38136 21440 38170 21452
rect 38236 21440 38270 21452
rect 38036 21418 38058 21440
rect 38058 21418 38070 21440
rect 38136 21418 38148 21440
rect 38148 21418 38170 21440
rect 38236 21418 38238 21440
rect 38238 21418 38270 21440
rect 38336 21418 38370 21452
rect 38436 21418 38470 21452
rect 38536 21440 38570 21452
rect 38536 21418 38564 21440
rect 38564 21418 38570 21440
rect 39765 21843 40159 22381
rect 41772 21843 42166 22381
rect 21097 21097 21131 21131
rect 26893 21097 26927 21131
rect 13277 20961 13311 20995
rect 8309 20893 8343 20927
rect 39765 20883 40159 21421
rect 41772 20883 42166 21421
rect 7863 20735 7897 20769
rect 8263 20735 8297 20769
rect 8663 20735 8697 20769
rect 9063 20735 9097 20769
rect 9463 20735 9497 20769
rect 9863 20735 9897 20769
rect 10263 20735 10297 20769
rect 10663 20735 10697 20769
rect 11063 20735 11097 20769
rect 11463 20735 11497 20769
rect 11863 20735 11897 20769
rect 12263 20735 12297 20769
rect 12663 20735 12697 20769
rect 13063 20735 13097 20769
rect 13745 20735 13779 20769
rect 14145 20735 14179 20769
rect 14545 20735 14579 20769
rect 14945 20735 14979 20769
rect 15345 20735 15379 20769
rect 15745 20735 15779 20769
rect 16145 20735 16179 20769
rect 16545 20735 16579 20769
rect 16945 20735 16979 20769
rect 17345 20735 17379 20769
rect 17745 20735 17779 20769
rect 18145 20735 18179 20769
rect 18545 20735 18579 20769
rect 18945 20735 18979 20769
rect 19345 20735 19379 20769
rect 19745 20735 19779 20769
rect 20145 20735 20179 20769
rect 20545 20735 20579 20769
rect 21191 20735 21225 20769
rect 21391 20735 21425 20769
rect 21591 20735 21625 20769
rect 21791 20735 21825 20769
rect 21991 20735 22025 20769
rect 22191 20735 22225 20769
rect 23151 20735 23185 20769
rect 23551 20735 23585 20769
rect 23951 20735 23985 20769
rect 24351 20735 24385 20769
rect 24751 20735 24785 20769
rect 25151 20735 25185 20769
rect 25551 20735 25585 20769
rect 25951 20735 25985 20769
rect 26351 20735 26385 20769
rect 26751 20735 26785 20769
rect 28443 20735 28477 20769
rect 28643 20735 28677 20769
rect 28843 20735 28877 20769
rect 29043 20735 29077 20769
rect 29243 20735 29277 20769
rect 29443 20735 29477 20769
rect 29643 20735 29677 20769
rect 29843 20735 29877 20769
rect 30043 20735 30077 20769
rect 30243 20735 30277 20769
rect 30443 20735 30477 20769
rect 30643 20735 30677 20769
rect 30843 20735 30877 20769
rect 31043 20735 31077 20769
rect 31243 20735 31277 20769
rect 31443 20735 31477 20769
rect 31643 20735 31677 20769
rect 31843 20735 31877 20769
rect 32043 20735 32077 20769
rect 32243 20735 32277 20769
rect 32443 20735 32477 20769
rect 32643 20735 32677 20769
rect 32843 20735 32877 20769
rect 33043 20735 33077 20769
rect 33243 20735 33277 20769
rect 33443 20735 33477 20769
rect 33643 20735 33677 20769
rect 33843 20735 33877 20769
rect 34043 20735 34077 20769
rect 34243 20735 34277 20769
rect 34443 20735 34477 20769
rect 34643 20735 34677 20769
rect 34843 20735 34877 20769
rect 35043 20735 35077 20769
rect 35243 20735 35277 20769
rect 35443 20735 35477 20769
rect 35643 20735 35677 20769
rect 35843 20735 35877 20769
rect 36043 20735 36077 20769
rect 36243 20735 36277 20769
rect 36443 20735 36477 20769
rect 36643 20735 36677 20769
rect 36843 20735 36877 20769
rect 37043 20735 37077 20769
rect 37243 20735 37277 20769
rect 37443 20735 37477 20769
rect 37643 20735 37677 20769
rect 37843 20735 37877 20769
rect 38043 20735 38077 20769
rect 38243 20735 38277 20769
rect 38443 20735 38477 20769
rect 38643 20735 38677 20769
rect 38843 20735 38877 20769
rect 39929 20735 39963 20769
rect 40129 20735 40163 20769
rect 40329 20735 40363 20769
rect 40529 20735 40563 20769
rect 40729 20735 40763 20769
rect 40929 20735 40963 20769
rect 41129 20735 41163 20769
rect 41329 20735 41363 20769
rect 41529 20735 41563 20769
rect 41729 20735 41763 20769
rect 41929 20735 41963 20769
rect 6197 18855 6231 18889
rect 6597 18855 6631 18889
rect 6997 18855 7031 18889
rect 7397 18855 7431 18889
rect 7797 18855 7831 18889
rect 8197 18855 8231 18889
rect 8597 18855 8631 18889
rect 8997 18855 9031 18889
rect 9397 18855 9431 18889
rect 9797 18855 9831 18889
rect 10823 18855 10857 18889
rect 11023 18855 11057 18889
rect 11223 18855 11257 18889
rect 11423 18855 11457 18889
rect 11623 18855 11657 18889
rect 11823 18855 11857 18889
rect 12023 18855 12057 18889
rect 12223 18855 12257 18889
rect 12423 18855 12457 18889
rect 12623 18855 12657 18889
rect 12823 18855 12857 18889
rect 13567 18855 13601 18889
rect 13767 18855 13801 18889
rect 13967 18855 14001 18889
rect 14167 18855 14201 18889
rect 14367 18855 14401 18889
rect 14567 18855 14601 18889
rect 14767 18855 14801 18889
rect 14967 18855 15001 18889
rect 15167 18855 15201 18889
rect 15367 18855 15401 18889
rect 15567 18855 15601 18889
rect 16293 18855 16327 18889
rect 16693 18855 16727 18889
rect 17093 18855 17127 18889
rect 17493 18855 17527 18889
rect 17893 18855 17927 18889
rect 18293 18855 18327 18889
rect 18693 18855 18727 18889
rect 19093 18855 19127 18889
rect 19493 18855 19527 18889
rect 19893 18855 19927 18889
rect 20293 18855 20327 18889
rect 20693 18855 20727 18889
rect 21093 18855 21127 18889
rect 21493 18855 21527 18889
rect 21893 18855 21927 18889
rect 22293 18855 22327 18889
rect 22693 18855 22727 18889
rect 23093 18855 23127 18889
rect 24131 18855 24165 18889
rect 24531 18855 24565 18889
rect 24931 18855 24965 18889
rect 25331 18855 25365 18889
rect 25731 18855 25765 18889
rect 26131 18855 26165 18889
rect 26531 18855 26565 18889
rect 28443 18855 28477 18889
rect 28643 18855 28677 18889
rect 28843 18855 28877 18889
rect 29043 18855 29077 18889
rect 29243 18855 29277 18889
rect 29443 18855 29477 18889
rect 29643 18855 29677 18889
rect 29843 18855 29877 18889
rect 30043 18855 30077 18889
rect 30243 18855 30277 18889
rect 30443 18855 30477 18889
rect 30643 18855 30677 18889
rect 30843 18855 30877 18889
rect 31043 18855 31077 18889
rect 31243 18855 31277 18889
rect 31443 18855 31477 18889
rect 31643 18855 31677 18889
rect 31843 18855 31877 18889
rect 32043 18855 32077 18889
rect 32243 18855 32277 18889
rect 32443 18855 32477 18889
rect 32643 18855 32677 18889
rect 32843 18855 32877 18889
rect 33043 18855 33077 18889
rect 33243 18855 33277 18889
rect 33443 18855 33477 18889
rect 33643 18855 33677 18889
rect 33843 18855 33877 18889
rect 34043 18855 34077 18889
rect 34243 18855 34277 18889
rect 34443 18855 34477 18889
rect 34643 18855 34677 18889
rect 34843 18855 34877 18889
rect 35043 18855 35077 18889
rect 35243 18855 35277 18889
rect 35443 18855 35477 18889
rect 35643 18855 35677 18889
rect 35843 18855 35877 18889
rect 36043 18855 36077 18889
rect 36243 18855 36277 18889
rect 36443 18855 36477 18889
rect 36643 18855 36677 18889
rect 36843 18855 36877 18889
rect 37043 18855 37077 18889
rect 37243 18855 37277 18889
rect 37443 18855 37477 18889
rect 37643 18855 37677 18889
rect 37843 18855 37877 18889
rect 38043 18855 38077 18889
rect 38243 18855 38277 18889
rect 38443 18855 38477 18889
rect 38643 18855 38677 18889
rect 38843 18855 38877 18889
rect 39439 18855 39473 18889
rect 39639 18855 39673 18889
rect 39839 18855 39873 18889
rect 40039 18855 40073 18889
rect 40239 18855 40273 18889
rect 40439 18855 40473 18889
rect 40639 18855 40673 18889
rect 40839 18855 40873 18889
rect 41039 18855 41073 18889
rect 41239 18855 41273 18889
rect 41439 18855 41473 18889
rect 6026 18349 6060 18369
rect 6026 18335 6060 18349
rect 6026 18281 6060 18297
rect 6026 18263 6060 18281
rect 6026 18213 6060 18225
rect 6026 18191 6060 18213
rect 6026 18145 6060 18153
rect 6026 18119 6060 18145
rect 6026 18077 6060 18081
rect 6026 18047 6060 18077
rect 6026 17975 6060 18009
rect 6026 17907 6060 17937
rect 6026 17903 6060 17907
rect 6026 17839 6060 17865
rect 6026 17831 6060 17839
rect 6026 17771 6060 17793
rect 6026 17759 6060 17771
rect 6026 17703 6060 17721
rect 6026 17687 6060 17703
rect 6026 17635 6060 17649
rect 6026 17615 6060 17635
rect 6484 18349 6518 18369
rect 6484 18335 6518 18349
rect 6484 18281 6518 18297
rect 6484 18263 6518 18281
rect 6484 18213 6518 18225
rect 6484 18191 6518 18213
rect 6484 18145 6518 18153
rect 6484 18119 6518 18145
rect 6484 18077 6518 18081
rect 6484 18047 6518 18077
rect 6484 17975 6518 18009
rect 6484 17907 6518 17937
rect 6484 17903 6518 17907
rect 6484 17839 6518 17865
rect 6484 17831 6518 17839
rect 6484 17771 6518 17793
rect 6484 17759 6518 17771
rect 6484 17703 6518 17721
rect 6484 17687 6518 17703
rect 6484 17635 6518 17649
rect 6942 18349 6976 18369
rect 6942 18335 6976 18349
rect 6942 18281 6976 18297
rect 6942 18263 6976 18281
rect 6942 18213 6976 18225
rect 6942 18191 6976 18213
rect 6942 18145 6976 18153
rect 6942 18119 6976 18145
rect 6942 18077 6976 18081
rect 6942 18047 6976 18077
rect 6942 17975 6976 18009
rect 6942 17907 6976 17937
rect 6942 17903 6976 17907
rect 6942 17839 6976 17865
rect 6942 17831 6976 17839
rect 6942 17771 6976 17793
rect 6942 17759 6976 17771
rect 6942 17703 6976 17721
rect 6942 17687 6976 17703
rect 6484 17615 6518 17635
rect 6942 17635 6976 17649
rect 6942 17615 6976 17635
rect 7400 18349 7434 18369
rect 7400 18335 7434 18349
rect 7400 18281 7434 18297
rect 7400 18263 7434 18281
rect 7400 18213 7434 18225
rect 7400 18191 7434 18213
rect 7400 18145 7434 18153
rect 7400 18119 7434 18145
rect 7400 18077 7434 18081
rect 7400 18047 7434 18077
rect 7400 17975 7434 18009
rect 7400 17907 7434 17937
rect 7400 17903 7434 17907
rect 7400 17839 7434 17865
rect 7400 17831 7434 17839
rect 7400 17771 7434 17793
rect 7400 17759 7434 17771
rect 7400 17703 7434 17721
rect 7400 17687 7434 17703
rect 7400 17635 7434 17649
rect 7858 18349 7892 18369
rect 7858 18335 7892 18349
rect 7858 18281 7892 18297
rect 7858 18263 7892 18281
rect 7858 18213 7892 18225
rect 7858 18191 7892 18213
rect 7858 18145 7892 18153
rect 7858 18119 7892 18145
rect 7858 18077 7892 18081
rect 7858 18047 7892 18077
rect 7858 17975 7892 18009
rect 7858 17907 7892 17937
rect 7858 17903 7892 17907
rect 7858 17839 7892 17865
rect 7858 17831 7892 17839
rect 7858 17771 7892 17793
rect 7858 17759 7892 17771
rect 7858 17703 7892 17721
rect 7858 17687 7892 17703
rect 7400 17615 7434 17635
rect 7858 17635 7892 17649
rect 7858 17615 7892 17635
rect 8316 18349 8350 18369
rect 8316 18335 8350 18349
rect 8316 18281 8350 18297
rect 8316 18263 8350 18281
rect 8316 18213 8350 18225
rect 8316 18191 8350 18213
rect 8316 18145 8350 18153
rect 8316 18119 8350 18145
rect 8316 18077 8350 18081
rect 8316 18047 8350 18077
rect 8316 17975 8350 18009
rect 8316 17907 8350 17937
rect 8316 17903 8350 17907
rect 8316 17839 8350 17865
rect 8316 17831 8350 17839
rect 8316 17771 8350 17793
rect 8316 17759 8350 17771
rect 8316 17703 8350 17721
rect 8316 17687 8350 17703
rect 8316 17635 8350 17649
rect 8774 18349 8808 18369
rect 8774 18335 8808 18349
rect 8774 18281 8808 18297
rect 8774 18263 8808 18281
rect 8774 18213 8808 18225
rect 8774 18191 8808 18213
rect 8774 18145 8808 18153
rect 8774 18119 8808 18145
rect 8774 18077 8808 18081
rect 8774 18047 8808 18077
rect 8774 17975 8808 18009
rect 8774 17907 8808 17937
rect 8774 17903 8808 17907
rect 8774 17839 8808 17865
rect 8774 17831 8808 17839
rect 8774 17771 8808 17793
rect 8774 17759 8808 17771
rect 8774 17703 8808 17721
rect 8774 17687 8808 17703
rect 8316 17615 8350 17635
rect 8774 17635 8808 17649
rect 8774 17615 8808 17635
rect 9232 18349 9266 18369
rect 9232 18335 9266 18349
rect 9232 18281 9266 18297
rect 9232 18263 9266 18281
rect 9232 18213 9266 18225
rect 9232 18191 9266 18213
rect 9232 18145 9266 18153
rect 9232 18119 9266 18145
rect 9232 18077 9266 18081
rect 9232 18047 9266 18077
rect 9232 17975 9266 18009
rect 9232 17907 9266 17937
rect 9232 17903 9266 17907
rect 9232 17839 9266 17865
rect 9232 17831 9266 17839
rect 9232 17771 9266 17793
rect 9232 17759 9266 17771
rect 9232 17703 9266 17721
rect 9232 17687 9266 17703
rect 9232 17635 9266 17649
rect 9690 18349 9724 18369
rect 9690 18335 9724 18349
rect 9690 18281 9724 18297
rect 9690 18263 9724 18281
rect 9690 18213 9724 18225
rect 9690 18191 9724 18213
rect 9690 18145 9724 18153
rect 9690 18119 9724 18145
rect 9690 18077 9724 18081
rect 9690 18047 9724 18077
rect 9690 17975 9724 18009
rect 9690 17907 9724 17937
rect 9690 17903 9724 17907
rect 9690 17839 9724 17865
rect 9690 17831 9724 17839
rect 9690 17771 9724 17793
rect 9690 17759 9724 17771
rect 9690 17703 9724 17721
rect 9690 17687 9724 17703
rect 9232 17615 9266 17635
rect 9690 17635 9724 17649
rect 9690 17615 9724 17635
rect 10148 18349 10182 18369
rect 10148 18335 10182 18349
rect 10148 18281 10182 18297
rect 10148 18263 10182 18281
rect 10148 18213 10182 18225
rect 10148 18191 10182 18213
rect 10148 18145 10182 18153
rect 10148 18119 10182 18145
rect 10148 18077 10182 18081
rect 10148 18047 10182 18077
rect 10659 18083 11053 18621
rect 12666 18083 13060 18621
rect 13403 18083 13797 18621
rect 26157 18683 26191 18717
rect 15410 18083 15804 18621
rect 10148 17975 10182 18009
rect 10148 17907 10182 17937
rect 10148 17903 10182 17907
rect 10148 17839 10182 17865
rect 10148 17831 10182 17839
rect 10148 17771 10182 17793
rect 10148 17759 10182 17771
rect 10148 17703 10182 17721
rect 10148 17687 10182 17703
rect 10148 17635 10182 17649
rect 10148 17615 10182 17635
rect 6101 17289 6135 17323
rect 10659 17123 11053 17661
rect 12666 17123 13060 17661
rect 13403 17123 13797 17661
rect 15410 17123 15804 17661
rect 23995 18587 24029 18621
rect 23995 18519 24029 18549
rect 23995 18515 24029 18519
rect 23995 18451 24029 18477
rect 23995 18443 24029 18451
rect 23995 18383 24029 18405
rect 23995 18371 24029 18383
rect 23995 18315 24029 18333
rect 23995 18299 24029 18315
rect 23995 18247 24029 18261
rect 23995 18227 24029 18247
rect 23995 18179 24029 18189
rect 23995 18155 24029 18179
rect 23995 18111 24029 18117
rect 23995 18083 24029 18111
rect 23995 18043 24029 18045
rect 23995 18011 24029 18043
rect 23995 17941 24029 17973
rect 23995 17939 24029 17941
rect 23995 17873 24029 17901
rect 23995 17867 24029 17873
rect 23995 17805 24029 17829
rect 23995 17795 24029 17805
rect 23995 17737 24029 17757
rect 23995 17723 24029 17737
rect 23995 17669 24029 17685
rect 23995 17651 24029 17669
rect 23995 17601 24029 17613
rect 23995 17579 24029 17601
rect 23995 17533 24029 17541
rect 23995 17507 24029 17533
rect 23995 17465 24029 17469
rect 23995 17435 24029 17465
rect 23995 17363 24029 17397
rect 24453 18587 24487 18621
rect 24453 18519 24487 18549
rect 24453 18515 24487 18519
rect 24453 18451 24487 18477
rect 24453 18443 24487 18451
rect 24453 18383 24487 18405
rect 24453 18371 24487 18383
rect 24453 18315 24487 18333
rect 24453 18299 24487 18315
rect 24453 18247 24487 18261
rect 24453 18227 24487 18247
rect 24453 18179 24487 18189
rect 24453 18155 24487 18179
rect 24453 18111 24487 18117
rect 24453 18083 24487 18111
rect 24453 18043 24487 18045
rect 24453 18011 24487 18043
rect 24453 17941 24487 17973
rect 24453 17939 24487 17941
rect 24453 17873 24487 17901
rect 24453 17867 24487 17873
rect 24453 17805 24487 17829
rect 24453 17795 24487 17805
rect 24453 17737 24487 17757
rect 24453 17723 24487 17737
rect 24453 17669 24487 17685
rect 24453 17651 24487 17669
rect 24453 17601 24487 17613
rect 24453 17579 24487 17601
rect 24453 17533 24487 17541
rect 24453 17507 24487 17533
rect 24453 17465 24487 17469
rect 24453 17435 24487 17465
rect 24453 17363 24487 17397
rect 24911 18587 24945 18621
rect 24911 18519 24945 18549
rect 24911 18515 24945 18519
rect 24911 18451 24945 18477
rect 24911 18443 24945 18451
rect 24911 18383 24945 18405
rect 24911 18371 24945 18383
rect 24911 18315 24945 18333
rect 24911 18299 24945 18315
rect 24911 18247 24945 18261
rect 24911 18227 24945 18247
rect 24911 18179 24945 18189
rect 24911 18155 24945 18179
rect 24911 18111 24945 18117
rect 24911 18083 24945 18111
rect 24911 18043 24945 18045
rect 24911 18011 24945 18043
rect 24911 17941 24945 17973
rect 24911 17939 24945 17941
rect 24911 17873 24945 17901
rect 24911 17867 24945 17873
rect 24911 17805 24945 17829
rect 24911 17795 24945 17805
rect 24911 17737 24945 17757
rect 24911 17723 24945 17737
rect 24911 17669 24945 17685
rect 24911 17651 24945 17669
rect 24911 17601 24945 17613
rect 24911 17579 24945 17601
rect 24911 17533 24945 17541
rect 24911 17507 24945 17533
rect 24911 17465 24945 17469
rect 24911 17435 24945 17465
rect 24911 17363 24945 17397
rect 25369 18587 25403 18621
rect 25369 18519 25403 18549
rect 25369 18515 25403 18519
rect 25369 18451 25403 18477
rect 25369 18443 25403 18451
rect 25369 18383 25403 18405
rect 25369 18371 25403 18383
rect 25369 18315 25403 18333
rect 25369 18299 25403 18315
rect 25369 18247 25403 18261
rect 25369 18227 25403 18247
rect 25369 18179 25403 18189
rect 25369 18155 25403 18179
rect 25369 18111 25403 18117
rect 25369 18083 25403 18111
rect 25369 18043 25403 18045
rect 25369 18011 25403 18043
rect 25369 17941 25403 17973
rect 25369 17939 25403 17941
rect 25369 17873 25403 17901
rect 25369 17867 25403 17873
rect 25369 17805 25403 17829
rect 25369 17795 25403 17805
rect 25369 17737 25403 17757
rect 25369 17723 25403 17737
rect 25369 17669 25403 17685
rect 25369 17651 25403 17669
rect 25369 17601 25403 17613
rect 25369 17579 25403 17601
rect 25369 17533 25403 17541
rect 25369 17507 25403 17533
rect 25369 17465 25403 17469
rect 25369 17435 25403 17465
rect 25369 17363 25403 17397
rect 25827 18587 25861 18621
rect 25827 18519 25861 18549
rect 25827 18515 25861 18519
rect 25827 18451 25861 18477
rect 25827 18443 25861 18451
rect 25827 18383 25861 18405
rect 25827 18371 25861 18383
rect 25827 18315 25861 18333
rect 25827 18299 25861 18315
rect 25827 18247 25861 18261
rect 25827 18227 25861 18247
rect 25827 18179 25861 18189
rect 25827 18155 25861 18179
rect 25827 18111 25861 18117
rect 25827 18083 25861 18111
rect 25827 18043 25861 18045
rect 25827 18011 25861 18043
rect 25827 17941 25861 17973
rect 25827 17939 25861 17941
rect 25827 17873 25861 17901
rect 25827 17867 25861 17873
rect 25827 17805 25861 17829
rect 25827 17795 25861 17805
rect 25827 17737 25861 17757
rect 25827 17723 25861 17737
rect 25827 17669 25861 17685
rect 25827 17651 25861 17669
rect 25827 17601 25861 17613
rect 25827 17579 25861 17601
rect 25827 17533 25861 17541
rect 25827 17507 25861 17533
rect 25827 17465 25861 17469
rect 25827 17435 25861 17465
rect 25827 17363 25861 17397
rect 26285 18587 26319 18621
rect 26285 18519 26319 18549
rect 26285 18515 26319 18519
rect 26285 18451 26319 18477
rect 26285 18443 26319 18451
rect 26285 18383 26319 18405
rect 26285 18371 26319 18383
rect 26285 18315 26319 18333
rect 26285 18299 26319 18315
rect 26285 18247 26319 18261
rect 26285 18227 26319 18247
rect 26285 18179 26319 18189
rect 26285 18155 26319 18179
rect 26285 18111 26319 18117
rect 26285 18083 26319 18111
rect 26285 18043 26319 18045
rect 26285 18011 26319 18043
rect 26285 17941 26319 17973
rect 26285 17939 26319 17941
rect 26285 17873 26319 17901
rect 26285 17867 26319 17873
rect 26285 17805 26319 17829
rect 26285 17795 26319 17805
rect 26285 17737 26319 17757
rect 26285 17723 26319 17737
rect 26285 17669 26319 17685
rect 26285 17651 26319 17669
rect 26285 17601 26319 17613
rect 26285 17579 26319 17601
rect 26285 17533 26319 17541
rect 26285 17507 26319 17533
rect 26285 17465 26319 17469
rect 26285 17435 26319 17465
rect 26285 17363 26319 17397
rect 26743 18587 26777 18621
rect 26743 18519 26777 18549
rect 26743 18515 26777 18519
rect 26743 18451 26777 18477
rect 26743 18443 26777 18451
rect 26743 18383 26777 18405
rect 26743 18371 26777 18383
rect 26743 18315 26777 18333
rect 26743 18299 26777 18315
rect 26743 18247 26777 18261
rect 26743 18227 26777 18247
rect 26743 18179 26777 18189
rect 26743 18155 26777 18179
rect 26743 18111 26777 18117
rect 26743 18083 26777 18111
rect 26743 18043 26777 18045
rect 26743 18011 26777 18043
rect 26743 17941 26777 17973
rect 26743 17939 26777 17941
rect 26743 17873 26777 17901
rect 26743 17867 26777 17873
rect 26743 17805 26777 17829
rect 26743 17795 26777 17805
rect 26743 17737 26777 17757
rect 26743 17723 26777 17737
rect 26743 17669 26777 17685
rect 26743 17651 26777 17669
rect 26743 17601 26777 17613
rect 26743 17579 26777 17601
rect 26743 17533 26777 17541
rect 26743 17507 26777 17533
rect 26743 17465 26777 17469
rect 26743 17435 26777 17465
rect 26743 17363 26777 17397
rect 28306 18522 28340 18556
rect 28396 18541 28430 18556
rect 28486 18541 28520 18556
rect 28576 18541 28610 18556
rect 28666 18541 28700 18556
rect 28756 18541 28790 18556
rect 28846 18541 28880 18556
rect 28936 18541 28970 18556
rect 29026 18541 29060 18556
rect 29116 18541 29150 18556
rect 29206 18541 29240 18556
rect 29296 18541 29330 18556
rect 29386 18541 29420 18556
rect 28396 18522 28416 18541
rect 28416 18522 28430 18541
rect 28486 18522 28506 18541
rect 28506 18522 28520 18541
rect 28576 18522 28596 18541
rect 28596 18522 28610 18541
rect 28666 18522 28686 18541
rect 28686 18522 28700 18541
rect 28756 18522 28776 18541
rect 28776 18522 28790 18541
rect 28846 18522 28866 18541
rect 28866 18522 28880 18541
rect 28936 18522 28956 18541
rect 28956 18522 28970 18541
rect 29026 18522 29046 18541
rect 29046 18522 29060 18541
rect 29116 18522 29136 18541
rect 29136 18522 29150 18541
rect 29206 18522 29226 18541
rect 29226 18522 29240 18541
rect 29296 18522 29316 18541
rect 29316 18522 29330 18541
rect 29386 18522 29406 18541
rect 29406 18522 29420 18541
rect 29476 18522 29510 18556
rect 29646 18522 29680 18556
rect 29736 18541 29770 18556
rect 29826 18541 29860 18556
rect 29916 18541 29950 18556
rect 30006 18541 30040 18556
rect 30096 18541 30130 18556
rect 30186 18541 30220 18556
rect 30276 18541 30310 18556
rect 30366 18541 30400 18556
rect 30456 18541 30490 18556
rect 30546 18541 30580 18556
rect 30636 18541 30670 18556
rect 30726 18541 30760 18556
rect 29736 18522 29756 18541
rect 29756 18522 29770 18541
rect 29826 18522 29846 18541
rect 29846 18522 29860 18541
rect 29916 18522 29936 18541
rect 29936 18522 29950 18541
rect 30006 18522 30026 18541
rect 30026 18522 30040 18541
rect 30096 18522 30116 18541
rect 30116 18522 30130 18541
rect 30186 18522 30206 18541
rect 30206 18522 30220 18541
rect 30276 18522 30296 18541
rect 30296 18522 30310 18541
rect 30366 18522 30386 18541
rect 30386 18522 30400 18541
rect 30456 18522 30476 18541
rect 30476 18522 30490 18541
rect 30546 18522 30566 18541
rect 30566 18522 30580 18541
rect 30636 18522 30656 18541
rect 30656 18522 30670 18541
rect 30726 18522 30746 18541
rect 30746 18522 30760 18541
rect 30816 18522 30850 18556
rect 30986 18522 31020 18556
rect 31076 18541 31110 18556
rect 31166 18541 31200 18556
rect 31256 18541 31290 18556
rect 31346 18541 31380 18556
rect 31436 18541 31470 18556
rect 31526 18541 31560 18556
rect 31616 18541 31650 18556
rect 31706 18541 31740 18556
rect 31796 18541 31830 18556
rect 31886 18541 31920 18556
rect 31976 18541 32010 18556
rect 32066 18541 32100 18556
rect 31076 18522 31096 18541
rect 31096 18522 31110 18541
rect 31166 18522 31186 18541
rect 31186 18522 31200 18541
rect 31256 18522 31276 18541
rect 31276 18522 31290 18541
rect 31346 18522 31366 18541
rect 31366 18522 31380 18541
rect 31436 18522 31456 18541
rect 31456 18522 31470 18541
rect 31526 18522 31546 18541
rect 31546 18522 31560 18541
rect 31616 18522 31636 18541
rect 31636 18522 31650 18541
rect 31706 18522 31726 18541
rect 31726 18522 31740 18541
rect 31796 18522 31816 18541
rect 31816 18522 31830 18541
rect 31886 18522 31906 18541
rect 31906 18522 31920 18541
rect 31976 18522 31996 18541
rect 31996 18522 32010 18541
rect 32066 18522 32086 18541
rect 32086 18522 32100 18541
rect 32156 18522 32190 18556
rect 32326 18522 32360 18556
rect 32416 18541 32450 18556
rect 32506 18541 32540 18556
rect 32596 18541 32630 18556
rect 32686 18541 32720 18556
rect 32776 18541 32810 18556
rect 32866 18541 32900 18556
rect 32956 18541 32990 18556
rect 33046 18541 33080 18556
rect 33136 18541 33170 18556
rect 33226 18541 33260 18556
rect 33316 18541 33350 18556
rect 33406 18541 33440 18556
rect 32416 18522 32436 18541
rect 32436 18522 32450 18541
rect 32506 18522 32526 18541
rect 32526 18522 32540 18541
rect 32596 18522 32616 18541
rect 32616 18522 32630 18541
rect 32686 18522 32706 18541
rect 32706 18522 32720 18541
rect 32776 18522 32796 18541
rect 32796 18522 32810 18541
rect 32866 18522 32886 18541
rect 32886 18522 32900 18541
rect 32956 18522 32976 18541
rect 32976 18522 32990 18541
rect 33046 18522 33066 18541
rect 33066 18522 33080 18541
rect 33136 18522 33156 18541
rect 33156 18522 33170 18541
rect 33226 18522 33246 18541
rect 33246 18522 33260 18541
rect 33316 18522 33336 18541
rect 33336 18522 33350 18541
rect 33406 18522 33426 18541
rect 33426 18522 33440 18541
rect 33496 18522 33530 18556
rect 33666 18522 33700 18556
rect 33756 18541 33790 18556
rect 33846 18541 33880 18556
rect 33936 18541 33970 18556
rect 34026 18541 34060 18556
rect 34116 18541 34150 18556
rect 34206 18541 34240 18556
rect 34296 18541 34330 18556
rect 34386 18541 34420 18556
rect 34476 18541 34510 18556
rect 34566 18541 34600 18556
rect 34656 18541 34690 18556
rect 34746 18541 34780 18556
rect 33756 18522 33776 18541
rect 33776 18522 33790 18541
rect 33846 18522 33866 18541
rect 33866 18522 33880 18541
rect 33936 18522 33956 18541
rect 33956 18522 33970 18541
rect 34026 18522 34046 18541
rect 34046 18522 34060 18541
rect 34116 18522 34136 18541
rect 34136 18522 34150 18541
rect 34206 18522 34226 18541
rect 34226 18522 34240 18541
rect 34296 18522 34316 18541
rect 34316 18522 34330 18541
rect 34386 18522 34406 18541
rect 34406 18522 34420 18541
rect 34476 18522 34496 18541
rect 34496 18522 34510 18541
rect 34566 18522 34586 18541
rect 34586 18522 34600 18541
rect 34656 18522 34676 18541
rect 34676 18522 34690 18541
rect 34746 18522 34766 18541
rect 34766 18522 34780 18541
rect 34836 18522 34870 18556
rect 35006 18522 35040 18556
rect 35096 18541 35130 18556
rect 35186 18541 35220 18556
rect 35276 18541 35310 18556
rect 35366 18541 35400 18556
rect 35456 18541 35490 18556
rect 35546 18541 35580 18556
rect 35636 18541 35670 18556
rect 35726 18541 35760 18556
rect 35816 18541 35850 18556
rect 35906 18541 35940 18556
rect 35996 18541 36030 18556
rect 36086 18541 36120 18556
rect 35096 18522 35116 18541
rect 35116 18522 35130 18541
rect 35186 18522 35206 18541
rect 35206 18522 35220 18541
rect 35276 18522 35296 18541
rect 35296 18522 35310 18541
rect 35366 18522 35386 18541
rect 35386 18522 35400 18541
rect 35456 18522 35476 18541
rect 35476 18522 35490 18541
rect 35546 18522 35566 18541
rect 35566 18522 35580 18541
rect 35636 18522 35656 18541
rect 35656 18522 35670 18541
rect 35726 18522 35746 18541
rect 35746 18522 35760 18541
rect 35816 18522 35836 18541
rect 35836 18522 35850 18541
rect 35906 18522 35926 18541
rect 35926 18522 35940 18541
rect 35996 18522 36016 18541
rect 36016 18522 36030 18541
rect 36086 18522 36106 18541
rect 36106 18522 36120 18541
rect 36176 18522 36210 18556
rect 36346 18522 36380 18556
rect 36436 18541 36470 18556
rect 36526 18541 36560 18556
rect 36616 18541 36650 18556
rect 36706 18541 36740 18556
rect 36796 18541 36830 18556
rect 36886 18541 36920 18556
rect 36976 18541 37010 18556
rect 37066 18541 37100 18556
rect 37156 18541 37190 18556
rect 37246 18541 37280 18556
rect 37336 18541 37370 18556
rect 37426 18541 37460 18556
rect 36436 18522 36456 18541
rect 36456 18522 36470 18541
rect 36526 18522 36546 18541
rect 36546 18522 36560 18541
rect 36616 18522 36636 18541
rect 36636 18522 36650 18541
rect 36706 18522 36726 18541
rect 36726 18522 36740 18541
rect 36796 18522 36816 18541
rect 36816 18522 36830 18541
rect 36886 18522 36906 18541
rect 36906 18522 36920 18541
rect 36976 18522 36996 18541
rect 36996 18522 37010 18541
rect 37066 18522 37086 18541
rect 37086 18522 37100 18541
rect 37156 18522 37176 18541
rect 37176 18522 37190 18541
rect 37246 18522 37266 18541
rect 37266 18522 37280 18541
rect 37336 18522 37356 18541
rect 37356 18522 37370 18541
rect 37426 18522 37446 18541
rect 37446 18522 37460 18541
rect 37516 18522 37550 18556
rect 37686 18522 37720 18556
rect 37776 18541 37810 18556
rect 37866 18541 37900 18556
rect 37956 18541 37990 18556
rect 38046 18541 38080 18556
rect 38136 18541 38170 18556
rect 38226 18541 38260 18556
rect 38316 18541 38350 18556
rect 38406 18541 38440 18556
rect 38496 18541 38530 18556
rect 38586 18541 38620 18556
rect 38676 18541 38710 18556
rect 38766 18541 38800 18556
rect 37776 18522 37796 18541
rect 37796 18522 37810 18541
rect 37866 18522 37886 18541
rect 37886 18522 37900 18541
rect 37956 18522 37976 18541
rect 37976 18522 37990 18541
rect 38046 18522 38066 18541
rect 38066 18522 38080 18541
rect 38136 18522 38156 18541
rect 38156 18522 38170 18541
rect 38226 18522 38246 18541
rect 38246 18522 38260 18541
rect 38316 18522 38336 18541
rect 38336 18522 38350 18541
rect 38406 18522 38426 18541
rect 38426 18522 38440 18541
rect 38496 18522 38516 18541
rect 38516 18522 38530 18541
rect 38586 18522 38606 18541
rect 38606 18522 38620 18541
rect 38676 18522 38696 18541
rect 38696 18522 38710 18541
rect 38766 18522 38786 18541
rect 38786 18522 38800 18541
rect 38856 18522 38890 18556
rect 28470 18362 28504 18396
rect 28560 18394 28594 18396
rect 28650 18394 28684 18396
rect 28740 18394 28774 18396
rect 28830 18394 28864 18396
rect 28920 18394 28954 18396
rect 29010 18394 29044 18396
rect 29100 18394 29134 18396
rect 29190 18394 29224 18396
rect 29280 18394 29314 18396
rect 28560 18362 28580 18394
rect 28580 18362 28594 18394
rect 28650 18362 28670 18394
rect 28670 18362 28684 18394
rect 28740 18362 28760 18394
rect 28760 18362 28774 18394
rect 28830 18362 28850 18394
rect 28850 18362 28864 18394
rect 28920 18362 28940 18394
rect 28940 18362 28954 18394
rect 29010 18362 29030 18394
rect 29030 18362 29044 18394
rect 29100 18362 29120 18394
rect 29120 18362 29134 18394
rect 29190 18362 29210 18394
rect 29210 18362 29224 18394
rect 29280 18362 29300 18394
rect 29300 18362 29314 18394
rect 29370 18362 29404 18396
rect 28656 18186 28678 18192
rect 28678 18186 28690 18192
rect 28756 18186 28768 18192
rect 28768 18186 28790 18192
rect 28856 18186 28858 18192
rect 28858 18186 28890 18192
rect 28656 18158 28690 18186
rect 28756 18158 28790 18186
rect 28856 18158 28890 18186
rect 28956 18158 28990 18192
rect 29056 18158 29090 18192
rect 29156 18186 29184 18192
rect 29184 18186 29190 18192
rect 29156 18158 29190 18186
rect 28656 18058 28690 18092
rect 28756 18058 28790 18092
rect 28856 18058 28890 18092
rect 28956 18058 28990 18092
rect 29056 18058 29090 18092
rect 29156 18058 29190 18092
rect 28656 17958 28690 17992
rect 28756 17958 28790 17992
rect 28856 17958 28890 17992
rect 28956 17958 28990 17992
rect 29056 17958 29090 17992
rect 29156 17958 29190 17992
rect 28656 17860 28690 17892
rect 28756 17860 28790 17892
rect 28856 17860 28890 17892
rect 28656 17858 28678 17860
rect 28678 17858 28690 17860
rect 28756 17858 28768 17860
rect 28768 17858 28790 17860
rect 28856 17858 28858 17860
rect 28858 17858 28890 17860
rect 28956 17858 28990 17892
rect 29056 17858 29090 17892
rect 29156 17860 29190 17892
rect 29156 17858 29184 17860
rect 29184 17858 29190 17860
rect 28656 17770 28690 17792
rect 28756 17770 28790 17792
rect 28856 17770 28890 17792
rect 28656 17758 28678 17770
rect 28678 17758 28690 17770
rect 28756 17758 28768 17770
rect 28768 17758 28790 17770
rect 28856 17758 28858 17770
rect 28858 17758 28890 17770
rect 28956 17758 28990 17792
rect 29056 17758 29090 17792
rect 29156 17770 29190 17792
rect 29156 17758 29184 17770
rect 29184 17758 29190 17770
rect 28656 17680 28690 17692
rect 28756 17680 28790 17692
rect 28856 17680 28890 17692
rect 28656 17658 28678 17680
rect 28678 17658 28690 17680
rect 28756 17658 28768 17680
rect 28768 17658 28790 17680
rect 28856 17658 28858 17680
rect 28858 17658 28890 17680
rect 28956 17658 28990 17692
rect 29056 17658 29090 17692
rect 29156 17680 29190 17692
rect 29156 17658 29184 17680
rect 29184 17658 29190 17680
rect 29810 18362 29844 18396
rect 29900 18394 29934 18396
rect 29990 18394 30024 18396
rect 30080 18394 30114 18396
rect 30170 18394 30204 18396
rect 30260 18394 30294 18396
rect 30350 18394 30384 18396
rect 30440 18394 30474 18396
rect 30530 18394 30564 18396
rect 30620 18394 30654 18396
rect 29900 18362 29920 18394
rect 29920 18362 29934 18394
rect 29990 18362 30010 18394
rect 30010 18362 30024 18394
rect 30080 18362 30100 18394
rect 30100 18362 30114 18394
rect 30170 18362 30190 18394
rect 30190 18362 30204 18394
rect 30260 18362 30280 18394
rect 30280 18362 30294 18394
rect 30350 18362 30370 18394
rect 30370 18362 30384 18394
rect 30440 18362 30460 18394
rect 30460 18362 30474 18394
rect 30530 18362 30550 18394
rect 30550 18362 30564 18394
rect 30620 18362 30640 18394
rect 30640 18362 30654 18394
rect 30710 18362 30744 18396
rect 29996 18186 30018 18192
rect 30018 18186 30030 18192
rect 30096 18186 30108 18192
rect 30108 18186 30130 18192
rect 30196 18186 30198 18192
rect 30198 18186 30230 18192
rect 29996 18158 30030 18186
rect 30096 18158 30130 18186
rect 30196 18158 30230 18186
rect 30296 18158 30330 18192
rect 30396 18158 30430 18192
rect 30496 18186 30524 18192
rect 30524 18186 30530 18192
rect 30496 18158 30530 18186
rect 29996 18058 30030 18092
rect 30096 18058 30130 18092
rect 30196 18058 30230 18092
rect 30296 18058 30330 18092
rect 30396 18058 30430 18092
rect 30496 18058 30530 18092
rect 29996 17958 30030 17992
rect 30096 17958 30130 17992
rect 30196 17958 30230 17992
rect 30296 17958 30330 17992
rect 30396 17958 30430 17992
rect 30496 17958 30530 17992
rect 29996 17860 30030 17892
rect 30096 17860 30130 17892
rect 30196 17860 30230 17892
rect 29996 17858 30018 17860
rect 30018 17858 30030 17860
rect 30096 17858 30108 17860
rect 30108 17858 30130 17860
rect 30196 17858 30198 17860
rect 30198 17858 30230 17860
rect 30296 17858 30330 17892
rect 30396 17858 30430 17892
rect 30496 17860 30530 17892
rect 30496 17858 30524 17860
rect 30524 17858 30530 17860
rect 29996 17770 30030 17792
rect 30096 17770 30130 17792
rect 30196 17770 30230 17792
rect 29996 17758 30018 17770
rect 30018 17758 30030 17770
rect 30096 17758 30108 17770
rect 30108 17758 30130 17770
rect 30196 17758 30198 17770
rect 30198 17758 30230 17770
rect 30296 17758 30330 17792
rect 30396 17758 30430 17792
rect 30496 17770 30530 17792
rect 30496 17758 30524 17770
rect 30524 17758 30530 17770
rect 29996 17680 30030 17692
rect 30096 17680 30130 17692
rect 30196 17680 30230 17692
rect 29996 17658 30018 17680
rect 30018 17658 30030 17680
rect 30096 17658 30108 17680
rect 30108 17658 30130 17680
rect 30196 17658 30198 17680
rect 30198 17658 30230 17680
rect 30296 17658 30330 17692
rect 30396 17658 30430 17692
rect 30496 17680 30530 17692
rect 30496 17658 30524 17680
rect 30524 17658 30530 17680
rect 31150 18362 31184 18396
rect 31240 18394 31274 18396
rect 31330 18394 31364 18396
rect 31420 18394 31454 18396
rect 31510 18394 31544 18396
rect 31600 18394 31634 18396
rect 31690 18394 31724 18396
rect 31780 18394 31814 18396
rect 31870 18394 31904 18396
rect 31960 18394 31994 18396
rect 31240 18362 31260 18394
rect 31260 18362 31274 18394
rect 31330 18362 31350 18394
rect 31350 18362 31364 18394
rect 31420 18362 31440 18394
rect 31440 18362 31454 18394
rect 31510 18362 31530 18394
rect 31530 18362 31544 18394
rect 31600 18362 31620 18394
rect 31620 18362 31634 18394
rect 31690 18362 31710 18394
rect 31710 18362 31724 18394
rect 31780 18362 31800 18394
rect 31800 18362 31814 18394
rect 31870 18362 31890 18394
rect 31890 18362 31904 18394
rect 31960 18362 31980 18394
rect 31980 18362 31994 18394
rect 32050 18362 32084 18396
rect 31336 18186 31358 18192
rect 31358 18186 31370 18192
rect 31436 18186 31448 18192
rect 31448 18186 31470 18192
rect 31536 18186 31538 18192
rect 31538 18186 31570 18192
rect 31336 18158 31370 18186
rect 31436 18158 31470 18186
rect 31536 18158 31570 18186
rect 31636 18158 31670 18192
rect 31736 18158 31770 18192
rect 31836 18186 31864 18192
rect 31864 18186 31870 18192
rect 31836 18158 31870 18186
rect 31336 18058 31370 18092
rect 31436 18058 31470 18092
rect 31536 18058 31570 18092
rect 31636 18058 31670 18092
rect 31736 18058 31770 18092
rect 31836 18058 31870 18092
rect 31336 17958 31370 17992
rect 31436 17958 31470 17992
rect 31536 17958 31570 17992
rect 31636 17958 31670 17992
rect 31736 17958 31770 17992
rect 31836 17958 31870 17992
rect 31336 17860 31370 17892
rect 31436 17860 31470 17892
rect 31536 17860 31570 17892
rect 31336 17858 31358 17860
rect 31358 17858 31370 17860
rect 31436 17858 31448 17860
rect 31448 17858 31470 17860
rect 31536 17858 31538 17860
rect 31538 17858 31570 17860
rect 31636 17858 31670 17892
rect 31736 17858 31770 17892
rect 31836 17860 31870 17892
rect 31836 17858 31864 17860
rect 31864 17858 31870 17860
rect 31336 17770 31370 17792
rect 31436 17770 31470 17792
rect 31536 17770 31570 17792
rect 31336 17758 31358 17770
rect 31358 17758 31370 17770
rect 31436 17758 31448 17770
rect 31448 17758 31470 17770
rect 31536 17758 31538 17770
rect 31538 17758 31570 17770
rect 31636 17758 31670 17792
rect 31736 17758 31770 17792
rect 31836 17770 31870 17792
rect 31836 17758 31864 17770
rect 31864 17758 31870 17770
rect 31336 17680 31370 17692
rect 31436 17680 31470 17692
rect 31536 17680 31570 17692
rect 31336 17658 31358 17680
rect 31358 17658 31370 17680
rect 31436 17658 31448 17680
rect 31448 17658 31470 17680
rect 31536 17658 31538 17680
rect 31538 17658 31570 17680
rect 31636 17658 31670 17692
rect 31736 17658 31770 17692
rect 31836 17680 31870 17692
rect 31836 17658 31864 17680
rect 31864 17658 31870 17680
rect 32490 18362 32524 18396
rect 32580 18394 32614 18396
rect 32670 18394 32704 18396
rect 32760 18394 32794 18396
rect 32850 18394 32884 18396
rect 32940 18394 32974 18396
rect 33030 18394 33064 18396
rect 33120 18394 33154 18396
rect 33210 18394 33244 18396
rect 33300 18394 33334 18396
rect 32580 18362 32600 18394
rect 32600 18362 32614 18394
rect 32670 18362 32690 18394
rect 32690 18362 32704 18394
rect 32760 18362 32780 18394
rect 32780 18362 32794 18394
rect 32850 18362 32870 18394
rect 32870 18362 32884 18394
rect 32940 18362 32960 18394
rect 32960 18362 32974 18394
rect 33030 18362 33050 18394
rect 33050 18362 33064 18394
rect 33120 18362 33140 18394
rect 33140 18362 33154 18394
rect 33210 18362 33230 18394
rect 33230 18362 33244 18394
rect 33300 18362 33320 18394
rect 33320 18362 33334 18394
rect 33390 18362 33424 18396
rect 32676 18186 32698 18192
rect 32698 18186 32710 18192
rect 32776 18186 32788 18192
rect 32788 18186 32810 18192
rect 32876 18186 32878 18192
rect 32878 18186 32910 18192
rect 32676 18158 32710 18186
rect 32776 18158 32810 18186
rect 32876 18158 32910 18186
rect 32976 18158 33010 18192
rect 33076 18158 33110 18192
rect 33176 18186 33204 18192
rect 33204 18186 33210 18192
rect 33176 18158 33210 18186
rect 32676 18058 32710 18092
rect 32776 18058 32810 18092
rect 32876 18058 32910 18092
rect 32976 18058 33010 18092
rect 33076 18058 33110 18092
rect 33176 18058 33210 18092
rect 32676 17958 32710 17992
rect 32776 17958 32810 17992
rect 32876 17958 32910 17992
rect 32976 17958 33010 17992
rect 33076 17958 33110 17992
rect 33176 17958 33210 17992
rect 32676 17860 32710 17892
rect 32776 17860 32810 17892
rect 32876 17860 32910 17892
rect 32676 17858 32698 17860
rect 32698 17858 32710 17860
rect 32776 17858 32788 17860
rect 32788 17858 32810 17860
rect 32876 17858 32878 17860
rect 32878 17858 32910 17860
rect 32976 17858 33010 17892
rect 33076 17858 33110 17892
rect 33176 17860 33210 17892
rect 33176 17858 33204 17860
rect 33204 17858 33210 17860
rect 32676 17770 32710 17792
rect 32776 17770 32810 17792
rect 32876 17770 32910 17792
rect 32676 17758 32698 17770
rect 32698 17758 32710 17770
rect 32776 17758 32788 17770
rect 32788 17758 32810 17770
rect 32876 17758 32878 17770
rect 32878 17758 32910 17770
rect 32976 17758 33010 17792
rect 33076 17758 33110 17792
rect 33176 17770 33210 17792
rect 33176 17758 33204 17770
rect 33204 17758 33210 17770
rect 32676 17680 32710 17692
rect 32776 17680 32810 17692
rect 32876 17680 32910 17692
rect 32676 17658 32698 17680
rect 32698 17658 32710 17680
rect 32776 17658 32788 17680
rect 32788 17658 32810 17680
rect 32876 17658 32878 17680
rect 32878 17658 32910 17680
rect 32976 17658 33010 17692
rect 33076 17658 33110 17692
rect 33176 17680 33210 17692
rect 33176 17658 33204 17680
rect 33204 17658 33210 17680
rect 33830 18362 33864 18396
rect 33920 18394 33954 18396
rect 34010 18394 34044 18396
rect 34100 18394 34134 18396
rect 34190 18394 34224 18396
rect 34280 18394 34314 18396
rect 34370 18394 34404 18396
rect 34460 18394 34494 18396
rect 34550 18394 34584 18396
rect 34640 18394 34674 18396
rect 33920 18362 33940 18394
rect 33940 18362 33954 18394
rect 34010 18362 34030 18394
rect 34030 18362 34044 18394
rect 34100 18362 34120 18394
rect 34120 18362 34134 18394
rect 34190 18362 34210 18394
rect 34210 18362 34224 18394
rect 34280 18362 34300 18394
rect 34300 18362 34314 18394
rect 34370 18362 34390 18394
rect 34390 18362 34404 18394
rect 34460 18362 34480 18394
rect 34480 18362 34494 18394
rect 34550 18362 34570 18394
rect 34570 18362 34584 18394
rect 34640 18362 34660 18394
rect 34660 18362 34674 18394
rect 34730 18362 34764 18396
rect 34016 18186 34038 18192
rect 34038 18186 34050 18192
rect 34116 18186 34128 18192
rect 34128 18186 34150 18192
rect 34216 18186 34218 18192
rect 34218 18186 34250 18192
rect 34016 18158 34050 18186
rect 34116 18158 34150 18186
rect 34216 18158 34250 18186
rect 34316 18158 34350 18192
rect 34416 18158 34450 18192
rect 34516 18186 34544 18192
rect 34544 18186 34550 18192
rect 34516 18158 34550 18186
rect 34016 18058 34050 18092
rect 34116 18058 34150 18092
rect 34216 18058 34250 18092
rect 34316 18058 34350 18092
rect 34416 18058 34450 18092
rect 34516 18058 34550 18092
rect 34016 17958 34050 17992
rect 34116 17958 34150 17992
rect 34216 17958 34250 17992
rect 34316 17958 34350 17992
rect 34416 17958 34450 17992
rect 34516 17958 34550 17992
rect 34016 17860 34050 17892
rect 34116 17860 34150 17892
rect 34216 17860 34250 17892
rect 34016 17858 34038 17860
rect 34038 17858 34050 17860
rect 34116 17858 34128 17860
rect 34128 17858 34150 17860
rect 34216 17858 34218 17860
rect 34218 17858 34250 17860
rect 34316 17858 34350 17892
rect 34416 17858 34450 17892
rect 34516 17860 34550 17892
rect 34516 17858 34544 17860
rect 34544 17858 34550 17860
rect 34016 17770 34050 17792
rect 34116 17770 34150 17792
rect 34216 17770 34250 17792
rect 34016 17758 34038 17770
rect 34038 17758 34050 17770
rect 34116 17758 34128 17770
rect 34128 17758 34150 17770
rect 34216 17758 34218 17770
rect 34218 17758 34250 17770
rect 34316 17758 34350 17792
rect 34416 17758 34450 17792
rect 34516 17770 34550 17792
rect 34516 17758 34544 17770
rect 34544 17758 34550 17770
rect 34016 17680 34050 17692
rect 34116 17680 34150 17692
rect 34216 17680 34250 17692
rect 34016 17658 34038 17680
rect 34038 17658 34050 17680
rect 34116 17658 34128 17680
rect 34128 17658 34150 17680
rect 34216 17658 34218 17680
rect 34218 17658 34250 17680
rect 34316 17658 34350 17692
rect 34416 17658 34450 17692
rect 34516 17680 34550 17692
rect 34516 17658 34544 17680
rect 34544 17658 34550 17680
rect 35170 18362 35204 18396
rect 35260 18394 35294 18396
rect 35350 18394 35384 18396
rect 35440 18394 35474 18396
rect 35530 18394 35564 18396
rect 35620 18394 35654 18396
rect 35710 18394 35744 18396
rect 35800 18394 35834 18396
rect 35890 18394 35924 18396
rect 35980 18394 36014 18396
rect 35260 18362 35280 18394
rect 35280 18362 35294 18394
rect 35350 18362 35370 18394
rect 35370 18362 35384 18394
rect 35440 18362 35460 18394
rect 35460 18362 35474 18394
rect 35530 18362 35550 18394
rect 35550 18362 35564 18394
rect 35620 18362 35640 18394
rect 35640 18362 35654 18394
rect 35710 18362 35730 18394
rect 35730 18362 35744 18394
rect 35800 18362 35820 18394
rect 35820 18362 35834 18394
rect 35890 18362 35910 18394
rect 35910 18362 35924 18394
rect 35980 18362 36000 18394
rect 36000 18362 36014 18394
rect 36070 18362 36104 18396
rect 35356 18186 35378 18192
rect 35378 18186 35390 18192
rect 35456 18186 35468 18192
rect 35468 18186 35490 18192
rect 35556 18186 35558 18192
rect 35558 18186 35590 18192
rect 35356 18158 35390 18186
rect 35456 18158 35490 18186
rect 35556 18158 35590 18186
rect 35656 18158 35690 18192
rect 35756 18158 35790 18192
rect 35856 18186 35884 18192
rect 35884 18186 35890 18192
rect 35856 18158 35890 18186
rect 35356 18058 35390 18092
rect 35456 18058 35490 18092
rect 35556 18058 35590 18092
rect 35656 18058 35690 18092
rect 35756 18058 35790 18092
rect 35856 18058 35890 18092
rect 35356 17958 35390 17992
rect 35456 17958 35490 17992
rect 35556 17958 35590 17992
rect 35656 17958 35690 17992
rect 35756 17958 35790 17992
rect 35856 17958 35890 17992
rect 35356 17860 35390 17892
rect 35456 17860 35490 17892
rect 35556 17860 35590 17892
rect 35356 17858 35378 17860
rect 35378 17858 35390 17860
rect 35456 17858 35468 17860
rect 35468 17858 35490 17860
rect 35556 17858 35558 17860
rect 35558 17858 35590 17860
rect 35656 17858 35690 17892
rect 35756 17858 35790 17892
rect 35856 17860 35890 17892
rect 35856 17858 35884 17860
rect 35884 17858 35890 17860
rect 35356 17770 35390 17792
rect 35456 17770 35490 17792
rect 35556 17770 35590 17792
rect 35356 17758 35378 17770
rect 35378 17758 35390 17770
rect 35456 17758 35468 17770
rect 35468 17758 35490 17770
rect 35556 17758 35558 17770
rect 35558 17758 35590 17770
rect 35656 17758 35690 17792
rect 35756 17758 35790 17792
rect 35856 17770 35890 17792
rect 35856 17758 35884 17770
rect 35884 17758 35890 17770
rect 35356 17680 35390 17692
rect 35456 17680 35490 17692
rect 35556 17680 35590 17692
rect 35356 17658 35378 17680
rect 35378 17658 35390 17680
rect 35456 17658 35468 17680
rect 35468 17658 35490 17680
rect 35556 17658 35558 17680
rect 35558 17658 35590 17680
rect 35656 17658 35690 17692
rect 35756 17658 35790 17692
rect 35856 17680 35890 17692
rect 35856 17658 35884 17680
rect 35884 17658 35890 17680
rect 36510 18362 36544 18396
rect 36600 18394 36634 18396
rect 36690 18394 36724 18396
rect 36780 18394 36814 18396
rect 36870 18394 36904 18396
rect 36960 18394 36994 18396
rect 37050 18394 37084 18396
rect 37140 18394 37174 18396
rect 37230 18394 37264 18396
rect 37320 18394 37354 18396
rect 36600 18362 36620 18394
rect 36620 18362 36634 18394
rect 36690 18362 36710 18394
rect 36710 18362 36724 18394
rect 36780 18362 36800 18394
rect 36800 18362 36814 18394
rect 36870 18362 36890 18394
rect 36890 18362 36904 18394
rect 36960 18362 36980 18394
rect 36980 18362 36994 18394
rect 37050 18362 37070 18394
rect 37070 18362 37084 18394
rect 37140 18362 37160 18394
rect 37160 18362 37174 18394
rect 37230 18362 37250 18394
rect 37250 18362 37264 18394
rect 37320 18362 37340 18394
rect 37340 18362 37354 18394
rect 37410 18362 37444 18396
rect 36696 18186 36718 18192
rect 36718 18186 36730 18192
rect 36796 18186 36808 18192
rect 36808 18186 36830 18192
rect 36896 18186 36898 18192
rect 36898 18186 36930 18192
rect 36696 18158 36730 18186
rect 36796 18158 36830 18186
rect 36896 18158 36930 18186
rect 36996 18158 37030 18192
rect 37096 18158 37130 18192
rect 37196 18186 37224 18192
rect 37224 18186 37230 18192
rect 37196 18158 37230 18186
rect 36696 18058 36730 18092
rect 36796 18058 36830 18092
rect 36896 18058 36930 18092
rect 36996 18058 37030 18092
rect 37096 18058 37130 18092
rect 37196 18058 37230 18092
rect 36696 17958 36730 17992
rect 36796 17958 36830 17992
rect 36896 17958 36930 17992
rect 36996 17958 37030 17992
rect 37096 17958 37130 17992
rect 37196 17958 37230 17992
rect 36696 17860 36730 17892
rect 36796 17860 36830 17892
rect 36896 17860 36930 17892
rect 36696 17858 36718 17860
rect 36718 17858 36730 17860
rect 36796 17858 36808 17860
rect 36808 17858 36830 17860
rect 36896 17858 36898 17860
rect 36898 17858 36930 17860
rect 36996 17858 37030 17892
rect 37096 17858 37130 17892
rect 37196 17860 37230 17892
rect 37196 17858 37224 17860
rect 37224 17858 37230 17860
rect 36696 17770 36730 17792
rect 36796 17770 36830 17792
rect 36896 17770 36930 17792
rect 36696 17758 36718 17770
rect 36718 17758 36730 17770
rect 36796 17758 36808 17770
rect 36808 17758 36830 17770
rect 36896 17758 36898 17770
rect 36898 17758 36930 17770
rect 36996 17758 37030 17792
rect 37096 17758 37130 17792
rect 37196 17770 37230 17792
rect 37196 17758 37224 17770
rect 37224 17758 37230 17770
rect 36696 17680 36730 17692
rect 36796 17680 36830 17692
rect 36896 17680 36930 17692
rect 36696 17658 36718 17680
rect 36718 17658 36730 17680
rect 36796 17658 36808 17680
rect 36808 17658 36830 17680
rect 36896 17658 36898 17680
rect 36898 17658 36930 17680
rect 36996 17658 37030 17692
rect 37096 17658 37130 17692
rect 37196 17680 37230 17692
rect 37196 17658 37224 17680
rect 37224 17658 37230 17680
rect 37850 18362 37884 18396
rect 37940 18394 37974 18396
rect 38030 18394 38064 18396
rect 38120 18394 38154 18396
rect 38210 18394 38244 18396
rect 38300 18394 38334 18396
rect 38390 18394 38424 18396
rect 38480 18394 38514 18396
rect 38570 18394 38604 18396
rect 38660 18394 38694 18396
rect 37940 18362 37960 18394
rect 37960 18362 37974 18394
rect 38030 18362 38050 18394
rect 38050 18362 38064 18394
rect 38120 18362 38140 18394
rect 38140 18362 38154 18394
rect 38210 18362 38230 18394
rect 38230 18362 38244 18394
rect 38300 18362 38320 18394
rect 38320 18362 38334 18394
rect 38390 18362 38410 18394
rect 38410 18362 38424 18394
rect 38480 18362 38500 18394
rect 38500 18362 38514 18394
rect 38570 18362 38590 18394
rect 38590 18362 38604 18394
rect 38660 18362 38680 18394
rect 38680 18362 38694 18394
rect 38750 18362 38784 18396
rect 38036 18186 38058 18192
rect 38058 18186 38070 18192
rect 38136 18186 38148 18192
rect 38148 18186 38170 18192
rect 38236 18186 38238 18192
rect 38238 18186 38270 18192
rect 38036 18158 38070 18186
rect 38136 18158 38170 18186
rect 38236 18158 38270 18186
rect 38336 18158 38370 18192
rect 38436 18158 38470 18192
rect 38536 18186 38564 18192
rect 38564 18186 38570 18192
rect 38536 18158 38570 18186
rect 38036 18058 38070 18092
rect 38136 18058 38170 18092
rect 38236 18058 38270 18092
rect 38336 18058 38370 18092
rect 38436 18058 38470 18092
rect 38536 18058 38570 18092
rect 38036 17958 38070 17992
rect 38136 17958 38170 17992
rect 38236 17958 38270 17992
rect 38336 17958 38370 17992
rect 38436 17958 38470 17992
rect 38536 17958 38570 17992
rect 38036 17860 38070 17892
rect 38136 17860 38170 17892
rect 38236 17860 38270 17892
rect 38036 17858 38058 17860
rect 38058 17858 38070 17860
rect 38136 17858 38148 17860
rect 38148 17858 38170 17860
rect 38236 17858 38238 17860
rect 38238 17858 38270 17860
rect 38336 17858 38370 17892
rect 38436 17858 38470 17892
rect 38536 17860 38570 17892
rect 38536 17858 38564 17860
rect 38564 17858 38570 17860
rect 38036 17770 38070 17792
rect 38136 17770 38170 17792
rect 38236 17770 38270 17792
rect 38036 17758 38058 17770
rect 38058 17758 38070 17770
rect 38136 17758 38148 17770
rect 38148 17758 38170 17770
rect 38236 17758 38238 17770
rect 38238 17758 38270 17770
rect 38336 17758 38370 17792
rect 38436 17758 38470 17792
rect 38536 17770 38570 17792
rect 38536 17758 38564 17770
rect 38564 17758 38570 17770
rect 38036 17680 38070 17692
rect 38136 17680 38170 17692
rect 38236 17680 38270 17692
rect 38036 17658 38058 17680
rect 38058 17658 38070 17680
rect 38136 17658 38148 17680
rect 38148 17658 38170 17680
rect 38236 17658 38238 17680
rect 38238 17658 38270 17680
rect 38336 17658 38370 17692
rect 38436 17658 38470 17692
rect 38536 17680 38570 17692
rect 38536 17658 38564 17680
rect 38564 17658 38570 17680
rect 39275 18083 39669 18621
rect 41282 18083 41676 18621
rect 23949 17221 23983 17255
rect 26525 17143 26559 17153
rect 26525 17119 26531 17143
rect 26531 17119 26559 17143
rect 39275 17123 39669 17661
rect 41282 17123 41676 17661
rect 6197 16975 6231 17009
rect 6597 16975 6631 17009
rect 6997 16975 7031 17009
rect 7397 16975 7431 17009
rect 7797 16975 7831 17009
rect 8197 16975 8231 17009
rect 8597 16975 8631 17009
rect 8997 16975 9031 17009
rect 9397 16975 9431 17009
rect 9797 16975 9831 17009
rect 10823 16975 10857 17009
rect 11023 16975 11057 17009
rect 11223 16975 11257 17009
rect 11423 16975 11457 17009
rect 11623 16975 11657 17009
rect 11823 16975 11857 17009
rect 12023 16975 12057 17009
rect 12223 16975 12257 17009
rect 12423 16975 12457 17009
rect 12623 16975 12657 17009
rect 12823 16975 12857 17009
rect 13567 16975 13601 17009
rect 13767 16975 13801 17009
rect 13967 16975 14001 17009
rect 14167 16975 14201 17009
rect 14367 16975 14401 17009
rect 14567 16975 14601 17009
rect 14767 16975 14801 17009
rect 14967 16975 15001 17009
rect 15167 16975 15201 17009
rect 15367 16975 15401 17009
rect 15567 16975 15601 17009
rect 16293 16975 16327 17009
rect 16693 16975 16727 17009
rect 17093 16975 17127 17009
rect 17493 16975 17527 17009
rect 17893 16975 17927 17009
rect 18293 16975 18327 17009
rect 18693 16975 18727 17009
rect 19093 16975 19127 17009
rect 19493 16975 19527 17009
rect 19893 16975 19927 17009
rect 20293 16975 20327 17009
rect 20693 16975 20727 17009
rect 21093 16975 21127 17009
rect 21493 16975 21527 17009
rect 21893 16975 21927 17009
rect 22293 16975 22327 17009
rect 22693 16975 22727 17009
rect 23093 16975 23127 17009
rect 24131 16975 24165 17009
rect 24531 16975 24565 17009
rect 24931 16975 24965 17009
rect 25331 16975 25365 17009
rect 25731 16975 25765 17009
rect 26131 16975 26165 17009
rect 26531 16975 26565 17009
rect 28443 16975 28477 17009
rect 28643 16975 28677 17009
rect 28843 16975 28877 17009
rect 29043 16975 29077 17009
rect 29243 16975 29277 17009
rect 29443 16975 29477 17009
rect 29643 16975 29677 17009
rect 29843 16975 29877 17009
rect 30043 16975 30077 17009
rect 30243 16975 30277 17009
rect 30443 16975 30477 17009
rect 30643 16975 30677 17009
rect 30843 16975 30877 17009
rect 31043 16975 31077 17009
rect 31243 16975 31277 17009
rect 31443 16975 31477 17009
rect 31643 16975 31677 17009
rect 31843 16975 31877 17009
rect 32043 16975 32077 17009
rect 32243 16975 32277 17009
rect 32443 16975 32477 17009
rect 32643 16975 32677 17009
rect 32843 16975 32877 17009
rect 33043 16975 33077 17009
rect 33243 16975 33277 17009
rect 33443 16975 33477 17009
rect 33643 16975 33677 17009
rect 33843 16975 33877 17009
rect 34043 16975 34077 17009
rect 34243 16975 34277 17009
rect 34443 16975 34477 17009
rect 34643 16975 34677 17009
rect 34843 16975 34877 17009
rect 35043 16975 35077 17009
rect 35243 16975 35277 17009
rect 35443 16975 35477 17009
rect 35643 16975 35677 17009
rect 35843 16975 35877 17009
rect 36043 16975 36077 17009
rect 36243 16975 36277 17009
rect 36443 16975 36477 17009
rect 36643 16975 36677 17009
rect 36843 16975 36877 17009
rect 37043 16975 37077 17009
rect 37243 16975 37277 17009
rect 37443 16975 37477 17009
rect 37643 16975 37677 17009
rect 37843 16975 37877 17009
rect 38043 16975 38077 17009
rect 38243 16975 38277 17009
rect 38443 16975 38477 17009
rect 38643 16975 38677 17009
rect 38843 16975 38877 17009
rect 39439 16975 39473 17009
rect 39639 16975 39673 17009
rect 39839 16975 39873 17009
rect 40039 16975 40073 17009
rect 40239 16975 40273 17009
rect 40439 16975 40473 17009
rect 40639 16975 40673 17009
rect 40839 16975 40873 17009
rect 41039 16975 41073 17009
rect 41239 16975 41273 17009
rect 41439 16975 41473 17009
rect 8079 15095 8113 15129
rect 8279 15095 8313 15129
rect 8479 15095 8513 15129
rect 8679 15095 8713 15129
rect 8879 15095 8913 15129
rect 9079 15095 9113 15129
rect 9279 15095 9313 15129
rect 9479 15095 9513 15129
rect 9679 15095 9713 15129
rect 9879 15095 9913 15129
rect 10079 15095 10113 15129
rect 10823 15095 10857 15129
rect 11023 15095 11057 15129
rect 11223 15095 11257 15129
rect 11423 15095 11457 15129
rect 11623 15095 11657 15129
rect 11823 15095 11857 15129
rect 12023 15095 12057 15129
rect 12223 15095 12257 15129
rect 12423 15095 12457 15129
rect 12623 15095 12657 15129
rect 12823 15095 12857 15129
rect 13567 15095 13601 15129
rect 13767 15095 13801 15129
rect 13967 15095 14001 15129
rect 14167 15095 14201 15129
rect 14367 15095 14401 15129
rect 14567 15095 14601 15129
rect 14767 15095 14801 15129
rect 14967 15095 15001 15129
rect 15167 15095 15201 15129
rect 15367 15095 15401 15129
rect 15567 15095 15601 15129
rect 16293 15095 16327 15129
rect 16693 15095 16727 15129
rect 17093 15095 17127 15129
rect 17493 15095 17527 15129
rect 17893 15095 17927 15129
rect 18293 15095 18327 15129
rect 18693 15095 18727 15129
rect 19093 15095 19127 15129
rect 19493 15095 19527 15129
rect 19893 15095 19927 15129
rect 20293 15095 20327 15129
rect 20693 15095 20727 15129
rect 21093 15095 21127 15129
rect 21493 15095 21527 15129
rect 21893 15095 21927 15129
rect 22293 15095 22327 15129
rect 22693 15095 22727 15129
rect 23093 15095 23127 15129
rect 23759 15095 23793 15129
rect 23959 15095 23993 15129
rect 24159 15095 24193 15129
rect 24359 15095 24393 15129
rect 24559 15095 24593 15129
rect 24759 15095 24793 15129
rect 24959 15095 24993 15129
rect 25159 15095 25193 15129
rect 25359 15095 25393 15129
rect 25559 15095 25593 15129
rect 25759 15095 25793 15129
rect 28443 15095 28477 15129
rect 28643 15095 28677 15129
rect 28843 15095 28877 15129
rect 29043 15095 29077 15129
rect 29243 15095 29277 15129
rect 29443 15095 29477 15129
rect 29643 15095 29677 15129
rect 29843 15095 29877 15129
rect 30043 15095 30077 15129
rect 30243 15095 30277 15129
rect 30443 15095 30477 15129
rect 30643 15095 30677 15129
rect 30843 15095 30877 15129
rect 31043 15095 31077 15129
rect 31243 15095 31277 15129
rect 31443 15095 31477 15129
rect 31643 15095 31677 15129
rect 31843 15095 31877 15129
rect 32043 15095 32077 15129
rect 32243 15095 32277 15129
rect 32443 15095 32477 15129
rect 32643 15095 32677 15129
rect 32843 15095 32877 15129
rect 33043 15095 33077 15129
rect 33243 15095 33277 15129
rect 33443 15095 33477 15129
rect 33643 15095 33677 15129
rect 33843 15095 33877 15129
rect 34043 15095 34077 15129
rect 34243 15095 34277 15129
rect 34443 15095 34477 15129
rect 34643 15095 34677 15129
rect 34843 15095 34877 15129
rect 35043 15095 35077 15129
rect 35243 15095 35277 15129
rect 35443 15095 35477 15129
rect 35643 15095 35677 15129
rect 35843 15095 35877 15129
rect 36043 15095 36077 15129
rect 36243 15095 36277 15129
rect 36443 15095 36477 15129
rect 36643 15095 36677 15129
rect 36843 15095 36877 15129
rect 37043 15095 37077 15129
rect 37243 15095 37277 15129
rect 37443 15095 37477 15129
rect 37643 15095 37677 15129
rect 37843 15095 37877 15129
rect 38043 15095 38077 15129
rect 38243 15095 38277 15129
rect 38443 15095 38477 15129
rect 38643 15095 38677 15129
rect 38843 15095 38877 15129
rect 39439 15095 39473 15129
rect 39639 15095 39673 15129
rect 39839 15095 39873 15129
rect 40039 15095 40073 15129
rect 40239 15095 40273 15129
rect 40439 15095 40473 15129
rect 40639 15095 40673 15129
rect 40839 15095 40873 15129
rect 41039 15095 41073 15129
rect 41239 15095 41273 15129
rect 41439 15095 41473 15129
rect 7915 14323 8309 14861
rect 9922 14323 10316 14861
rect 10659 14323 11053 14861
rect 12666 14323 13060 14861
rect 13403 14323 13797 14861
rect 15410 14323 15804 14861
rect 23595 14323 23989 14861
rect 25602 14323 25996 14861
rect 7915 13363 8309 13901
rect 9922 13363 10316 13901
rect 10659 13363 11053 13901
rect 12666 13363 13060 13901
rect 13403 13363 13797 13901
rect 15410 13363 15804 13901
rect 23595 13363 23989 13901
rect 25602 13363 25996 13901
rect 28306 14762 28340 14796
rect 28396 14781 28430 14796
rect 28486 14781 28520 14796
rect 28576 14781 28610 14796
rect 28666 14781 28700 14796
rect 28756 14781 28790 14796
rect 28846 14781 28880 14796
rect 28936 14781 28970 14796
rect 29026 14781 29060 14796
rect 29116 14781 29150 14796
rect 29206 14781 29240 14796
rect 29296 14781 29330 14796
rect 29386 14781 29420 14796
rect 28396 14762 28416 14781
rect 28416 14762 28430 14781
rect 28486 14762 28506 14781
rect 28506 14762 28520 14781
rect 28576 14762 28596 14781
rect 28596 14762 28610 14781
rect 28666 14762 28686 14781
rect 28686 14762 28700 14781
rect 28756 14762 28776 14781
rect 28776 14762 28790 14781
rect 28846 14762 28866 14781
rect 28866 14762 28880 14781
rect 28936 14762 28956 14781
rect 28956 14762 28970 14781
rect 29026 14762 29046 14781
rect 29046 14762 29060 14781
rect 29116 14762 29136 14781
rect 29136 14762 29150 14781
rect 29206 14762 29226 14781
rect 29226 14762 29240 14781
rect 29296 14762 29316 14781
rect 29316 14762 29330 14781
rect 29386 14762 29406 14781
rect 29406 14762 29420 14781
rect 29476 14762 29510 14796
rect 29646 14762 29680 14796
rect 29736 14781 29770 14796
rect 29826 14781 29860 14796
rect 29916 14781 29950 14796
rect 30006 14781 30040 14796
rect 30096 14781 30130 14796
rect 30186 14781 30220 14796
rect 30276 14781 30310 14796
rect 30366 14781 30400 14796
rect 30456 14781 30490 14796
rect 30546 14781 30580 14796
rect 30636 14781 30670 14796
rect 30726 14781 30760 14796
rect 29736 14762 29756 14781
rect 29756 14762 29770 14781
rect 29826 14762 29846 14781
rect 29846 14762 29860 14781
rect 29916 14762 29936 14781
rect 29936 14762 29950 14781
rect 30006 14762 30026 14781
rect 30026 14762 30040 14781
rect 30096 14762 30116 14781
rect 30116 14762 30130 14781
rect 30186 14762 30206 14781
rect 30206 14762 30220 14781
rect 30276 14762 30296 14781
rect 30296 14762 30310 14781
rect 30366 14762 30386 14781
rect 30386 14762 30400 14781
rect 30456 14762 30476 14781
rect 30476 14762 30490 14781
rect 30546 14762 30566 14781
rect 30566 14762 30580 14781
rect 30636 14762 30656 14781
rect 30656 14762 30670 14781
rect 30726 14762 30746 14781
rect 30746 14762 30760 14781
rect 30816 14762 30850 14796
rect 30986 14762 31020 14796
rect 31076 14781 31110 14796
rect 31166 14781 31200 14796
rect 31256 14781 31290 14796
rect 31346 14781 31380 14796
rect 31436 14781 31470 14796
rect 31526 14781 31560 14796
rect 31616 14781 31650 14796
rect 31706 14781 31740 14796
rect 31796 14781 31830 14796
rect 31886 14781 31920 14796
rect 31976 14781 32010 14796
rect 32066 14781 32100 14796
rect 31076 14762 31096 14781
rect 31096 14762 31110 14781
rect 31166 14762 31186 14781
rect 31186 14762 31200 14781
rect 31256 14762 31276 14781
rect 31276 14762 31290 14781
rect 31346 14762 31366 14781
rect 31366 14762 31380 14781
rect 31436 14762 31456 14781
rect 31456 14762 31470 14781
rect 31526 14762 31546 14781
rect 31546 14762 31560 14781
rect 31616 14762 31636 14781
rect 31636 14762 31650 14781
rect 31706 14762 31726 14781
rect 31726 14762 31740 14781
rect 31796 14762 31816 14781
rect 31816 14762 31830 14781
rect 31886 14762 31906 14781
rect 31906 14762 31920 14781
rect 31976 14762 31996 14781
rect 31996 14762 32010 14781
rect 32066 14762 32086 14781
rect 32086 14762 32100 14781
rect 32156 14762 32190 14796
rect 32326 14762 32360 14796
rect 32416 14781 32450 14796
rect 32506 14781 32540 14796
rect 32596 14781 32630 14796
rect 32686 14781 32720 14796
rect 32776 14781 32810 14796
rect 32866 14781 32900 14796
rect 32956 14781 32990 14796
rect 33046 14781 33080 14796
rect 33136 14781 33170 14796
rect 33226 14781 33260 14796
rect 33316 14781 33350 14796
rect 33406 14781 33440 14796
rect 32416 14762 32436 14781
rect 32436 14762 32450 14781
rect 32506 14762 32526 14781
rect 32526 14762 32540 14781
rect 32596 14762 32616 14781
rect 32616 14762 32630 14781
rect 32686 14762 32706 14781
rect 32706 14762 32720 14781
rect 32776 14762 32796 14781
rect 32796 14762 32810 14781
rect 32866 14762 32886 14781
rect 32886 14762 32900 14781
rect 32956 14762 32976 14781
rect 32976 14762 32990 14781
rect 33046 14762 33066 14781
rect 33066 14762 33080 14781
rect 33136 14762 33156 14781
rect 33156 14762 33170 14781
rect 33226 14762 33246 14781
rect 33246 14762 33260 14781
rect 33316 14762 33336 14781
rect 33336 14762 33350 14781
rect 33406 14762 33426 14781
rect 33426 14762 33440 14781
rect 33496 14762 33530 14796
rect 33666 14762 33700 14796
rect 33756 14781 33790 14796
rect 33846 14781 33880 14796
rect 33936 14781 33970 14796
rect 34026 14781 34060 14796
rect 34116 14781 34150 14796
rect 34206 14781 34240 14796
rect 34296 14781 34330 14796
rect 34386 14781 34420 14796
rect 34476 14781 34510 14796
rect 34566 14781 34600 14796
rect 34656 14781 34690 14796
rect 34746 14781 34780 14796
rect 33756 14762 33776 14781
rect 33776 14762 33790 14781
rect 33846 14762 33866 14781
rect 33866 14762 33880 14781
rect 33936 14762 33956 14781
rect 33956 14762 33970 14781
rect 34026 14762 34046 14781
rect 34046 14762 34060 14781
rect 34116 14762 34136 14781
rect 34136 14762 34150 14781
rect 34206 14762 34226 14781
rect 34226 14762 34240 14781
rect 34296 14762 34316 14781
rect 34316 14762 34330 14781
rect 34386 14762 34406 14781
rect 34406 14762 34420 14781
rect 34476 14762 34496 14781
rect 34496 14762 34510 14781
rect 34566 14762 34586 14781
rect 34586 14762 34600 14781
rect 34656 14762 34676 14781
rect 34676 14762 34690 14781
rect 34746 14762 34766 14781
rect 34766 14762 34780 14781
rect 34836 14762 34870 14796
rect 35006 14762 35040 14796
rect 35096 14781 35130 14796
rect 35186 14781 35220 14796
rect 35276 14781 35310 14796
rect 35366 14781 35400 14796
rect 35456 14781 35490 14796
rect 35546 14781 35580 14796
rect 35636 14781 35670 14796
rect 35726 14781 35760 14796
rect 35816 14781 35850 14796
rect 35906 14781 35940 14796
rect 35996 14781 36030 14796
rect 36086 14781 36120 14796
rect 35096 14762 35116 14781
rect 35116 14762 35130 14781
rect 35186 14762 35206 14781
rect 35206 14762 35220 14781
rect 35276 14762 35296 14781
rect 35296 14762 35310 14781
rect 35366 14762 35386 14781
rect 35386 14762 35400 14781
rect 35456 14762 35476 14781
rect 35476 14762 35490 14781
rect 35546 14762 35566 14781
rect 35566 14762 35580 14781
rect 35636 14762 35656 14781
rect 35656 14762 35670 14781
rect 35726 14762 35746 14781
rect 35746 14762 35760 14781
rect 35816 14762 35836 14781
rect 35836 14762 35850 14781
rect 35906 14762 35926 14781
rect 35926 14762 35940 14781
rect 35996 14762 36016 14781
rect 36016 14762 36030 14781
rect 36086 14762 36106 14781
rect 36106 14762 36120 14781
rect 36176 14762 36210 14796
rect 36346 14762 36380 14796
rect 36436 14781 36470 14796
rect 36526 14781 36560 14796
rect 36616 14781 36650 14796
rect 36706 14781 36740 14796
rect 36796 14781 36830 14796
rect 36886 14781 36920 14796
rect 36976 14781 37010 14796
rect 37066 14781 37100 14796
rect 37156 14781 37190 14796
rect 37246 14781 37280 14796
rect 37336 14781 37370 14796
rect 37426 14781 37460 14796
rect 36436 14762 36456 14781
rect 36456 14762 36470 14781
rect 36526 14762 36546 14781
rect 36546 14762 36560 14781
rect 36616 14762 36636 14781
rect 36636 14762 36650 14781
rect 36706 14762 36726 14781
rect 36726 14762 36740 14781
rect 36796 14762 36816 14781
rect 36816 14762 36830 14781
rect 36886 14762 36906 14781
rect 36906 14762 36920 14781
rect 36976 14762 36996 14781
rect 36996 14762 37010 14781
rect 37066 14762 37086 14781
rect 37086 14762 37100 14781
rect 37156 14762 37176 14781
rect 37176 14762 37190 14781
rect 37246 14762 37266 14781
rect 37266 14762 37280 14781
rect 37336 14762 37356 14781
rect 37356 14762 37370 14781
rect 37426 14762 37446 14781
rect 37446 14762 37460 14781
rect 37516 14762 37550 14796
rect 37686 14762 37720 14796
rect 37776 14781 37810 14796
rect 37866 14781 37900 14796
rect 37956 14781 37990 14796
rect 38046 14781 38080 14796
rect 38136 14781 38170 14796
rect 38226 14781 38260 14796
rect 38316 14781 38350 14796
rect 38406 14781 38440 14796
rect 38496 14781 38530 14796
rect 38586 14781 38620 14796
rect 38676 14781 38710 14796
rect 38766 14781 38800 14796
rect 37776 14762 37796 14781
rect 37796 14762 37810 14781
rect 37866 14762 37886 14781
rect 37886 14762 37900 14781
rect 37956 14762 37976 14781
rect 37976 14762 37990 14781
rect 38046 14762 38066 14781
rect 38066 14762 38080 14781
rect 38136 14762 38156 14781
rect 38156 14762 38170 14781
rect 38226 14762 38246 14781
rect 38246 14762 38260 14781
rect 38316 14762 38336 14781
rect 38336 14762 38350 14781
rect 38406 14762 38426 14781
rect 38426 14762 38440 14781
rect 38496 14762 38516 14781
rect 38516 14762 38530 14781
rect 38586 14762 38606 14781
rect 38606 14762 38620 14781
rect 38676 14762 38696 14781
rect 38696 14762 38710 14781
rect 38766 14762 38786 14781
rect 38786 14762 38800 14781
rect 38856 14762 38890 14796
rect 28470 14602 28504 14636
rect 28560 14634 28594 14636
rect 28650 14634 28684 14636
rect 28740 14634 28774 14636
rect 28830 14634 28864 14636
rect 28920 14634 28954 14636
rect 29010 14634 29044 14636
rect 29100 14634 29134 14636
rect 29190 14634 29224 14636
rect 29280 14634 29314 14636
rect 28560 14602 28580 14634
rect 28580 14602 28594 14634
rect 28650 14602 28670 14634
rect 28670 14602 28684 14634
rect 28740 14602 28760 14634
rect 28760 14602 28774 14634
rect 28830 14602 28850 14634
rect 28850 14602 28864 14634
rect 28920 14602 28940 14634
rect 28940 14602 28954 14634
rect 29010 14602 29030 14634
rect 29030 14602 29044 14634
rect 29100 14602 29120 14634
rect 29120 14602 29134 14634
rect 29190 14602 29210 14634
rect 29210 14602 29224 14634
rect 29280 14602 29300 14634
rect 29300 14602 29314 14634
rect 29370 14602 29404 14636
rect 28656 14426 28678 14432
rect 28678 14426 28690 14432
rect 28756 14426 28768 14432
rect 28768 14426 28790 14432
rect 28856 14426 28858 14432
rect 28858 14426 28890 14432
rect 28656 14398 28690 14426
rect 28756 14398 28790 14426
rect 28856 14398 28890 14426
rect 28956 14398 28990 14432
rect 29056 14398 29090 14432
rect 29156 14426 29184 14432
rect 29184 14426 29190 14432
rect 29156 14398 29190 14426
rect 28656 14298 28690 14332
rect 28756 14298 28790 14332
rect 28856 14298 28890 14332
rect 28956 14298 28990 14332
rect 29056 14298 29090 14332
rect 29156 14298 29190 14332
rect 28656 14198 28690 14232
rect 28756 14198 28790 14232
rect 28856 14198 28890 14232
rect 28956 14198 28990 14232
rect 29056 14198 29090 14232
rect 29156 14198 29190 14232
rect 28656 14100 28690 14132
rect 28756 14100 28790 14132
rect 28856 14100 28890 14132
rect 28656 14098 28678 14100
rect 28678 14098 28690 14100
rect 28756 14098 28768 14100
rect 28768 14098 28790 14100
rect 28856 14098 28858 14100
rect 28858 14098 28890 14100
rect 28956 14098 28990 14132
rect 29056 14098 29090 14132
rect 29156 14100 29190 14132
rect 29156 14098 29184 14100
rect 29184 14098 29190 14100
rect 28656 14010 28690 14032
rect 28756 14010 28790 14032
rect 28856 14010 28890 14032
rect 28656 13998 28678 14010
rect 28678 13998 28690 14010
rect 28756 13998 28768 14010
rect 28768 13998 28790 14010
rect 28856 13998 28858 14010
rect 28858 13998 28890 14010
rect 28956 13998 28990 14032
rect 29056 13998 29090 14032
rect 29156 14010 29190 14032
rect 29156 13998 29184 14010
rect 29184 13998 29190 14010
rect 28656 13920 28690 13932
rect 28756 13920 28790 13932
rect 28856 13920 28890 13932
rect 28656 13898 28678 13920
rect 28678 13898 28690 13920
rect 28756 13898 28768 13920
rect 28768 13898 28790 13920
rect 28856 13898 28858 13920
rect 28858 13898 28890 13920
rect 28956 13898 28990 13932
rect 29056 13898 29090 13932
rect 29156 13920 29190 13932
rect 29156 13898 29184 13920
rect 29184 13898 29190 13920
rect 29810 14602 29844 14636
rect 29900 14634 29934 14636
rect 29990 14634 30024 14636
rect 30080 14634 30114 14636
rect 30170 14634 30204 14636
rect 30260 14634 30294 14636
rect 30350 14634 30384 14636
rect 30440 14634 30474 14636
rect 30530 14634 30564 14636
rect 30620 14634 30654 14636
rect 29900 14602 29920 14634
rect 29920 14602 29934 14634
rect 29990 14602 30010 14634
rect 30010 14602 30024 14634
rect 30080 14602 30100 14634
rect 30100 14602 30114 14634
rect 30170 14602 30190 14634
rect 30190 14602 30204 14634
rect 30260 14602 30280 14634
rect 30280 14602 30294 14634
rect 30350 14602 30370 14634
rect 30370 14602 30384 14634
rect 30440 14602 30460 14634
rect 30460 14602 30474 14634
rect 30530 14602 30550 14634
rect 30550 14602 30564 14634
rect 30620 14602 30640 14634
rect 30640 14602 30654 14634
rect 30710 14602 30744 14636
rect 29996 14426 30018 14432
rect 30018 14426 30030 14432
rect 30096 14426 30108 14432
rect 30108 14426 30130 14432
rect 30196 14426 30198 14432
rect 30198 14426 30230 14432
rect 29996 14398 30030 14426
rect 30096 14398 30130 14426
rect 30196 14398 30230 14426
rect 30296 14398 30330 14432
rect 30396 14398 30430 14432
rect 30496 14426 30524 14432
rect 30524 14426 30530 14432
rect 30496 14398 30530 14426
rect 29996 14298 30030 14332
rect 30096 14298 30130 14332
rect 30196 14298 30230 14332
rect 30296 14298 30330 14332
rect 30396 14298 30430 14332
rect 30496 14298 30530 14332
rect 29996 14198 30030 14232
rect 30096 14198 30130 14232
rect 30196 14198 30230 14232
rect 30296 14198 30330 14232
rect 30396 14198 30430 14232
rect 30496 14198 30530 14232
rect 29996 14100 30030 14132
rect 30096 14100 30130 14132
rect 30196 14100 30230 14132
rect 29996 14098 30018 14100
rect 30018 14098 30030 14100
rect 30096 14098 30108 14100
rect 30108 14098 30130 14100
rect 30196 14098 30198 14100
rect 30198 14098 30230 14100
rect 30296 14098 30330 14132
rect 30396 14098 30430 14132
rect 30496 14100 30530 14132
rect 30496 14098 30524 14100
rect 30524 14098 30530 14100
rect 29996 14010 30030 14032
rect 30096 14010 30130 14032
rect 30196 14010 30230 14032
rect 29996 13998 30018 14010
rect 30018 13998 30030 14010
rect 30096 13998 30108 14010
rect 30108 13998 30130 14010
rect 30196 13998 30198 14010
rect 30198 13998 30230 14010
rect 30296 13998 30330 14032
rect 30396 13998 30430 14032
rect 30496 14010 30530 14032
rect 30496 13998 30524 14010
rect 30524 13998 30530 14010
rect 29996 13920 30030 13932
rect 30096 13920 30130 13932
rect 30196 13920 30230 13932
rect 29996 13898 30018 13920
rect 30018 13898 30030 13920
rect 30096 13898 30108 13920
rect 30108 13898 30130 13920
rect 30196 13898 30198 13920
rect 30198 13898 30230 13920
rect 30296 13898 30330 13932
rect 30396 13898 30430 13932
rect 30496 13920 30530 13932
rect 30496 13898 30524 13920
rect 30524 13898 30530 13920
rect 31150 14602 31184 14636
rect 31240 14634 31274 14636
rect 31330 14634 31364 14636
rect 31420 14634 31454 14636
rect 31510 14634 31544 14636
rect 31600 14634 31634 14636
rect 31690 14634 31724 14636
rect 31780 14634 31814 14636
rect 31870 14634 31904 14636
rect 31960 14634 31994 14636
rect 31240 14602 31260 14634
rect 31260 14602 31274 14634
rect 31330 14602 31350 14634
rect 31350 14602 31364 14634
rect 31420 14602 31440 14634
rect 31440 14602 31454 14634
rect 31510 14602 31530 14634
rect 31530 14602 31544 14634
rect 31600 14602 31620 14634
rect 31620 14602 31634 14634
rect 31690 14602 31710 14634
rect 31710 14602 31724 14634
rect 31780 14602 31800 14634
rect 31800 14602 31814 14634
rect 31870 14602 31890 14634
rect 31890 14602 31904 14634
rect 31960 14602 31980 14634
rect 31980 14602 31994 14634
rect 32050 14602 32084 14636
rect 31336 14426 31358 14432
rect 31358 14426 31370 14432
rect 31436 14426 31448 14432
rect 31448 14426 31470 14432
rect 31536 14426 31538 14432
rect 31538 14426 31570 14432
rect 31336 14398 31370 14426
rect 31436 14398 31470 14426
rect 31536 14398 31570 14426
rect 31636 14398 31670 14432
rect 31736 14398 31770 14432
rect 31836 14426 31864 14432
rect 31864 14426 31870 14432
rect 31836 14398 31870 14426
rect 31336 14298 31370 14332
rect 31436 14298 31470 14332
rect 31536 14298 31570 14332
rect 31636 14298 31670 14332
rect 31736 14298 31770 14332
rect 31836 14298 31870 14332
rect 31336 14198 31370 14232
rect 31436 14198 31470 14232
rect 31536 14198 31570 14232
rect 31636 14198 31670 14232
rect 31736 14198 31770 14232
rect 31836 14198 31870 14232
rect 31336 14100 31370 14132
rect 31436 14100 31470 14132
rect 31536 14100 31570 14132
rect 31336 14098 31358 14100
rect 31358 14098 31370 14100
rect 31436 14098 31448 14100
rect 31448 14098 31470 14100
rect 31536 14098 31538 14100
rect 31538 14098 31570 14100
rect 31636 14098 31670 14132
rect 31736 14098 31770 14132
rect 31836 14100 31870 14132
rect 31836 14098 31864 14100
rect 31864 14098 31870 14100
rect 31336 14010 31370 14032
rect 31436 14010 31470 14032
rect 31536 14010 31570 14032
rect 31336 13998 31358 14010
rect 31358 13998 31370 14010
rect 31436 13998 31448 14010
rect 31448 13998 31470 14010
rect 31536 13998 31538 14010
rect 31538 13998 31570 14010
rect 31636 13998 31670 14032
rect 31736 13998 31770 14032
rect 31836 14010 31870 14032
rect 31836 13998 31864 14010
rect 31864 13998 31870 14010
rect 31336 13920 31370 13932
rect 31436 13920 31470 13932
rect 31536 13920 31570 13932
rect 31336 13898 31358 13920
rect 31358 13898 31370 13920
rect 31436 13898 31448 13920
rect 31448 13898 31470 13920
rect 31536 13898 31538 13920
rect 31538 13898 31570 13920
rect 31636 13898 31670 13932
rect 31736 13898 31770 13932
rect 31836 13920 31870 13932
rect 31836 13898 31864 13920
rect 31864 13898 31870 13920
rect 32490 14602 32524 14636
rect 32580 14634 32614 14636
rect 32670 14634 32704 14636
rect 32760 14634 32794 14636
rect 32850 14634 32884 14636
rect 32940 14634 32974 14636
rect 33030 14634 33064 14636
rect 33120 14634 33154 14636
rect 33210 14634 33244 14636
rect 33300 14634 33334 14636
rect 32580 14602 32600 14634
rect 32600 14602 32614 14634
rect 32670 14602 32690 14634
rect 32690 14602 32704 14634
rect 32760 14602 32780 14634
rect 32780 14602 32794 14634
rect 32850 14602 32870 14634
rect 32870 14602 32884 14634
rect 32940 14602 32960 14634
rect 32960 14602 32974 14634
rect 33030 14602 33050 14634
rect 33050 14602 33064 14634
rect 33120 14602 33140 14634
rect 33140 14602 33154 14634
rect 33210 14602 33230 14634
rect 33230 14602 33244 14634
rect 33300 14602 33320 14634
rect 33320 14602 33334 14634
rect 33390 14602 33424 14636
rect 32676 14426 32698 14432
rect 32698 14426 32710 14432
rect 32776 14426 32788 14432
rect 32788 14426 32810 14432
rect 32876 14426 32878 14432
rect 32878 14426 32910 14432
rect 32676 14398 32710 14426
rect 32776 14398 32810 14426
rect 32876 14398 32910 14426
rect 32976 14398 33010 14432
rect 33076 14398 33110 14432
rect 33176 14426 33204 14432
rect 33204 14426 33210 14432
rect 33176 14398 33210 14426
rect 32676 14298 32710 14332
rect 32776 14298 32810 14332
rect 32876 14298 32910 14332
rect 32976 14298 33010 14332
rect 33076 14298 33110 14332
rect 33176 14298 33210 14332
rect 32676 14198 32710 14232
rect 32776 14198 32810 14232
rect 32876 14198 32910 14232
rect 32976 14198 33010 14232
rect 33076 14198 33110 14232
rect 33176 14198 33210 14232
rect 32676 14100 32710 14132
rect 32776 14100 32810 14132
rect 32876 14100 32910 14132
rect 32676 14098 32698 14100
rect 32698 14098 32710 14100
rect 32776 14098 32788 14100
rect 32788 14098 32810 14100
rect 32876 14098 32878 14100
rect 32878 14098 32910 14100
rect 32976 14098 33010 14132
rect 33076 14098 33110 14132
rect 33176 14100 33210 14132
rect 33176 14098 33204 14100
rect 33204 14098 33210 14100
rect 32676 14010 32710 14032
rect 32776 14010 32810 14032
rect 32876 14010 32910 14032
rect 32676 13998 32698 14010
rect 32698 13998 32710 14010
rect 32776 13998 32788 14010
rect 32788 13998 32810 14010
rect 32876 13998 32878 14010
rect 32878 13998 32910 14010
rect 32976 13998 33010 14032
rect 33076 13998 33110 14032
rect 33176 14010 33210 14032
rect 33176 13998 33204 14010
rect 33204 13998 33210 14010
rect 32676 13920 32710 13932
rect 32776 13920 32810 13932
rect 32876 13920 32910 13932
rect 32676 13898 32698 13920
rect 32698 13898 32710 13920
rect 32776 13898 32788 13920
rect 32788 13898 32810 13920
rect 32876 13898 32878 13920
rect 32878 13898 32910 13920
rect 32976 13898 33010 13932
rect 33076 13898 33110 13932
rect 33176 13920 33210 13932
rect 33176 13898 33204 13920
rect 33204 13898 33210 13920
rect 33830 14602 33864 14636
rect 33920 14634 33954 14636
rect 34010 14634 34044 14636
rect 34100 14634 34134 14636
rect 34190 14634 34224 14636
rect 34280 14634 34314 14636
rect 34370 14634 34404 14636
rect 34460 14634 34494 14636
rect 34550 14634 34584 14636
rect 34640 14634 34674 14636
rect 33920 14602 33940 14634
rect 33940 14602 33954 14634
rect 34010 14602 34030 14634
rect 34030 14602 34044 14634
rect 34100 14602 34120 14634
rect 34120 14602 34134 14634
rect 34190 14602 34210 14634
rect 34210 14602 34224 14634
rect 34280 14602 34300 14634
rect 34300 14602 34314 14634
rect 34370 14602 34390 14634
rect 34390 14602 34404 14634
rect 34460 14602 34480 14634
rect 34480 14602 34494 14634
rect 34550 14602 34570 14634
rect 34570 14602 34584 14634
rect 34640 14602 34660 14634
rect 34660 14602 34674 14634
rect 34730 14602 34764 14636
rect 34016 14426 34038 14432
rect 34038 14426 34050 14432
rect 34116 14426 34128 14432
rect 34128 14426 34150 14432
rect 34216 14426 34218 14432
rect 34218 14426 34250 14432
rect 34016 14398 34050 14426
rect 34116 14398 34150 14426
rect 34216 14398 34250 14426
rect 34316 14398 34350 14432
rect 34416 14398 34450 14432
rect 34516 14426 34544 14432
rect 34544 14426 34550 14432
rect 34516 14398 34550 14426
rect 34016 14298 34050 14332
rect 34116 14298 34150 14332
rect 34216 14298 34250 14332
rect 34316 14298 34350 14332
rect 34416 14298 34450 14332
rect 34516 14298 34550 14332
rect 34016 14198 34050 14232
rect 34116 14198 34150 14232
rect 34216 14198 34250 14232
rect 34316 14198 34350 14232
rect 34416 14198 34450 14232
rect 34516 14198 34550 14232
rect 34016 14100 34050 14132
rect 34116 14100 34150 14132
rect 34216 14100 34250 14132
rect 34016 14098 34038 14100
rect 34038 14098 34050 14100
rect 34116 14098 34128 14100
rect 34128 14098 34150 14100
rect 34216 14098 34218 14100
rect 34218 14098 34250 14100
rect 34316 14098 34350 14132
rect 34416 14098 34450 14132
rect 34516 14100 34550 14132
rect 34516 14098 34544 14100
rect 34544 14098 34550 14100
rect 34016 14010 34050 14032
rect 34116 14010 34150 14032
rect 34216 14010 34250 14032
rect 34016 13998 34038 14010
rect 34038 13998 34050 14010
rect 34116 13998 34128 14010
rect 34128 13998 34150 14010
rect 34216 13998 34218 14010
rect 34218 13998 34250 14010
rect 34316 13998 34350 14032
rect 34416 13998 34450 14032
rect 34516 14010 34550 14032
rect 34516 13998 34544 14010
rect 34544 13998 34550 14010
rect 34016 13920 34050 13932
rect 34116 13920 34150 13932
rect 34216 13920 34250 13932
rect 34016 13898 34038 13920
rect 34038 13898 34050 13920
rect 34116 13898 34128 13920
rect 34128 13898 34150 13920
rect 34216 13898 34218 13920
rect 34218 13898 34250 13920
rect 34316 13898 34350 13932
rect 34416 13898 34450 13932
rect 34516 13920 34550 13932
rect 34516 13898 34544 13920
rect 34544 13898 34550 13920
rect 35170 14602 35204 14636
rect 35260 14634 35294 14636
rect 35350 14634 35384 14636
rect 35440 14634 35474 14636
rect 35530 14634 35564 14636
rect 35620 14634 35654 14636
rect 35710 14634 35744 14636
rect 35800 14634 35834 14636
rect 35890 14634 35924 14636
rect 35980 14634 36014 14636
rect 35260 14602 35280 14634
rect 35280 14602 35294 14634
rect 35350 14602 35370 14634
rect 35370 14602 35384 14634
rect 35440 14602 35460 14634
rect 35460 14602 35474 14634
rect 35530 14602 35550 14634
rect 35550 14602 35564 14634
rect 35620 14602 35640 14634
rect 35640 14602 35654 14634
rect 35710 14602 35730 14634
rect 35730 14602 35744 14634
rect 35800 14602 35820 14634
rect 35820 14602 35834 14634
rect 35890 14602 35910 14634
rect 35910 14602 35924 14634
rect 35980 14602 36000 14634
rect 36000 14602 36014 14634
rect 36070 14602 36104 14636
rect 35356 14426 35378 14432
rect 35378 14426 35390 14432
rect 35456 14426 35468 14432
rect 35468 14426 35490 14432
rect 35556 14426 35558 14432
rect 35558 14426 35590 14432
rect 35356 14398 35390 14426
rect 35456 14398 35490 14426
rect 35556 14398 35590 14426
rect 35656 14398 35690 14432
rect 35756 14398 35790 14432
rect 35856 14426 35884 14432
rect 35884 14426 35890 14432
rect 35856 14398 35890 14426
rect 35356 14298 35390 14332
rect 35456 14298 35490 14332
rect 35556 14298 35590 14332
rect 35656 14298 35690 14332
rect 35756 14298 35790 14332
rect 35856 14298 35890 14332
rect 35356 14198 35390 14232
rect 35456 14198 35490 14232
rect 35556 14198 35590 14232
rect 35656 14198 35690 14232
rect 35756 14198 35790 14232
rect 35856 14198 35890 14232
rect 35356 14100 35390 14132
rect 35456 14100 35490 14132
rect 35556 14100 35590 14132
rect 35356 14098 35378 14100
rect 35378 14098 35390 14100
rect 35456 14098 35468 14100
rect 35468 14098 35490 14100
rect 35556 14098 35558 14100
rect 35558 14098 35590 14100
rect 35656 14098 35690 14132
rect 35756 14098 35790 14132
rect 35856 14100 35890 14132
rect 35856 14098 35884 14100
rect 35884 14098 35890 14100
rect 35356 14010 35390 14032
rect 35456 14010 35490 14032
rect 35556 14010 35590 14032
rect 35356 13998 35378 14010
rect 35378 13998 35390 14010
rect 35456 13998 35468 14010
rect 35468 13998 35490 14010
rect 35556 13998 35558 14010
rect 35558 13998 35590 14010
rect 35656 13998 35690 14032
rect 35756 13998 35790 14032
rect 35856 14010 35890 14032
rect 35856 13998 35884 14010
rect 35884 13998 35890 14010
rect 35356 13920 35390 13932
rect 35456 13920 35490 13932
rect 35556 13920 35590 13932
rect 35356 13898 35378 13920
rect 35378 13898 35390 13920
rect 35456 13898 35468 13920
rect 35468 13898 35490 13920
rect 35556 13898 35558 13920
rect 35558 13898 35590 13920
rect 35656 13898 35690 13932
rect 35756 13898 35790 13932
rect 35856 13920 35890 13932
rect 35856 13898 35884 13920
rect 35884 13898 35890 13920
rect 36510 14602 36544 14636
rect 36600 14634 36634 14636
rect 36690 14634 36724 14636
rect 36780 14634 36814 14636
rect 36870 14634 36904 14636
rect 36960 14634 36994 14636
rect 37050 14634 37084 14636
rect 37140 14634 37174 14636
rect 37230 14634 37264 14636
rect 37320 14634 37354 14636
rect 36600 14602 36620 14634
rect 36620 14602 36634 14634
rect 36690 14602 36710 14634
rect 36710 14602 36724 14634
rect 36780 14602 36800 14634
rect 36800 14602 36814 14634
rect 36870 14602 36890 14634
rect 36890 14602 36904 14634
rect 36960 14602 36980 14634
rect 36980 14602 36994 14634
rect 37050 14602 37070 14634
rect 37070 14602 37084 14634
rect 37140 14602 37160 14634
rect 37160 14602 37174 14634
rect 37230 14602 37250 14634
rect 37250 14602 37264 14634
rect 37320 14602 37340 14634
rect 37340 14602 37354 14634
rect 37410 14602 37444 14636
rect 36696 14426 36718 14432
rect 36718 14426 36730 14432
rect 36796 14426 36808 14432
rect 36808 14426 36830 14432
rect 36896 14426 36898 14432
rect 36898 14426 36930 14432
rect 36696 14398 36730 14426
rect 36796 14398 36830 14426
rect 36896 14398 36930 14426
rect 36996 14398 37030 14432
rect 37096 14398 37130 14432
rect 37196 14426 37224 14432
rect 37224 14426 37230 14432
rect 37196 14398 37230 14426
rect 36696 14298 36730 14332
rect 36796 14298 36830 14332
rect 36896 14298 36930 14332
rect 36996 14298 37030 14332
rect 37096 14298 37130 14332
rect 37196 14298 37230 14332
rect 36696 14198 36730 14232
rect 36796 14198 36830 14232
rect 36896 14198 36930 14232
rect 36996 14198 37030 14232
rect 37096 14198 37130 14232
rect 37196 14198 37230 14232
rect 36696 14100 36730 14132
rect 36796 14100 36830 14132
rect 36896 14100 36930 14132
rect 36696 14098 36718 14100
rect 36718 14098 36730 14100
rect 36796 14098 36808 14100
rect 36808 14098 36830 14100
rect 36896 14098 36898 14100
rect 36898 14098 36930 14100
rect 36996 14098 37030 14132
rect 37096 14098 37130 14132
rect 37196 14100 37230 14132
rect 37196 14098 37224 14100
rect 37224 14098 37230 14100
rect 36696 14010 36730 14032
rect 36796 14010 36830 14032
rect 36896 14010 36930 14032
rect 36696 13998 36718 14010
rect 36718 13998 36730 14010
rect 36796 13998 36808 14010
rect 36808 13998 36830 14010
rect 36896 13998 36898 14010
rect 36898 13998 36930 14010
rect 36996 13998 37030 14032
rect 37096 13998 37130 14032
rect 37196 14010 37230 14032
rect 37196 13998 37224 14010
rect 37224 13998 37230 14010
rect 36696 13920 36730 13932
rect 36796 13920 36830 13932
rect 36896 13920 36930 13932
rect 36696 13898 36718 13920
rect 36718 13898 36730 13920
rect 36796 13898 36808 13920
rect 36808 13898 36830 13920
rect 36896 13898 36898 13920
rect 36898 13898 36930 13920
rect 36996 13898 37030 13932
rect 37096 13898 37130 13932
rect 37196 13920 37230 13932
rect 37196 13898 37224 13920
rect 37224 13898 37230 13920
rect 37850 14602 37884 14636
rect 37940 14634 37974 14636
rect 38030 14634 38064 14636
rect 38120 14634 38154 14636
rect 38210 14634 38244 14636
rect 38300 14634 38334 14636
rect 38390 14634 38424 14636
rect 38480 14634 38514 14636
rect 38570 14634 38604 14636
rect 38660 14634 38694 14636
rect 37940 14602 37960 14634
rect 37960 14602 37974 14634
rect 38030 14602 38050 14634
rect 38050 14602 38064 14634
rect 38120 14602 38140 14634
rect 38140 14602 38154 14634
rect 38210 14602 38230 14634
rect 38230 14602 38244 14634
rect 38300 14602 38320 14634
rect 38320 14602 38334 14634
rect 38390 14602 38410 14634
rect 38410 14602 38424 14634
rect 38480 14602 38500 14634
rect 38500 14602 38514 14634
rect 38570 14602 38590 14634
rect 38590 14602 38604 14634
rect 38660 14602 38680 14634
rect 38680 14602 38694 14634
rect 38750 14602 38784 14636
rect 38036 14426 38058 14432
rect 38058 14426 38070 14432
rect 38136 14426 38148 14432
rect 38148 14426 38170 14432
rect 38236 14426 38238 14432
rect 38238 14426 38270 14432
rect 38036 14398 38070 14426
rect 38136 14398 38170 14426
rect 38236 14398 38270 14426
rect 38336 14398 38370 14432
rect 38436 14398 38470 14432
rect 38536 14426 38564 14432
rect 38564 14426 38570 14432
rect 38536 14398 38570 14426
rect 38036 14298 38070 14332
rect 38136 14298 38170 14332
rect 38236 14298 38270 14332
rect 38336 14298 38370 14332
rect 38436 14298 38470 14332
rect 38536 14298 38570 14332
rect 38036 14198 38070 14232
rect 38136 14198 38170 14232
rect 38236 14198 38270 14232
rect 38336 14198 38370 14232
rect 38436 14198 38470 14232
rect 38536 14198 38570 14232
rect 38036 14100 38070 14132
rect 38136 14100 38170 14132
rect 38236 14100 38270 14132
rect 38036 14098 38058 14100
rect 38058 14098 38070 14100
rect 38136 14098 38148 14100
rect 38148 14098 38170 14100
rect 38236 14098 38238 14100
rect 38238 14098 38270 14100
rect 38336 14098 38370 14132
rect 38436 14098 38470 14132
rect 38536 14100 38570 14132
rect 38536 14098 38564 14100
rect 38564 14098 38570 14100
rect 38036 14010 38070 14032
rect 38136 14010 38170 14032
rect 38236 14010 38270 14032
rect 38036 13998 38058 14010
rect 38058 13998 38070 14010
rect 38136 13998 38148 14010
rect 38148 13998 38170 14010
rect 38236 13998 38238 14010
rect 38238 13998 38270 14010
rect 38336 13998 38370 14032
rect 38436 13998 38470 14032
rect 38536 14010 38570 14032
rect 38536 13998 38564 14010
rect 38564 13998 38570 14010
rect 38036 13920 38070 13932
rect 38136 13920 38170 13932
rect 38236 13920 38270 13932
rect 38036 13898 38058 13920
rect 38058 13898 38070 13920
rect 38136 13898 38148 13920
rect 38148 13898 38170 13920
rect 38236 13898 38238 13920
rect 38238 13898 38270 13920
rect 38336 13898 38370 13932
rect 38436 13898 38470 13932
rect 38536 13920 38570 13932
rect 38536 13898 38564 13920
rect 38564 13898 38570 13920
rect 39275 14323 39669 14861
rect 41282 14323 41676 14861
rect 39275 13363 39669 13901
rect 41282 13363 41676 13901
rect 8079 13215 8113 13249
rect 8279 13215 8313 13249
rect 8479 13215 8513 13249
rect 8679 13215 8713 13249
rect 8879 13215 8913 13249
rect 9079 13215 9113 13249
rect 9279 13215 9313 13249
rect 9479 13215 9513 13249
rect 9679 13215 9713 13249
rect 9879 13215 9913 13249
rect 10079 13215 10113 13249
rect 10823 13215 10857 13249
rect 11023 13215 11057 13249
rect 11223 13215 11257 13249
rect 11423 13215 11457 13249
rect 11623 13215 11657 13249
rect 11823 13215 11857 13249
rect 12023 13215 12057 13249
rect 12223 13215 12257 13249
rect 12423 13215 12457 13249
rect 12623 13215 12657 13249
rect 12823 13215 12857 13249
rect 13567 13215 13601 13249
rect 13767 13215 13801 13249
rect 13967 13215 14001 13249
rect 14167 13215 14201 13249
rect 14367 13215 14401 13249
rect 14567 13215 14601 13249
rect 14767 13215 14801 13249
rect 14967 13215 15001 13249
rect 15167 13215 15201 13249
rect 15367 13215 15401 13249
rect 15567 13215 15601 13249
rect 16293 13215 16327 13249
rect 16693 13215 16727 13249
rect 17093 13215 17127 13249
rect 17493 13215 17527 13249
rect 17893 13215 17927 13249
rect 18293 13215 18327 13249
rect 18693 13215 18727 13249
rect 19093 13215 19127 13249
rect 19493 13215 19527 13249
rect 19893 13215 19927 13249
rect 20293 13215 20327 13249
rect 20693 13215 20727 13249
rect 21093 13215 21127 13249
rect 21493 13215 21527 13249
rect 21893 13215 21927 13249
rect 22293 13215 22327 13249
rect 22693 13215 22727 13249
rect 23093 13215 23127 13249
rect 23759 13215 23793 13249
rect 23959 13215 23993 13249
rect 24159 13215 24193 13249
rect 24359 13215 24393 13249
rect 24559 13215 24593 13249
rect 24759 13215 24793 13249
rect 24959 13215 24993 13249
rect 25159 13215 25193 13249
rect 25359 13215 25393 13249
rect 25559 13215 25593 13249
rect 25759 13215 25793 13249
rect 28443 13215 28477 13249
rect 28643 13215 28677 13249
rect 28843 13215 28877 13249
rect 29043 13215 29077 13249
rect 29243 13215 29277 13249
rect 29443 13215 29477 13249
rect 29643 13215 29677 13249
rect 29843 13215 29877 13249
rect 30043 13215 30077 13249
rect 30243 13215 30277 13249
rect 30443 13215 30477 13249
rect 30643 13215 30677 13249
rect 30843 13215 30877 13249
rect 31043 13215 31077 13249
rect 31243 13215 31277 13249
rect 31443 13215 31477 13249
rect 31643 13215 31677 13249
rect 31843 13215 31877 13249
rect 32043 13215 32077 13249
rect 32243 13215 32277 13249
rect 32443 13215 32477 13249
rect 32643 13215 32677 13249
rect 32843 13215 32877 13249
rect 33043 13215 33077 13249
rect 33243 13215 33277 13249
rect 33443 13215 33477 13249
rect 33643 13215 33677 13249
rect 33843 13215 33877 13249
rect 34043 13215 34077 13249
rect 34243 13215 34277 13249
rect 34443 13215 34477 13249
rect 34643 13215 34677 13249
rect 34843 13215 34877 13249
rect 35043 13215 35077 13249
rect 35243 13215 35277 13249
rect 35443 13215 35477 13249
rect 35643 13215 35677 13249
rect 35843 13215 35877 13249
rect 36043 13215 36077 13249
rect 36243 13215 36277 13249
rect 36443 13215 36477 13249
rect 36643 13215 36677 13249
rect 36843 13215 36877 13249
rect 37043 13215 37077 13249
rect 37243 13215 37277 13249
rect 37443 13215 37477 13249
rect 37643 13215 37677 13249
rect 37843 13215 37877 13249
rect 38043 13215 38077 13249
rect 38243 13215 38277 13249
rect 38443 13215 38477 13249
rect 38643 13215 38677 13249
rect 38843 13215 38877 13249
rect 39439 13215 39473 13249
rect 39639 13215 39673 13249
rect 39839 13215 39873 13249
rect 40039 13215 40073 13249
rect 40239 13215 40273 13249
rect 40439 13215 40473 13249
rect 40639 13215 40673 13249
rect 40839 13215 40873 13249
rect 41039 13215 41073 13249
rect 41239 13215 41273 13249
rect 41439 13215 41473 13249
rect 8079 11335 8113 11369
rect 8279 11335 8313 11369
rect 8479 11335 8513 11369
rect 8679 11335 8713 11369
rect 8879 11335 8913 11369
rect 9079 11335 9113 11369
rect 9279 11335 9313 11369
rect 9479 11335 9513 11369
rect 9679 11335 9713 11369
rect 9879 11335 9913 11369
rect 10079 11335 10113 11369
rect 10823 11335 10857 11369
rect 11023 11335 11057 11369
rect 11223 11335 11257 11369
rect 11423 11335 11457 11369
rect 11623 11335 11657 11369
rect 11823 11335 11857 11369
rect 12023 11335 12057 11369
rect 12223 11335 12257 11369
rect 12423 11335 12457 11369
rect 12623 11335 12657 11369
rect 12823 11335 12857 11369
rect 13567 11335 13601 11369
rect 13767 11335 13801 11369
rect 13967 11335 14001 11369
rect 14167 11335 14201 11369
rect 14367 11335 14401 11369
rect 14567 11335 14601 11369
rect 14767 11335 14801 11369
rect 14967 11335 15001 11369
rect 15167 11335 15201 11369
rect 15367 11335 15401 11369
rect 15567 11335 15601 11369
rect 16293 11335 16327 11369
rect 16693 11335 16727 11369
rect 17093 11335 17127 11369
rect 17493 11335 17527 11369
rect 17893 11335 17927 11369
rect 18293 11335 18327 11369
rect 18693 11335 18727 11369
rect 19093 11335 19127 11369
rect 19493 11335 19527 11369
rect 19893 11335 19927 11369
rect 20293 11335 20327 11369
rect 20693 11335 20727 11369
rect 21093 11335 21127 11369
rect 21493 11335 21527 11369
rect 21893 11335 21927 11369
rect 22293 11335 22327 11369
rect 22693 11335 22727 11369
rect 23093 11335 23127 11369
rect 23761 11335 23795 11369
rect 23961 11335 23995 11369
rect 24161 11335 24195 11369
rect 24361 11335 24395 11369
rect 24561 11335 24595 11369
rect 24761 11335 24795 11369
rect 24961 11335 24995 11369
rect 25161 11335 25195 11369
rect 25361 11335 25395 11369
rect 25561 11335 25595 11369
rect 25761 11335 25795 11369
rect 25961 11335 25995 11369
rect 26161 11335 26195 11369
rect 26361 11335 26395 11369
rect 27091 11335 27125 11369
rect 27291 11335 27325 11369
rect 27491 11335 27525 11369
rect 27691 11335 27725 11369
rect 27891 11335 27925 11369
rect 28091 11335 28125 11369
rect 28291 11335 28325 11369
rect 28491 11335 28525 11369
rect 28691 11335 28725 11369
rect 28891 11335 28925 11369
rect 29091 11335 29125 11369
rect 29835 11335 29869 11369
rect 30035 11335 30069 11369
rect 30235 11335 30269 11369
rect 30435 11335 30469 11369
rect 30635 11335 30669 11369
rect 30835 11335 30869 11369
rect 31035 11335 31069 11369
rect 31235 11335 31269 11369
rect 31435 11335 31469 11369
rect 31635 11335 31669 11369
rect 31835 11335 31869 11369
rect 32579 11335 32613 11369
rect 32779 11335 32813 11369
rect 32979 11335 33013 11369
rect 33179 11335 33213 11369
rect 33379 11335 33413 11369
rect 33579 11335 33613 11369
rect 33779 11335 33813 11369
rect 33979 11335 34013 11369
rect 34179 11335 34213 11369
rect 34379 11335 34413 11369
rect 34579 11335 34613 11369
rect 35323 11335 35357 11369
rect 35523 11335 35557 11369
rect 35723 11335 35757 11369
rect 35923 11335 35957 11369
rect 36123 11335 36157 11369
rect 36323 11335 36357 11369
rect 36523 11335 36557 11369
rect 36723 11335 36757 11369
rect 36923 11335 36957 11369
rect 37123 11335 37157 11369
rect 37323 11335 37357 11369
rect 38067 11335 38101 11369
rect 38267 11335 38301 11369
rect 38467 11335 38501 11369
rect 38667 11335 38701 11369
rect 38867 11335 38901 11369
rect 39067 11335 39101 11369
rect 39267 11335 39301 11369
rect 39467 11335 39501 11369
rect 39667 11335 39701 11369
rect 39867 11335 39901 11369
rect 40067 11335 40101 11369
rect 7915 10563 8309 11101
rect 9922 10563 10316 11101
rect 10659 10563 11053 11101
rect 12666 10563 13060 11101
rect 13403 10563 13797 11101
rect 15410 10563 15804 11101
rect 23596 10563 23990 11101
rect 26177 10563 26571 11101
rect 26927 10563 27321 11101
rect 28934 10563 29328 11101
rect 29671 10563 30065 11101
rect 31678 10563 32072 11101
rect 32415 10563 32809 11101
rect 34422 10563 34816 11101
rect 35159 10563 35553 11101
rect 37166 10563 37560 11101
rect 37903 10563 38297 11101
rect 39910 10563 40304 11101
rect 7915 9603 8309 10141
rect 9922 9603 10316 10141
rect 10659 9603 11053 10141
rect 12666 9603 13060 10141
rect 13403 9603 13797 10141
rect 15410 9603 15804 10141
rect 23596 9603 23990 10141
rect 26177 9603 26571 10141
rect 26927 9603 27321 10141
rect 28934 9603 29328 10141
rect 29671 9603 30065 10141
rect 31678 9603 32072 10141
rect 32415 9603 32809 10141
rect 34422 9603 34816 10141
rect 35159 9603 35553 10141
rect 37166 9603 37560 10141
rect 37903 9603 38297 10141
rect 39910 9603 40304 10141
rect 8079 9455 8113 9489
rect 8279 9455 8313 9489
rect 8479 9455 8513 9489
rect 8679 9455 8713 9489
rect 8879 9455 8913 9489
rect 9079 9455 9113 9489
rect 9279 9455 9313 9489
rect 9479 9455 9513 9489
rect 9679 9455 9713 9489
rect 9879 9455 9913 9489
rect 10079 9455 10113 9489
rect 10823 9455 10857 9489
rect 11023 9455 11057 9489
rect 11223 9455 11257 9489
rect 11423 9455 11457 9489
rect 11623 9455 11657 9489
rect 11823 9455 11857 9489
rect 12023 9455 12057 9489
rect 12223 9455 12257 9489
rect 12423 9455 12457 9489
rect 12623 9455 12657 9489
rect 12823 9455 12857 9489
rect 13567 9455 13601 9489
rect 13767 9455 13801 9489
rect 13967 9455 14001 9489
rect 14167 9455 14201 9489
rect 14367 9455 14401 9489
rect 14567 9455 14601 9489
rect 14767 9455 14801 9489
rect 14967 9455 15001 9489
rect 15167 9455 15201 9489
rect 15367 9455 15401 9489
rect 15567 9455 15601 9489
rect 16293 9455 16327 9489
rect 16693 9455 16727 9489
rect 17093 9455 17127 9489
rect 17493 9455 17527 9489
rect 17893 9455 17927 9489
rect 18293 9455 18327 9489
rect 18693 9455 18727 9489
rect 19093 9455 19127 9489
rect 19493 9455 19527 9489
rect 19893 9455 19927 9489
rect 20293 9455 20327 9489
rect 20693 9455 20727 9489
rect 21093 9455 21127 9489
rect 21493 9455 21527 9489
rect 21893 9455 21927 9489
rect 22293 9455 22327 9489
rect 22693 9455 22727 9489
rect 23093 9455 23127 9489
rect 23761 9455 23795 9489
rect 23961 9455 23995 9489
rect 24161 9455 24195 9489
rect 24361 9455 24395 9489
rect 24561 9455 24595 9489
rect 24761 9455 24795 9489
rect 24961 9455 24995 9489
rect 25161 9455 25195 9489
rect 25361 9455 25395 9489
rect 25561 9455 25595 9489
rect 25761 9455 25795 9489
rect 25961 9455 25995 9489
rect 26161 9455 26195 9489
rect 26361 9455 26395 9489
rect 27091 9455 27125 9489
rect 27291 9455 27325 9489
rect 27491 9455 27525 9489
rect 27691 9455 27725 9489
rect 27891 9455 27925 9489
rect 28091 9455 28125 9489
rect 28291 9455 28325 9489
rect 28491 9455 28525 9489
rect 28691 9455 28725 9489
rect 28891 9455 28925 9489
rect 29091 9455 29125 9489
rect 29835 9455 29869 9489
rect 30035 9455 30069 9489
rect 30235 9455 30269 9489
rect 30435 9455 30469 9489
rect 30635 9455 30669 9489
rect 30835 9455 30869 9489
rect 31035 9455 31069 9489
rect 31235 9455 31269 9489
rect 31435 9455 31469 9489
rect 31635 9455 31669 9489
rect 31835 9455 31869 9489
rect 32579 9455 32613 9489
rect 32779 9455 32813 9489
rect 32979 9455 33013 9489
rect 33179 9455 33213 9489
rect 33379 9455 33413 9489
rect 33579 9455 33613 9489
rect 33779 9455 33813 9489
rect 33979 9455 34013 9489
rect 34179 9455 34213 9489
rect 34379 9455 34413 9489
rect 34579 9455 34613 9489
rect 35323 9455 35357 9489
rect 35523 9455 35557 9489
rect 35723 9455 35757 9489
rect 35923 9455 35957 9489
rect 36123 9455 36157 9489
rect 36323 9455 36357 9489
rect 36523 9455 36557 9489
rect 36723 9455 36757 9489
rect 36923 9455 36957 9489
rect 37123 9455 37157 9489
rect 37323 9455 37357 9489
rect 38067 9455 38101 9489
rect 38267 9455 38301 9489
rect 38467 9455 38501 9489
rect 38667 9455 38701 9489
rect 38867 9455 38901 9489
rect 39067 9455 39101 9489
rect 39267 9455 39301 9489
rect 39467 9455 39501 9489
rect 39667 9455 39701 9489
rect 39867 9455 39901 9489
rect 40067 9455 40101 9489
rect 8079 7575 8113 7609
rect 8279 7575 8313 7609
rect 8479 7575 8513 7609
rect 8679 7575 8713 7609
rect 8879 7575 8913 7609
rect 9079 7575 9113 7609
rect 9279 7575 9313 7609
rect 9479 7575 9513 7609
rect 9679 7575 9713 7609
rect 9879 7575 9913 7609
rect 10079 7575 10113 7609
rect 14451 7575 14485 7609
rect 14651 7575 14685 7609
rect 14851 7575 14885 7609
rect 15051 7575 15085 7609
rect 15251 7575 15285 7609
rect 15451 7575 15485 7609
rect 15651 7575 15685 7609
rect 15851 7575 15885 7609
rect 16051 7575 16085 7609
rect 16251 7575 16285 7609
rect 16451 7575 16485 7609
rect 16651 7575 16685 7609
rect 16851 7575 16885 7609
rect 17051 7575 17085 7609
rect 17781 7575 17815 7609
rect 17981 7575 18015 7609
rect 18181 7575 18215 7609
rect 18381 7575 18415 7609
rect 18581 7575 18615 7609
rect 18781 7575 18815 7609
rect 18981 7575 19015 7609
rect 19181 7575 19215 7609
rect 19381 7575 19415 7609
rect 19581 7575 19615 7609
rect 19781 7575 19815 7609
rect 20525 7575 20559 7609
rect 20725 7575 20759 7609
rect 20925 7575 20959 7609
rect 21125 7575 21159 7609
rect 21325 7575 21359 7609
rect 21525 7575 21559 7609
rect 21725 7575 21759 7609
rect 21925 7575 21959 7609
rect 22125 7575 22159 7609
rect 22325 7575 22359 7609
rect 22525 7575 22559 7609
rect 23269 7575 23303 7609
rect 23469 7575 23503 7609
rect 23669 7575 23703 7609
rect 23869 7575 23903 7609
rect 24069 7575 24103 7609
rect 24269 7575 24303 7609
rect 24469 7575 24503 7609
rect 24669 7575 24703 7609
rect 24869 7575 24903 7609
rect 25069 7575 25103 7609
rect 25269 7575 25303 7609
rect 26013 7575 26047 7609
rect 26213 7575 26247 7609
rect 26413 7575 26447 7609
rect 26613 7575 26647 7609
rect 26813 7575 26847 7609
rect 27013 7575 27047 7609
rect 27213 7575 27247 7609
rect 27413 7575 27447 7609
rect 27613 7575 27647 7609
rect 27813 7575 27847 7609
rect 28013 7575 28047 7609
rect 28757 7575 28791 7609
rect 28957 7575 28991 7609
rect 29157 7575 29191 7609
rect 29357 7575 29391 7609
rect 29557 7575 29591 7609
rect 29757 7575 29791 7609
rect 29957 7575 29991 7609
rect 30157 7575 30191 7609
rect 30357 7575 30391 7609
rect 30557 7575 30591 7609
rect 30757 7575 30791 7609
rect 31501 7575 31535 7609
rect 31701 7575 31735 7609
rect 31901 7575 31935 7609
rect 32101 7575 32135 7609
rect 32301 7575 32335 7609
rect 32501 7575 32535 7609
rect 32701 7575 32735 7609
rect 32901 7575 32935 7609
rect 33101 7575 33135 7609
rect 33301 7575 33335 7609
rect 33501 7575 33535 7609
rect 35323 7575 35357 7609
rect 35523 7575 35557 7609
rect 35723 7575 35757 7609
rect 35923 7575 35957 7609
rect 36123 7575 36157 7609
rect 36323 7575 36357 7609
rect 36523 7575 36557 7609
rect 36723 7575 36757 7609
rect 36923 7575 36957 7609
rect 37123 7575 37157 7609
rect 37323 7575 37357 7609
rect 38067 7575 38101 7609
rect 38267 7575 38301 7609
rect 38467 7575 38501 7609
rect 38667 7575 38701 7609
rect 38867 7575 38901 7609
rect 39067 7575 39101 7609
rect 39267 7575 39301 7609
rect 39467 7575 39501 7609
rect 39667 7575 39701 7609
rect 39867 7575 39901 7609
rect 40067 7575 40101 7609
rect 7915 6803 8309 7341
rect 9922 6803 10316 7341
rect 14286 6803 14680 7341
rect 16867 6803 17261 7341
rect 17617 6803 18011 7341
rect 19624 6803 20018 7341
rect 20361 6803 20755 7341
rect 22368 6803 22762 7341
rect 23105 6803 23499 7341
rect 25112 6803 25506 7341
rect 25849 6803 26243 7341
rect 27856 6803 28250 7341
rect 28593 6803 28987 7341
rect 30600 6803 30994 7341
rect 31337 6803 31731 7341
rect 33344 6803 33738 7341
rect 35159 6803 35553 7341
rect 37166 6803 37560 7341
rect 37903 6803 38297 7341
rect 39910 6803 40304 7341
rect 7915 5843 8309 6381
rect 9922 5843 10316 6381
rect 14286 5843 14680 6381
rect 16867 5843 17261 6381
rect 17617 5843 18011 6381
rect 19624 5843 20018 6381
rect 20361 5843 20755 6381
rect 22368 5843 22762 6381
rect 23105 5843 23499 6381
rect 25112 5843 25506 6381
rect 25849 5843 26243 6381
rect 27856 5843 28250 6381
rect 28593 5843 28987 6381
rect 30600 5843 30994 6381
rect 31337 5843 31731 6381
rect 33344 5843 33738 6381
rect 35159 5843 35553 6381
rect 37166 5843 37560 6381
rect 37903 5843 38297 6381
rect 39910 5843 40304 6381
rect 8079 5695 8113 5729
rect 8279 5695 8313 5729
rect 8479 5695 8513 5729
rect 8679 5695 8713 5729
rect 8879 5695 8913 5729
rect 9079 5695 9113 5729
rect 9279 5695 9313 5729
rect 9479 5695 9513 5729
rect 9679 5695 9713 5729
rect 9879 5695 9913 5729
rect 10079 5695 10113 5729
rect 14451 5695 14485 5729
rect 14651 5695 14685 5729
rect 14851 5695 14885 5729
rect 15051 5695 15085 5729
rect 15251 5695 15285 5729
rect 15451 5695 15485 5729
rect 15651 5695 15685 5729
rect 15851 5695 15885 5729
rect 16051 5695 16085 5729
rect 16251 5695 16285 5729
rect 16451 5695 16485 5729
rect 16651 5695 16685 5729
rect 16851 5695 16885 5729
rect 17051 5695 17085 5729
rect 17781 5695 17815 5729
rect 17981 5695 18015 5729
rect 18181 5695 18215 5729
rect 18381 5695 18415 5729
rect 18581 5695 18615 5729
rect 18781 5695 18815 5729
rect 18981 5695 19015 5729
rect 19181 5695 19215 5729
rect 19381 5695 19415 5729
rect 19581 5695 19615 5729
rect 19781 5695 19815 5729
rect 20525 5695 20559 5729
rect 20725 5695 20759 5729
rect 20925 5695 20959 5729
rect 21125 5695 21159 5729
rect 21325 5695 21359 5729
rect 21525 5695 21559 5729
rect 21725 5695 21759 5729
rect 21925 5695 21959 5729
rect 22125 5695 22159 5729
rect 22325 5695 22359 5729
rect 22525 5695 22559 5729
rect 23269 5695 23303 5729
rect 23469 5695 23503 5729
rect 23669 5695 23703 5729
rect 23869 5695 23903 5729
rect 24069 5695 24103 5729
rect 24269 5695 24303 5729
rect 24469 5695 24503 5729
rect 24669 5695 24703 5729
rect 24869 5695 24903 5729
rect 25069 5695 25103 5729
rect 25269 5695 25303 5729
rect 26013 5695 26047 5729
rect 26213 5695 26247 5729
rect 26413 5695 26447 5729
rect 26613 5695 26647 5729
rect 26813 5695 26847 5729
rect 27013 5695 27047 5729
rect 27213 5695 27247 5729
rect 27413 5695 27447 5729
rect 27613 5695 27647 5729
rect 27813 5695 27847 5729
rect 28013 5695 28047 5729
rect 28757 5695 28791 5729
rect 28957 5695 28991 5729
rect 29157 5695 29191 5729
rect 29357 5695 29391 5729
rect 29557 5695 29591 5729
rect 29757 5695 29791 5729
rect 29957 5695 29991 5729
rect 30157 5695 30191 5729
rect 30357 5695 30391 5729
rect 30557 5695 30591 5729
rect 30757 5695 30791 5729
rect 31501 5695 31535 5729
rect 31701 5695 31735 5729
rect 31901 5695 31935 5729
rect 32101 5695 32135 5729
rect 32301 5695 32335 5729
rect 32501 5695 32535 5729
rect 32701 5695 32735 5729
rect 32901 5695 32935 5729
rect 33101 5695 33135 5729
rect 33301 5695 33335 5729
rect 33501 5695 33535 5729
rect 35323 5695 35357 5729
rect 35523 5695 35557 5729
rect 35723 5695 35757 5729
rect 35923 5695 35957 5729
rect 36123 5695 36157 5729
rect 36323 5695 36357 5729
rect 36523 5695 36557 5729
rect 36723 5695 36757 5729
rect 36923 5695 36957 5729
rect 37123 5695 37157 5729
rect 37323 5695 37357 5729
rect 38067 5695 38101 5729
rect 38267 5695 38301 5729
rect 38467 5695 38501 5729
rect 38667 5695 38701 5729
rect 38867 5695 38901 5729
rect 39067 5695 39101 5729
rect 39267 5695 39301 5729
rect 39467 5695 39501 5729
rect 39667 5695 39701 5729
rect 39867 5695 39901 5729
rect 40067 5695 40101 5729
<< metal1 >>
rect 3348 41490 45288 41492
rect 3348 41374 3370 41490
rect 4958 41472 43678 41490
rect 4958 41449 12440 41472
rect 4958 41415 6167 41449
rect 6201 41415 6983 41449
rect 7017 41415 7383 41449
rect 7417 41415 7783 41449
rect 7817 41415 8183 41449
rect 8217 41415 8583 41449
rect 8617 41415 8983 41449
rect 9017 41415 9383 41449
rect 9417 41415 9783 41449
rect 9817 41415 10183 41449
rect 10217 41415 10583 41449
rect 10617 41415 10983 41449
rect 11017 41415 11383 41449
rect 11417 41415 11783 41449
rect 11817 41415 12183 41449
rect 12217 41420 12440 41449
rect 12492 41449 43678 41472
rect 12492 41420 12583 41449
rect 12217 41415 12583 41420
rect 12617 41415 12983 41449
rect 13017 41415 13383 41449
rect 13417 41415 13783 41449
rect 13817 41415 15213 41449
rect 15247 41415 15613 41449
rect 15647 41415 16013 41449
rect 16047 41415 16413 41449
rect 16447 41415 16813 41449
rect 16847 41415 17213 41449
rect 17247 41415 17613 41449
rect 17647 41415 18013 41449
rect 18047 41415 18413 41449
rect 18447 41415 18813 41449
rect 18847 41415 19213 41449
rect 19247 41415 19613 41449
rect 19647 41415 20013 41449
rect 20047 41415 20413 41449
rect 20447 41415 20813 41449
rect 20847 41415 21213 41449
rect 21247 41415 21613 41449
rect 21647 41415 22013 41449
rect 22047 41415 22413 41449
rect 22447 41415 22813 41449
rect 22847 41415 23213 41449
rect 23247 41415 23613 41449
rect 23647 41415 24013 41449
rect 24047 41415 24413 41449
rect 24447 41415 24813 41449
rect 24847 41415 25213 41449
rect 25247 41415 25613 41449
rect 25647 41415 26013 41449
rect 26047 41415 26413 41449
rect 26447 41415 26813 41449
rect 26847 41415 27213 41449
rect 27247 41415 27613 41449
rect 27647 41415 28013 41449
rect 28047 41415 28413 41449
rect 28447 41415 28813 41449
rect 28847 41415 29213 41449
rect 29247 41415 29613 41449
rect 29647 41415 30013 41449
rect 30047 41415 30413 41449
rect 30447 41415 30813 41449
rect 30847 41415 31213 41449
rect 31247 41415 31613 41449
rect 31647 41415 32013 41449
rect 32047 41415 32413 41449
rect 32447 41415 32813 41449
rect 32847 41415 33213 41449
rect 33247 41415 33613 41449
rect 33647 41415 34013 41449
rect 34047 41415 34413 41449
rect 34447 41415 34813 41449
rect 34847 41415 35213 41449
rect 35247 41415 35613 41449
rect 35647 41415 36013 41449
rect 36047 41415 36413 41449
rect 36447 41415 36813 41449
rect 36847 41415 37213 41449
rect 37247 41415 37613 41449
rect 37647 41415 38013 41449
rect 38047 41415 38413 41449
rect 38447 41415 38813 41449
rect 38847 41415 39213 41449
rect 39247 41415 39613 41449
rect 39647 41415 40013 41449
rect 40047 41415 40413 41449
rect 40447 41415 40813 41449
rect 40847 41415 41213 41449
rect 41247 41415 41613 41449
rect 41647 41415 42013 41449
rect 42047 41415 42413 41449
rect 42447 41415 43678 41449
rect 4958 41374 43678 41415
rect 45266 41374 45288 41490
rect 3348 41372 45288 41374
rect 25608 41197 25636 41372
rect 15071 41181 15117 41197
rect 15071 41147 15077 41181
rect 15111 41147 15117 41181
rect 15071 41109 15117 41147
rect 15071 41075 15077 41109
rect 15111 41075 15117 41109
rect 15071 41037 15117 41075
rect 15071 41003 15077 41037
rect 15111 41003 15117 41037
rect 15071 40965 15117 41003
rect 5990 40929 6036 40952
rect 5990 40895 5996 40929
rect 6030 40895 6036 40929
rect 5990 40857 6036 40895
rect 5990 40823 5996 40857
rect 6030 40823 6036 40857
rect 5990 40785 6036 40823
rect 5990 40751 5996 40785
rect 6030 40751 6036 40785
rect 5990 40713 6036 40751
rect 5990 40679 5996 40713
rect 6030 40679 6036 40713
rect 5990 40641 6036 40679
rect 5990 40607 5996 40641
rect 6030 40607 6036 40641
rect 5990 40569 6036 40607
rect 5990 40535 5996 40569
rect 6030 40535 6036 40569
rect 5990 40497 6036 40535
rect 5990 40463 5996 40497
rect 6030 40463 6036 40497
rect 5990 40425 6036 40463
rect 5990 40391 5996 40425
rect 6030 40391 6036 40425
rect 5990 40353 6036 40391
rect 5990 40319 5996 40353
rect 6030 40319 6036 40353
rect 5990 40281 6036 40319
rect 5990 40247 5996 40281
rect 6030 40247 6036 40281
rect 5990 40209 6036 40247
rect 6448 40929 6494 40952
rect 6448 40895 6454 40929
rect 6488 40895 6494 40929
rect 6448 40857 6494 40895
rect 6448 40823 6454 40857
rect 6488 40823 6494 40857
rect 6448 40785 6494 40823
rect 6448 40751 6454 40785
rect 6488 40751 6494 40785
rect 6448 40713 6494 40751
rect 6448 40679 6454 40713
rect 6488 40679 6494 40713
rect 6448 40641 6494 40679
rect 6448 40607 6454 40641
rect 6488 40607 6494 40641
rect 6448 40569 6494 40607
rect 6448 40535 6454 40569
rect 6488 40535 6494 40569
rect 6448 40497 6494 40535
rect 6448 40463 6454 40497
rect 6488 40463 6494 40497
rect 6448 40425 6494 40463
rect 6448 40391 6454 40425
rect 6488 40391 6494 40425
rect 6448 40353 6494 40391
rect 6448 40319 6454 40353
rect 6488 40319 6494 40353
rect 6448 40281 6494 40319
rect 6448 40247 6454 40281
rect 6488 40247 6494 40281
rect 6448 40236 6494 40247
rect 5990 40175 5996 40209
rect 6030 40175 6036 40209
rect 5990 40152 6036 40175
rect 6380 40209 6494 40236
rect 6380 40208 6454 40209
rect 6380 39612 6408 40208
rect 6448 40175 6454 40208
rect 6488 40175 6494 40209
rect 6448 40152 6494 40175
rect 15071 40931 15077 40965
rect 15111 40931 15117 40965
rect 15071 40893 15117 40931
rect 15071 40859 15077 40893
rect 15111 40859 15117 40893
rect 15071 40821 15117 40859
rect 15071 40787 15077 40821
rect 15111 40787 15117 40821
rect 15071 40749 15117 40787
rect 15071 40715 15077 40749
rect 15111 40715 15117 40749
rect 15071 40677 15117 40715
rect 15071 40643 15077 40677
rect 15111 40643 15117 40677
rect 15071 40605 15117 40643
rect 15071 40571 15077 40605
rect 15111 40571 15117 40605
rect 15071 40533 15117 40571
rect 15071 40499 15077 40533
rect 15111 40499 15117 40533
rect 15071 40461 15117 40499
rect 15071 40427 15077 40461
rect 15111 40427 15117 40461
rect 15071 40389 15117 40427
rect 15071 40355 15077 40389
rect 15111 40355 15117 40389
rect 15071 40317 15117 40355
rect 15071 40283 15077 40317
rect 15111 40283 15117 40317
rect 15071 40245 15117 40283
rect 15071 40211 15077 40245
rect 15111 40211 15117 40245
rect 15071 40173 15117 40211
rect 15071 40139 15077 40173
rect 15111 40139 15117 40173
rect 15071 40101 15117 40139
rect 15071 40067 15077 40101
rect 15111 40067 15117 40101
rect 15071 40029 15117 40067
rect 15071 39995 15077 40029
rect 15111 39995 15117 40029
rect 6457 39967 6515 39973
rect 6457 39933 6469 39967
rect 6503 39933 6515 39967
rect 6457 39927 6515 39933
rect 15071 39957 15117 39995
rect 6472 39769 6500 39927
rect 15071 39923 15077 39957
rect 15111 39923 15117 39957
rect 15071 39907 15117 39923
rect 15529 41181 15575 41197
rect 15529 41147 15535 41181
rect 15569 41147 15575 41181
rect 15529 41109 15575 41147
rect 15529 41075 15535 41109
rect 15569 41075 15575 41109
rect 15529 41037 15575 41075
rect 15529 41003 15535 41037
rect 15569 41003 15575 41037
rect 15529 40965 15575 41003
rect 15529 40931 15535 40965
rect 15569 40931 15575 40965
rect 15529 40893 15575 40931
rect 15529 40859 15535 40893
rect 15569 40859 15575 40893
rect 15529 40821 15575 40859
rect 15529 40787 15535 40821
rect 15569 40787 15575 40821
rect 15529 40749 15575 40787
rect 15529 40715 15535 40749
rect 15569 40715 15575 40749
rect 15529 40677 15575 40715
rect 15529 40643 15535 40677
rect 15569 40643 15575 40677
rect 15529 40605 15575 40643
rect 15529 40571 15535 40605
rect 15569 40571 15575 40605
rect 15529 40533 15575 40571
rect 15529 40499 15535 40533
rect 15569 40499 15575 40533
rect 15529 40461 15575 40499
rect 15529 40427 15535 40461
rect 15569 40427 15575 40461
rect 15529 40389 15575 40427
rect 15529 40355 15535 40389
rect 15569 40355 15575 40389
rect 15529 40317 15575 40355
rect 15529 40283 15535 40317
rect 15569 40283 15575 40317
rect 15529 40245 15575 40283
rect 15529 40211 15535 40245
rect 15569 40211 15575 40245
rect 15529 40173 15575 40211
rect 15529 40139 15535 40173
rect 15569 40139 15575 40173
rect 15529 40101 15575 40139
rect 15529 40067 15535 40101
rect 15569 40067 15575 40101
rect 15529 40029 15575 40067
rect 15529 39995 15535 40029
rect 15569 39995 15575 40029
rect 15529 39957 15575 39995
rect 15529 39923 15535 39957
rect 15569 39923 15575 39957
rect 15529 39907 15575 39923
rect 15987 41181 16033 41197
rect 15987 41147 15993 41181
rect 16027 41147 16033 41181
rect 15987 41109 16033 41147
rect 15987 41075 15993 41109
rect 16027 41075 16033 41109
rect 15987 41037 16033 41075
rect 15987 41003 15993 41037
rect 16027 41003 16033 41037
rect 15987 40965 16033 41003
rect 15987 40931 15993 40965
rect 16027 40931 16033 40965
rect 15987 40893 16033 40931
rect 15987 40859 15993 40893
rect 16027 40859 16033 40893
rect 15987 40821 16033 40859
rect 15987 40787 15993 40821
rect 16027 40787 16033 40821
rect 15987 40749 16033 40787
rect 15987 40715 15993 40749
rect 16027 40715 16033 40749
rect 15987 40677 16033 40715
rect 15987 40643 15993 40677
rect 16027 40643 16033 40677
rect 15987 40605 16033 40643
rect 15987 40571 15993 40605
rect 16027 40571 16033 40605
rect 15987 40533 16033 40571
rect 15987 40499 15993 40533
rect 16027 40499 16033 40533
rect 15987 40461 16033 40499
rect 15987 40427 15993 40461
rect 16027 40427 16033 40461
rect 15987 40389 16033 40427
rect 15987 40355 15993 40389
rect 16027 40355 16033 40389
rect 15987 40317 16033 40355
rect 15987 40283 15993 40317
rect 16027 40283 16033 40317
rect 15987 40245 16033 40283
rect 15987 40211 15993 40245
rect 16027 40211 16033 40245
rect 15987 40173 16033 40211
rect 15987 40139 15993 40173
rect 16027 40139 16033 40173
rect 15987 40101 16033 40139
rect 15987 40067 15993 40101
rect 16027 40067 16033 40101
rect 15987 40029 16033 40067
rect 15987 39995 15993 40029
rect 16027 39995 16033 40029
rect 15987 39957 16033 39995
rect 15987 39923 15993 39957
rect 16027 39923 16033 39957
rect 15987 39907 16033 39923
rect 16445 41181 16491 41197
rect 16445 41147 16451 41181
rect 16485 41147 16491 41181
rect 16445 41109 16491 41147
rect 16445 41075 16451 41109
rect 16485 41075 16491 41109
rect 16445 41037 16491 41075
rect 16445 41003 16451 41037
rect 16485 41003 16491 41037
rect 16445 40965 16491 41003
rect 16445 40931 16451 40965
rect 16485 40931 16491 40965
rect 16445 40893 16491 40931
rect 16445 40859 16451 40893
rect 16485 40859 16491 40893
rect 16445 40821 16491 40859
rect 16445 40787 16451 40821
rect 16485 40787 16491 40821
rect 16445 40749 16491 40787
rect 16445 40715 16451 40749
rect 16485 40715 16491 40749
rect 16445 40677 16491 40715
rect 16445 40643 16451 40677
rect 16485 40643 16491 40677
rect 16445 40605 16491 40643
rect 16445 40571 16451 40605
rect 16485 40571 16491 40605
rect 16445 40533 16491 40571
rect 16445 40499 16451 40533
rect 16485 40499 16491 40533
rect 16445 40461 16491 40499
rect 16445 40427 16451 40461
rect 16485 40427 16491 40461
rect 16445 40389 16491 40427
rect 16445 40355 16451 40389
rect 16485 40355 16491 40389
rect 16445 40317 16491 40355
rect 16445 40283 16451 40317
rect 16485 40283 16491 40317
rect 16445 40245 16491 40283
rect 16445 40211 16451 40245
rect 16485 40211 16491 40245
rect 16445 40173 16491 40211
rect 16445 40139 16451 40173
rect 16485 40139 16491 40173
rect 16445 40101 16491 40139
rect 16445 40067 16451 40101
rect 16485 40067 16491 40101
rect 16445 40029 16491 40067
rect 16445 39995 16451 40029
rect 16485 39995 16491 40029
rect 16445 39957 16491 39995
rect 16445 39923 16451 39957
rect 16485 39923 16491 39957
rect 16445 39907 16491 39923
rect 16903 41181 16949 41197
rect 16903 41147 16909 41181
rect 16943 41147 16949 41181
rect 16903 41109 16949 41147
rect 16903 41075 16909 41109
rect 16943 41075 16949 41109
rect 16903 41037 16949 41075
rect 16903 41003 16909 41037
rect 16943 41003 16949 41037
rect 16903 40965 16949 41003
rect 16903 40931 16909 40965
rect 16943 40931 16949 40965
rect 16903 40893 16949 40931
rect 16903 40859 16909 40893
rect 16943 40859 16949 40893
rect 16903 40821 16949 40859
rect 16903 40787 16909 40821
rect 16943 40787 16949 40821
rect 16903 40749 16949 40787
rect 16903 40715 16909 40749
rect 16943 40715 16949 40749
rect 16903 40677 16949 40715
rect 16903 40643 16909 40677
rect 16943 40643 16949 40677
rect 16903 40605 16949 40643
rect 16903 40571 16909 40605
rect 16943 40571 16949 40605
rect 16903 40533 16949 40571
rect 16903 40499 16909 40533
rect 16943 40499 16949 40533
rect 16903 40461 16949 40499
rect 16903 40427 16909 40461
rect 16943 40427 16949 40461
rect 16903 40389 16949 40427
rect 16903 40355 16909 40389
rect 16943 40355 16949 40389
rect 16903 40317 16949 40355
rect 16903 40283 16909 40317
rect 16943 40283 16949 40317
rect 16903 40245 16949 40283
rect 16903 40211 16909 40245
rect 16943 40211 16949 40245
rect 16903 40173 16949 40211
rect 16903 40139 16909 40173
rect 16943 40139 16949 40173
rect 16903 40101 16949 40139
rect 16903 40067 16909 40101
rect 16943 40067 16949 40101
rect 16903 40029 16949 40067
rect 16903 39995 16909 40029
rect 16943 39995 16949 40029
rect 16903 39957 16949 39995
rect 16903 39923 16909 39957
rect 16943 39923 16949 39957
rect 16903 39907 16949 39923
rect 17361 41181 17407 41197
rect 17361 41147 17367 41181
rect 17401 41147 17407 41181
rect 17361 41109 17407 41147
rect 17361 41075 17367 41109
rect 17401 41075 17407 41109
rect 17361 41037 17407 41075
rect 17361 41003 17367 41037
rect 17401 41003 17407 41037
rect 17361 40965 17407 41003
rect 17361 40931 17367 40965
rect 17401 40931 17407 40965
rect 17361 40893 17407 40931
rect 17361 40859 17367 40893
rect 17401 40859 17407 40893
rect 17361 40821 17407 40859
rect 17361 40787 17367 40821
rect 17401 40787 17407 40821
rect 17361 40749 17407 40787
rect 17361 40715 17367 40749
rect 17401 40715 17407 40749
rect 17361 40677 17407 40715
rect 17361 40643 17367 40677
rect 17401 40643 17407 40677
rect 17361 40605 17407 40643
rect 17361 40571 17367 40605
rect 17401 40571 17407 40605
rect 17361 40533 17407 40571
rect 17361 40499 17367 40533
rect 17401 40499 17407 40533
rect 17361 40461 17407 40499
rect 17361 40427 17367 40461
rect 17401 40427 17407 40461
rect 17361 40389 17407 40427
rect 17361 40355 17367 40389
rect 17401 40355 17407 40389
rect 17361 40317 17407 40355
rect 17361 40283 17367 40317
rect 17401 40283 17407 40317
rect 17361 40245 17407 40283
rect 17361 40211 17367 40245
rect 17401 40211 17407 40245
rect 17361 40173 17407 40211
rect 17361 40139 17367 40173
rect 17401 40139 17407 40173
rect 17361 40101 17407 40139
rect 17361 40067 17367 40101
rect 17401 40067 17407 40101
rect 17361 40029 17407 40067
rect 17361 39995 17367 40029
rect 17401 39995 17407 40029
rect 17361 39957 17407 39995
rect 17361 39923 17367 39957
rect 17401 39923 17407 39957
rect 17361 39907 17407 39923
rect 17819 41181 17865 41197
rect 17819 41147 17825 41181
rect 17859 41147 17865 41181
rect 17819 41109 17865 41147
rect 17819 41075 17825 41109
rect 17859 41075 17865 41109
rect 17819 41037 17865 41075
rect 17819 41003 17825 41037
rect 17859 41003 17865 41037
rect 17819 40965 17865 41003
rect 17819 40931 17825 40965
rect 17859 40931 17865 40965
rect 17819 40893 17865 40931
rect 17819 40859 17825 40893
rect 17859 40859 17865 40893
rect 17819 40821 17865 40859
rect 17819 40787 17825 40821
rect 17859 40787 17865 40821
rect 17819 40749 17865 40787
rect 17819 40715 17825 40749
rect 17859 40715 17865 40749
rect 17819 40677 17865 40715
rect 17819 40643 17825 40677
rect 17859 40643 17865 40677
rect 17819 40605 17865 40643
rect 17819 40571 17825 40605
rect 17859 40571 17865 40605
rect 17819 40533 17865 40571
rect 17819 40499 17825 40533
rect 17859 40499 17865 40533
rect 17819 40461 17865 40499
rect 17819 40427 17825 40461
rect 17859 40427 17865 40461
rect 17819 40389 17865 40427
rect 17819 40355 17825 40389
rect 17859 40355 17865 40389
rect 17819 40317 17865 40355
rect 17819 40283 17825 40317
rect 17859 40283 17865 40317
rect 17819 40245 17865 40283
rect 17819 40211 17825 40245
rect 17859 40211 17865 40245
rect 17819 40173 17865 40211
rect 17819 40139 17825 40173
rect 17859 40139 17865 40173
rect 17819 40101 17865 40139
rect 17819 40067 17825 40101
rect 17859 40067 17865 40101
rect 17819 40029 17865 40067
rect 17819 39995 17825 40029
rect 17859 39995 17865 40029
rect 17819 39957 17865 39995
rect 17819 39923 17825 39957
rect 17859 39923 17865 39957
rect 17819 39907 17865 39923
rect 18277 41181 18323 41197
rect 18277 41147 18283 41181
rect 18317 41147 18323 41181
rect 18277 41109 18323 41147
rect 18277 41075 18283 41109
rect 18317 41075 18323 41109
rect 18277 41037 18323 41075
rect 18277 41003 18283 41037
rect 18317 41003 18323 41037
rect 18277 40965 18323 41003
rect 18277 40931 18283 40965
rect 18317 40931 18323 40965
rect 18277 40893 18323 40931
rect 18277 40859 18283 40893
rect 18317 40859 18323 40893
rect 18277 40821 18323 40859
rect 18277 40787 18283 40821
rect 18317 40787 18323 40821
rect 18277 40749 18323 40787
rect 18277 40715 18283 40749
rect 18317 40715 18323 40749
rect 18277 40677 18323 40715
rect 18277 40643 18283 40677
rect 18317 40643 18323 40677
rect 18277 40605 18323 40643
rect 18277 40571 18283 40605
rect 18317 40571 18323 40605
rect 18277 40533 18323 40571
rect 18277 40499 18283 40533
rect 18317 40499 18323 40533
rect 18277 40461 18323 40499
rect 18277 40427 18283 40461
rect 18317 40427 18323 40461
rect 18277 40389 18323 40427
rect 18277 40355 18283 40389
rect 18317 40355 18323 40389
rect 18277 40317 18323 40355
rect 18277 40283 18283 40317
rect 18317 40283 18323 40317
rect 18277 40245 18323 40283
rect 18277 40211 18283 40245
rect 18317 40211 18323 40245
rect 18277 40173 18323 40211
rect 18277 40139 18283 40173
rect 18317 40139 18323 40173
rect 18277 40101 18323 40139
rect 18277 40067 18283 40101
rect 18317 40067 18323 40101
rect 18277 40029 18323 40067
rect 18277 39995 18283 40029
rect 18317 39995 18323 40029
rect 18277 39957 18323 39995
rect 18277 39923 18283 39957
rect 18317 39923 18323 39957
rect 18277 39907 18323 39923
rect 18735 41181 18781 41197
rect 18735 41147 18741 41181
rect 18775 41147 18781 41181
rect 18735 41109 18781 41147
rect 18735 41075 18741 41109
rect 18775 41075 18781 41109
rect 18735 41037 18781 41075
rect 18735 41003 18741 41037
rect 18775 41003 18781 41037
rect 18735 40965 18781 41003
rect 18735 40931 18741 40965
rect 18775 40931 18781 40965
rect 18735 40893 18781 40931
rect 18735 40859 18741 40893
rect 18775 40859 18781 40893
rect 18735 40821 18781 40859
rect 18735 40787 18741 40821
rect 18775 40787 18781 40821
rect 18735 40749 18781 40787
rect 18735 40715 18741 40749
rect 18775 40715 18781 40749
rect 18735 40677 18781 40715
rect 18735 40643 18741 40677
rect 18775 40643 18781 40677
rect 18735 40605 18781 40643
rect 18735 40571 18741 40605
rect 18775 40571 18781 40605
rect 18735 40533 18781 40571
rect 18735 40499 18741 40533
rect 18775 40499 18781 40533
rect 18735 40461 18781 40499
rect 18735 40427 18741 40461
rect 18775 40427 18781 40461
rect 18735 40389 18781 40427
rect 18735 40355 18741 40389
rect 18775 40355 18781 40389
rect 18735 40317 18781 40355
rect 18735 40283 18741 40317
rect 18775 40283 18781 40317
rect 18735 40245 18781 40283
rect 18735 40211 18741 40245
rect 18775 40211 18781 40245
rect 18735 40173 18781 40211
rect 18735 40139 18741 40173
rect 18775 40139 18781 40173
rect 18735 40101 18781 40139
rect 18735 40067 18741 40101
rect 18775 40067 18781 40101
rect 18735 40029 18781 40067
rect 18735 39995 18741 40029
rect 18775 39995 18781 40029
rect 18735 39957 18781 39995
rect 18735 39923 18741 39957
rect 18775 39923 18781 39957
rect 18735 39907 18781 39923
rect 19193 41181 19239 41197
rect 19193 41147 19199 41181
rect 19233 41147 19239 41181
rect 19193 41109 19239 41147
rect 19193 41075 19199 41109
rect 19233 41075 19239 41109
rect 19193 41037 19239 41075
rect 19193 41003 19199 41037
rect 19233 41003 19239 41037
rect 19193 40965 19239 41003
rect 19193 40931 19199 40965
rect 19233 40931 19239 40965
rect 19193 40893 19239 40931
rect 19193 40859 19199 40893
rect 19233 40859 19239 40893
rect 19193 40821 19239 40859
rect 19193 40787 19199 40821
rect 19233 40787 19239 40821
rect 19193 40749 19239 40787
rect 19193 40715 19199 40749
rect 19233 40715 19239 40749
rect 19193 40677 19239 40715
rect 19193 40643 19199 40677
rect 19233 40643 19239 40677
rect 19193 40605 19239 40643
rect 19193 40571 19199 40605
rect 19233 40571 19239 40605
rect 19193 40533 19239 40571
rect 19193 40499 19199 40533
rect 19233 40499 19239 40533
rect 19193 40461 19239 40499
rect 19193 40427 19199 40461
rect 19233 40427 19239 40461
rect 19193 40389 19239 40427
rect 19193 40355 19199 40389
rect 19233 40355 19239 40389
rect 19193 40317 19239 40355
rect 19193 40283 19199 40317
rect 19233 40283 19239 40317
rect 19193 40245 19239 40283
rect 19193 40211 19199 40245
rect 19233 40211 19239 40245
rect 19193 40173 19239 40211
rect 19193 40139 19199 40173
rect 19233 40139 19239 40173
rect 19193 40101 19239 40139
rect 19193 40067 19199 40101
rect 19233 40067 19239 40101
rect 19193 40029 19239 40067
rect 19193 39995 19199 40029
rect 19233 39995 19239 40029
rect 19193 39957 19239 39995
rect 19193 39923 19199 39957
rect 19233 39923 19239 39957
rect 19193 39907 19239 39923
rect 19651 41181 19697 41197
rect 19651 41147 19657 41181
rect 19691 41147 19697 41181
rect 19651 41109 19697 41147
rect 19651 41075 19657 41109
rect 19691 41075 19697 41109
rect 19651 41037 19697 41075
rect 19651 41003 19657 41037
rect 19691 41003 19697 41037
rect 19651 40965 19697 41003
rect 19651 40931 19657 40965
rect 19691 40931 19697 40965
rect 19651 40893 19697 40931
rect 19651 40859 19657 40893
rect 19691 40859 19697 40893
rect 19651 40821 19697 40859
rect 19651 40787 19657 40821
rect 19691 40787 19697 40821
rect 19651 40749 19697 40787
rect 19651 40715 19657 40749
rect 19691 40715 19697 40749
rect 19651 40677 19697 40715
rect 19651 40643 19657 40677
rect 19691 40643 19697 40677
rect 19651 40605 19697 40643
rect 19651 40571 19657 40605
rect 19691 40571 19697 40605
rect 19651 40533 19697 40571
rect 19651 40499 19657 40533
rect 19691 40499 19697 40533
rect 19651 40461 19697 40499
rect 19651 40427 19657 40461
rect 19691 40427 19697 40461
rect 19651 40389 19697 40427
rect 19651 40355 19657 40389
rect 19691 40355 19697 40389
rect 19651 40317 19697 40355
rect 19651 40283 19657 40317
rect 19691 40283 19697 40317
rect 19651 40245 19697 40283
rect 19651 40211 19657 40245
rect 19691 40211 19697 40245
rect 19651 40173 19697 40211
rect 19651 40139 19657 40173
rect 19691 40139 19697 40173
rect 19651 40101 19697 40139
rect 19651 40067 19657 40101
rect 19691 40067 19697 40101
rect 19651 40029 19697 40067
rect 19651 39995 19657 40029
rect 19691 39995 19697 40029
rect 19651 39957 19697 39995
rect 19651 39923 19657 39957
rect 19691 39923 19697 39957
rect 19651 39907 19697 39923
rect 20109 41181 20155 41197
rect 20109 41147 20115 41181
rect 20149 41147 20155 41181
rect 20109 41109 20155 41147
rect 20109 41075 20115 41109
rect 20149 41075 20155 41109
rect 20109 41037 20155 41075
rect 20109 41003 20115 41037
rect 20149 41003 20155 41037
rect 20109 40965 20155 41003
rect 20109 40931 20115 40965
rect 20149 40931 20155 40965
rect 20109 40893 20155 40931
rect 20109 40859 20115 40893
rect 20149 40859 20155 40893
rect 20109 40821 20155 40859
rect 20109 40787 20115 40821
rect 20149 40787 20155 40821
rect 20109 40749 20155 40787
rect 20109 40715 20115 40749
rect 20149 40715 20155 40749
rect 20109 40677 20155 40715
rect 20109 40643 20115 40677
rect 20149 40643 20155 40677
rect 20109 40605 20155 40643
rect 20109 40571 20115 40605
rect 20149 40571 20155 40605
rect 20109 40533 20155 40571
rect 20109 40499 20115 40533
rect 20149 40499 20155 40533
rect 20109 40461 20155 40499
rect 20109 40427 20115 40461
rect 20149 40427 20155 40461
rect 20109 40389 20155 40427
rect 20109 40355 20115 40389
rect 20149 40355 20155 40389
rect 20109 40317 20155 40355
rect 20109 40283 20115 40317
rect 20149 40283 20155 40317
rect 20109 40245 20155 40283
rect 20109 40211 20115 40245
rect 20149 40211 20155 40245
rect 20109 40173 20155 40211
rect 20109 40139 20115 40173
rect 20149 40139 20155 40173
rect 20109 40101 20155 40139
rect 20109 40067 20115 40101
rect 20149 40067 20155 40101
rect 20109 40029 20155 40067
rect 20109 39995 20115 40029
rect 20149 39995 20155 40029
rect 20109 39957 20155 39995
rect 20109 39923 20115 39957
rect 20149 39923 20155 39957
rect 20109 39907 20155 39923
rect 20567 41181 20613 41197
rect 20567 41147 20573 41181
rect 20607 41147 20613 41181
rect 20567 41109 20613 41147
rect 20567 41075 20573 41109
rect 20607 41075 20613 41109
rect 20567 41037 20613 41075
rect 20567 41003 20573 41037
rect 20607 41003 20613 41037
rect 20567 40965 20613 41003
rect 20567 40931 20573 40965
rect 20607 40931 20613 40965
rect 20567 40893 20613 40931
rect 20567 40859 20573 40893
rect 20607 40859 20613 40893
rect 20567 40821 20613 40859
rect 20567 40787 20573 40821
rect 20607 40787 20613 40821
rect 20567 40749 20613 40787
rect 20567 40715 20573 40749
rect 20607 40715 20613 40749
rect 20567 40677 20613 40715
rect 20567 40643 20573 40677
rect 20607 40643 20613 40677
rect 20567 40605 20613 40643
rect 20567 40571 20573 40605
rect 20607 40571 20613 40605
rect 20567 40533 20613 40571
rect 20567 40499 20573 40533
rect 20607 40499 20613 40533
rect 20567 40461 20613 40499
rect 20567 40427 20573 40461
rect 20607 40427 20613 40461
rect 20567 40389 20613 40427
rect 20567 40355 20573 40389
rect 20607 40355 20613 40389
rect 20567 40317 20613 40355
rect 20567 40283 20573 40317
rect 20607 40283 20613 40317
rect 20567 40245 20613 40283
rect 20567 40211 20573 40245
rect 20607 40211 20613 40245
rect 20567 40173 20613 40211
rect 20567 40139 20573 40173
rect 20607 40139 20613 40173
rect 20567 40101 20613 40139
rect 20567 40067 20573 40101
rect 20607 40067 20613 40101
rect 20567 40029 20613 40067
rect 20567 39995 20573 40029
rect 20607 39995 20613 40029
rect 20567 39957 20613 39995
rect 20567 39923 20573 39957
rect 20607 39923 20613 39957
rect 20567 39907 20613 39923
rect 21025 41181 21071 41197
rect 21025 41147 21031 41181
rect 21065 41147 21071 41181
rect 21025 41109 21071 41147
rect 21025 41075 21031 41109
rect 21065 41075 21071 41109
rect 21025 41037 21071 41075
rect 21025 41003 21031 41037
rect 21065 41003 21071 41037
rect 21025 40965 21071 41003
rect 21025 40931 21031 40965
rect 21065 40931 21071 40965
rect 21025 40893 21071 40931
rect 21025 40859 21031 40893
rect 21065 40859 21071 40893
rect 21025 40821 21071 40859
rect 21025 40787 21031 40821
rect 21065 40787 21071 40821
rect 21025 40749 21071 40787
rect 21025 40715 21031 40749
rect 21065 40715 21071 40749
rect 21025 40677 21071 40715
rect 21025 40643 21031 40677
rect 21065 40643 21071 40677
rect 21025 40605 21071 40643
rect 21025 40571 21031 40605
rect 21065 40571 21071 40605
rect 21025 40533 21071 40571
rect 21025 40499 21031 40533
rect 21065 40499 21071 40533
rect 21025 40461 21071 40499
rect 21025 40427 21031 40461
rect 21065 40427 21071 40461
rect 21025 40389 21071 40427
rect 21025 40355 21031 40389
rect 21065 40355 21071 40389
rect 21025 40317 21071 40355
rect 21025 40283 21031 40317
rect 21065 40283 21071 40317
rect 21025 40245 21071 40283
rect 21025 40211 21031 40245
rect 21065 40211 21071 40245
rect 21025 40173 21071 40211
rect 21025 40139 21031 40173
rect 21065 40139 21071 40173
rect 21025 40101 21071 40139
rect 21025 40067 21031 40101
rect 21065 40067 21071 40101
rect 21025 40029 21071 40067
rect 21025 39995 21031 40029
rect 21065 39995 21071 40029
rect 21025 39957 21071 39995
rect 21025 39923 21031 39957
rect 21065 39923 21071 39957
rect 21025 39907 21071 39923
rect 21483 41181 21529 41197
rect 21483 41147 21489 41181
rect 21523 41147 21529 41181
rect 21483 41109 21529 41147
rect 21483 41075 21489 41109
rect 21523 41075 21529 41109
rect 21483 41037 21529 41075
rect 21483 41003 21489 41037
rect 21523 41003 21529 41037
rect 21483 40965 21529 41003
rect 21483 40931 21489 40965
rect 21523 40931 21529 40965
rect 21483 40893 21529 40931
rect 21483 40859 21489 40893
rect 21523 40859 21529 40893
rect 21483 40821 21529 40859
rect 21483 40787 21489 40821
rect 21523 40787 21529 40821
rect 21483 40749 21529 40787
rect 21483 40715 21489 40749
rect 21523 40715 21529 40749
rect 21483 40677 21529 40715
rect 21483 40643 21489 40677
rect 21523 40643 21529 40677
rect 21483 40605 21529 40643
rect 21483 40571 21489 40605
rect 21523 40571 21529 40605
rect 21483 40533 21529 40571
rect 21483 40499 21489 40533
rect 21523 40499 21529 40533
rect 21483 40461 21529 40499
rect 21483 40427 21489 40461
rect 21523 40427 21529 40461
rect 21483 40389 21529 40427
rect 21483 40355 21489 40389
rect 21523 40355 21529 40389
rect 21483 40317 21529 40355
rect 21483 40283 21489 40317
rect 21523 40283 21529 40317
rect 21483 40245 21529 40283
rect 21483 40211 21489 40245
rect 21523 40211 21529 40245
rect 21483 40173 21529 40211
rect 21483 40139 21489 40173
rect 21523 40139 21529 40173
rect 21483 40101 21529 40139
rect 21483 40067 21489 40101
rect 21523 40067 21529 40101
rect 21483 40029 21529 40067
rect 21483 39995 21489 40029
rect 21523 39995 21529 40029
rect 21483 39957 21529 39995
rect 21483 39923 21489 39957
rect 21523 39923 21529 39957
rect 21483 39907 21529 39923
rect 21941 41181 21987 41197
rect 21941 41147 21947 41181
rect 21981 41147 21987 41181
rect 21941 41109 21987 41147
rect 21941 41075 21947 41109
rect 21981 41075 21987 41109
rect 21941 41037 21987 41075
rect 21941 41003 21947 41037
rect 21981 41003 21987 41037
rect 21941 40965 21987 41003
rect 21941 40931 21947 40965
rect 21981 40931 21987 40965
rect 21941 40893 21987 40931
rect 21941 40859 21947 40893
rect 21981 40859 21987 40893
rect 21941 40821 21987 40859
rect 21941 40787 21947 40821
rect 21981 40787 21987 40821
rect 21941 40749 21987 40787
rect 21941 40715 21947 40749
rect 21981 40715 21987 40749
rect 21941 40677 21987 40715
rect 21941 40643 21947 40677
rect 21981 40643 21987 40677
rect 21941 40605 21987 40643
rect 21941 40571 21947 40605
rect 21981 40571 21987 40605
rect 21941 40533 21987 40571
rect 21941 40499 21947 40533
rect 21981 40499 21987 40533
rect 21941 40461 21987 40499
rect 21941 40427 21947 40461
rect 21981 40427 21987 40461
rect 21941 40389 21987 40427
rect 21941 40355 21947 40389
rect 21981 40355 21987 40389
rect 21941 40317 21987 40355
rect 21941 40283 21947 40317
rect 21981 40283 21987 40317
rect 21941 40245 21987 40283
rect 21941 40211 21947 40245
rect 21981 40211 21987 40245
rect 21941 40173 21987 40211
rect 21941 40139 21947 40173
rect 21981 40139 21987 40173
rect 21941 40101 21987 40139
rect 21941 40067 21947 40101
rect 21981 40067 21987 40101
rect 21941 40029 21987 40067
rect 21941 39995 21947 40029
rect 21981 39995 21987 40029
rect 21941 39957 21987 39995
rect 21941 39923 21947 39957
rect 21981 39923 21987 39957
rect 21941 39907 21987 39923
rect 22399 41181 22445 41197
rect 22399 41147 22405 41181
rect 22439 41147 22445 41181
rect 22399 41109 22445 41147
rect 22399 41075 22405 41109
rect 22439 41075 22445 41109
rect 22399 41037 22445 41075
rect 22399 41003 22405 41037
rect 22439 41003 22445 41037
rect 22399 40965 22445 41003
rect 22399 40931 22405 40965
rect 22439 40931 22445 40965
rect 22399 40893 22445 40931
rect 22399 40859 22405 40893
rect 22439 40859 22445 40893
rect 22399 40821 22445 40859
rect 22399 40787 22405 40821
rect 22439 40787 22445 40821
rect 22399 40749 22445 40787
rect 22399 40715 22405 40749
rect 22439 40715 22445 40749
rect 22399 40677 22445 40715
rect 22399 40643 22405 40677
rect 22439 40643 22445 40677
rect 22399 40605 22445 40643
rect 22399 40571 22405 40605
rect 22439 40571 22445 40605
rect 22399 40533 22445 40571
rect 22399 40499 22405 40533
rect 22439 40499 22445 40533
rect 22399 40461 22445 40499
rect 22399 40427 22405 40461
rect 22439 40427 22445 40461
rect 22399 40389 22445 40427
rect 22399 40355 22405 40389
rect 22439 40355 22445 40389
rect 22399 40317 22445 40355
rect 22399 40283 22405 40317
rect 22439 40283 22445 40317
rect 22399 40245 22445 40283
rect 22399 40211 22405 40245
rect 22439 40211 22445 40245
rect 22399 40173 22445 40211
rect 22399 40139 22405 40173
rect 22439 40139 22445 40173
rect 22399 40101 22445 40139
rect 22399 40067 22405 40101
rect 22439 40067 22445 40101
rect 22399 40029 22445 40067
rect 22399 39995 22405 40029
rect 22439 39995 22445 40029
rect 22399 39957 22445 39995
rect 22399 39923 22405 39957
rect 22439 39923 22445 39957
rect 22399 39907 22445 39923
rect 22857 41181 22903 41197
rect 22857 41147 22863 41181
rect 22897 41147 22903 41181
rect 22857 41109 22903 41147
rect 22857 41075 22863 41109
rect 22897 41075 22903 41109
rect 22857 41037 22903 41075
rect 22857 41003 22863 41037
rect 22897 41003 22903 41037
rect 22857 40965 22903 41003
rect 22857 40931 22863 40965
rect 22897 40931 22903 40965
rect 22857 40893 22903 40931
rect 22857 40859 22863 40893
rect 22897 40859 22903 40893
rect 22857 40821 22903 40859
rect 22857 40787 22863 40821
rect 22897 40787 22903 40821
rect 22857 40749 22903 40787
rect 22857 40715 22863 40749
rect 22897 40715 22903 40749
rect 22857 40677 22903 40715
rect 22857 40643 22863 40677
rect 22897 40643 22903 40677
rect 22857 40605 22903 40643
rect 22857 40571 22863 40605
rect 22897 40571 22903 40605
rect 22857 40533 22903 40571
rect 22857 40499 22863 40533
rect 22897 40499 22903 40533
rect 22857 40461 22903 40499
rect 22857 40427 22863 40461
rect 22897 40427 22903 40461
rect 22857 40389 22903 40427
rect 22857 40355 22863 40389
rect 22897 40355 22903 40389
rect 22857 40317 22903 40355
rect 22857 40283 22863 40317
rect 22897 40283 22903 40317
rect 22857 40245 22903 40283
rect 22857 40211 22863 40245
rect 22897 40211 22903 40245
rect 22857 40173 22903 40211
rect 22857 40139 22863 40173
rect 22897 40139 22903 40173
rect 22857 40101 22903 40139
rect 22857 40067 22863 40101
rect 22897 40067 22903 40101
rect 22857 40029 22903 40067
rect 22857 39995 22863 40029
rect 22897 39995 22903 40029
rect 22857 39957 22903 39995
rect 22857 39923 22863 39957
rect 22897 39923 22903 39957
rect 22857 39907 22903 39923
rect 23315 41181 23361 41197
rect 23315 41147 23321 41181
rect 23355 41147 23361 41181
rect 23315 41109 23361 41147
rect 23315 41075 23321 41109
rect 23355 41075 23361 41109
rect 23315 41037 23361 41075
rect 23315 41003 23321 41037
rect 23355 41003 23361 41037
rect 23315 40965 23361 41003
rect 23315 40931 23321 40965
rect 23355 40931 23361 40965
rect 23315 40893 23361 40931
rect 23315 40859 23321 40893
rect 23355 40859 23361 40893
rect 23315 40821 23361 40859
rect 23315 40787 23321 40821
rect 23355 40787 23361 40821
rect 23315 40749 23361 40787
rect 23315 40715 23321 40749
rect 23355 40715 23361 40749
rect 23315 40677 23361 40715
rect 23315 40643 23321 40677
rect 23355 40643 23361 40677
rect 23315 40605 23361 40643
rect 23315 40571 23321 40605
rect 23355 40571 23361 40605
rect 23315 40533 23361 40571
rect 23315 40499 23321 40533
rect 23355 40499 23361 40533
rect 23315 40461 23361 40499
rect 23315 40427 23321 40461
rect 23355 40427 23361 40461
rect 23315 40389 23361 40427
rect 23315 40355 23321 40389
rect 23355 40355 23361 40389
rect 23315 40317 23361 40355
rect 23315 40283 23321 40317
rect 23355 40283 23361 40317
rect 23315 40245 23361 40283
rect 23315 40211 23321 40245
rect 23355 40211 23361 40245
rect 23315 40173 23361 40211
rect 23315 40139 23321 40173
rect 23355 40139 23361 40173
rect 23315 40101 23361 40139
rect 23315 40067 23321 40101
rect 23355 40067 23361 40101
rect 23315 40029 23361 40067
rect 23315 39995 23321 40029
rect 23355 39995 23361 40029
rect 23315 39957 23361 39995
rect 23315 39923 23321 39957
rect 23355 39923 23361 39957
rect 23315 39907 23361 39923
rect 23773 41181 23819 41197
rect 23773 41147 23779 41181
rect 23813 41147 23819 41181
rect 23773 41109 23819 41147
rect 23773 41075 23779 41109
rect 23813 41075 23819 41109
rect 23773 41037 23819 41075
rect 23773 41003 23779 41037
rect 23813 41003 23819 41037
rect 23773 40965 23819 41003
rect 23773 40931 23779 40965
rect 23813 40931 23819 40965
rect 23773 40893 23819 40931
rect 23773 40859 23779 40893
rect 23813 40859 23819 40893
rect 23773 40821 23819 40859
rect 23773 40787 23779 40821
rect 23813 40787 23819 40821
rect 23773 40749 23819 40787
rect 23773 40715 23779 40749
rect 23813 40715 23819 40749
rect 23773 40677 23819 40715
rect 23773 40643 23779 40677
rect 23813 40643 23819 40677
rect 23773 40605 23819 40643
rect 23773 40571 23779 40605
rect 23813 40571 23819 40605
rect 23773 40533 23819 40571
rect 23773 40499 23779 40533
rect 23813 40499 23819 40533
rect 23773 40461 23819 40499
rect 23773 40427 23779 40461
rect 23813 40427 23819 40461
rect 23773 40389 23819 40427
rect 23773 40355 23779 40389
rect 23813 40355 23819 40389
rect 23773 40317 23819 40355
rect 23773 40283 23779 40317
rect 23813 40283 23819 40317
rect 23773 40245 23819 40283
rect 23773 40211 23779 40245
rect 23813 40211 23819 40245
rect 23773 40173 23819 40211
rect 23773 40139 23779 40173
rect 23813 40139 23819 40173
rect 23773 40101 23819 40139
rect 23773 40067 23779 40101
rect 23813 40067 23819 40101
rect 23773 40029 23819 40067
rect 23773 39995 23779 40029
rect 23813 39995 23819 40029
rect 23773 39957 23819 39995
rect 23773 39923 23779 39957
rect 23813 39923 23819 39957
rect 23773 39907 23819 39923
rect 24231 41181 24277 41197
rect 24231 41147 24237 41181
rect 24271 41147 24277 41181
rect 24231 41109 24277 41147
rect 24231 41075 24237 41109
rect 24271 41075 24277 41109
rect 24231 41037 24277 41075
rect 24231 41003 24237 41037
rect 24271 41003 24277 41037
rect 24231 40965 24277 41003
rect 24231 40931 24237 40965
rect 24271 40931 24277 40965
rect 24231 40893 24277 40931
rect 24231 40859 24237 40893
rect 24271 40859 24277 40893
rect 24231 40821 24277 40859
rect 24231 40787 24237 40821
rect 24271 40787 24277 40821
rect 24231 40749 24277 40787
rect 24231 40715 24237 40749
rect 24271 40715 24277 40749
rect 24231 40677 24277 40715
rect 24231 40643 24237 40677
rect 24271 40643 24277 40677
rect 24231 40605 24277 40643
rect 24231 40571 24237 40605
rect 24271 40571 24277 40605
rect 24231 40533 24277 40571
rect 24231 40499 24237 40533
rect 24271 40499 24277 40533
rect 24231 40461 24277 40499
rect 24231 40427 24237 40461
rect 24271 40427 24277 40461
rect 24231 40389 24277 40427
rect 24231 40355 24237 40389
rect 24271 40355 24277 40389
rect 24231 40317 24277 40355
rect 24231 40283 24237 40317
rect 24271 40283 24277 40317
rect 24231 40245 24277 40283
rect 24231 40211 24237 40245
rect 24271 40211 24277 40245
rect 24231 40173 24277 40211
rect 24231 40139 24237 40173
rect 24271 40139 24277 40173
rect 24231 40101 24277 40139
rect 24231 40067 24237 40101
rect 24271 40067 24277 40101
rect 24231 40029 24277 40067
rect 24231 39995 24237 40029
rect 24271 39995 24277 40029
rect 24231 39957 24277 39995
rect 24231 39923 24237 39957
rect 24271 39923 24277 39957
rect 24231 39907 24277 39923
rect 24689 41181 24735 41197
rect 24689 41147 24695 41181
rect 24729 41147 24735 41181
rect 24689 41109 24735 41147
rect 24689 41075 24695 41109
rect 24729 41075 24735 41109
rect 24689 41037 24735 41075
rect 24689 41003 24695 41037
rect 24729 41003 24735 41037
rect 24689 40965 24735 41003
rect 24689 40931 24695 40965
rect 24729 40931 24735 40965
rect 24689 40893 24735 40931
rect 24689 40859 24695 40893
rect 24729 40859 24735 40893
rect 24689 40821 24735 40859
rect 24689 40787 24695 40821
rect 24729 40787 24735 40821
rect 24689 40749 24735 40787
rect 24689 40715 24695 40749
rect 24729 40715 24735 40749
rect 24689 40677 24735 40715
rect 24689 40643 24695 40677
rect 24729 40643 24735 40677
rect 24689 40605 24735 40643
rect 24689 40571 24695 40605
rect 24729 40571 24735 40605
rect 24689 40533 24735 40571
rect 24689 40499 24695 40533
rect 24729 40499 24735 40533
rect 24689 40461 24735 40499
rect 24689 40427 24695 40461
rect 24729 40427 24735 40461
rect 24689 40389 24735 40427
rect 24689 40355 24695 40389
rect 24729 40355 24735 40389
rect 24689 40317 24735 40355
rect 24689 40283 24695 40317
rect 24729 40283 24735 40317
rect 24689 40245 24735 40283
rect 24689 40211 24695 40245
rect 24729 40211 24735 40245
rect 24689 40173 24735 40211
rect 24689 40139 24695 40173
rect 24729 40139 24735 40173
rect 24689 40101 24735 40139
rect 24689 40067 24695 40101
rect 24729 40067 24735 40101
rect 24689 40029 24735 40067
rect 24689 39995 24695 40029
rect 24729 39995 24735 40029
rect 24689 39957 24735 39995
rect 24689 39923 24695 39957
rect 24729 39923 24735 39957
rect 24689 39907 24735 39923
rect 25147 41181 25193 41197
rect 25147 41147 25153 41181
rect 25187 41147 25193 41181
rect 25147 41109 25193 41147
rect 25147 41075 25153 41109
rect 25187 41075 25193 41109
rect 25147 41037 25193 41075
rect 25147 41003 25153 41037
rect 25187 41003 25193 41037
rect 25147 40965 25193 41003
rect 25147 40931 25153 40965
rect 25187 40931 25193 40965
rect 25147 40893 25193 40931
rect 25147 40859 25153 40893
rect 25187 40859 25193 40893
rect 25147 40821 25193 40859
rect 25147 40787 25153 40821
rect 25187 40787 25193 40821
rect 25147 40749 25193 40787
rect 25147 40715 25153 40749
rect 25187 40715 25193 40749
rect 25147 40677 25193 40715
rect 25147 40643 25153 40677
rect 25187 40643 25193 40677
rect 25147 40605 25193 40643
rect 25147 40571 25153 40605
rect 25187 40571 25193 40605
rect 25147 40533 25193 40571
rect 25147 40499 25153 40533
rect 25187 40499 25193 40533
rect 25147 40461 25193 40499
rect 25147 40427 25153 40461
rect 25187 40427 25193 40461
rect 25147 40389 25193 40427
rect 25147 40355 25153 40389
rect 25187 40355 25193 40389
rect 25147 40317 25193 40355
rect 25147 40283 25153 40317
rect 25187 40283 25193 40317
rect 25147 40245 25193 40283
rect 25147 40211 25153 40245
rect 25187 40211 25193 40245
rect 25147 40173 25193 40211
rect 25147 40139 25153 40173
rect 25187 40139 25193 40173
rect 25147 40101 25193 40139
rect 25147 40067 25153 40101
rect 25187 40067 25193 40101
rect 25147 40029 25193 40067
rect 25147 39995 25153 40029
rect 25187 39995 25193 40029
rect 25147 39957 25193 39995
rect 25147 39923 25153 39957
rect 25187 39923 25193 39957
rect 25147 39907 25193 39923
rect 25605 41181 25651 41197
rect 25605 41147 25611 41181
rect 25645 41147 25651 41181
rect 25605 41109 25651 41147
rect 25605 41075 25611 41109
rect 25645 41075 25651 41109
rect 25605 41037 25651 41075
rect 25605 41003 25611 41037
rect 25645 41003 25651 41037
rect 25605 40965 25651 41003
rect 25605 40931 25611 40965
rect 25645 40931 25651 40965
rect 25605 40893 25651 40931
rect 25605 40859 25611 40893
rect 25645 40859 25651 40893
rect 25605 40821 25651 40859
rect 25605 40787 25611 40821
rect 25645 40787 25651 40821
rect 25605 40749 25651 40787
rect 25605 40715 25611 40749
rect 25645 40715 25651 40749
rect 25605 40677 25651 40715
rect 25605 40643 25611 40677
rect 25645 40643 25651 40677
rect 25605 40605 25651 40643
rect 25605 40571 25611 40605
rect 25645 40571 25651 40605
rect 25605 40533 25651 40571
rect 25605 40499 25611 40533
rect 25645 40499 25651 40533
rect 25605 40461 25651 40499
rect 25605 40427 25611 40461
rect 25645 40427 25651 40461
rect 25605 40389 25651 40427
rect 25605 40355 25611 40389
rect 25645 40355 25651 40389
rect 25605 40317 25651 40355
rect 25605 40283 25611 40317
rect 25645 40283 25651 40317
rect 25605 40245 25651 40283
rect 25605 40211 25611 40245
rect 25645 40211 25651 40245
rect 25605 40173 25651 40211
rect 25605 40139 25611 40173
rect 25645 40139 25651 40173
rect 25605 40101 25651 40139
rect 25605 40067 25611 40101
rect 25645 40067 25651 40101
rect 25605 40029 25651 40067
rect 25605 39995 25611 40029
rect 25645 39995 25651 40029
rect 25605 39957 25651 39995
rect 25605 39923 25611 39957
rect 25645 39923 25651 39957
rect 25605 39907 25651 39923
rect 26063 41181 26109 41197
rect 26063 41147 26069 41181
rect 26103 41147 26109 41181
rect 26063 41109 26109 41147
rect 26063 41075 26069 41109
rect 26103 41075 26109 41109
rect 26063 41037 26109 41075
rect 26063 41003 26069 41037
rect 26103 41003 26109 41037
rect 26063 40965 26109 41003
rect 26063 40931 26069 40965
rect 26103 40931 26109 40965
rect 26063 40893 26109 40931
rect 26063 40859 26069 40893
rect 26103 40859 26109 40893
rect 26063 40821 26109 40859
rect 26063 40787 26069 40821
rect 26103 40787 26109 40821
rect 26063 40749 26109 40787
rect 26063 40715 26069 40749
rect 26103 40715 26109 40749
rect 26063 40677 26109 40715
rect 26063 40643 26069 40677
rect 26103 40643 26109 40677
rect 26063 40605 26109 40643
rect 26063 40571 26069 40605
rect 26103 40571 26109 40605
rect 26063 40533 26109 40571
rect 26063 40499 26069 40533
rect 26103 40499 26109 40533
rect 26063 40461 26109 40499
rect 26063 40427 26069 40461
rect 26103 40427 26109 40461
rect 26063 40389 26109 40427
rect 26063 40355 26069 40389
rect 26103 40355 26109 40389
rect 26063 40317 26109 40355
rect 26063 40283 26069 40317
rect 26103 40283 26109 40317
rect 26063 40245 26109 40283
rect 26063 40211 26069 40245
rect 26103 40211 26109 40245
rect 26063 40173 26109 40211
rect 26063 40139 26069 40173
rect 26103 40139 26109 40173
rect 26063 40101 26109 40139
rect 26063 40067 26069 40101
rect 26103 40067 26109 40101
rect 26063 40029 26109 40067
rect 26063 39995 26069 40029
rect 26103 39995 26109 40029
rect 26063 39957 26109 39995
rect 26063 39923 26069 39957
rect 26103 39923 26109 39957
rect 26063 39907 26109 39923
rect 26521 41181 26567 41197
rect 26521 41147 26527 41181
rect 26561 41147 26567 41181
rect 26521 41109 26567 41147
rect 26521 41075 26527 41109
rect 26561 41075 26567 41109
rect 26521 41037 26567 41075
rect 26521 41003 26527 41037
rect 26561 41003 26567 41037
rect 26521 40965 26567 41003
rect 26521 40931 26527 40965
rect 26561 40931 26567 40965
rect 26521 40893 26567 40931
rect 26521 40859 26527 40893
rect 26561 40859 26567 40893
rect 26521 40821 26567 40859
rect 26521 40787 26527 40821
rect 26561 40787 26567 40821
rect 26521 40749 26567 40787
rect 26521 40715 26527 40749
rect 26561 40715 26567 40749
rect 26521 40677 26567 40715
rect 26521 40643 26527 40677
rect 26561 40643 26567 40677
rect 26521 40605 26567 40643
rect 26521 40571 26527 40605
rect 26561 40571 26567 40605
rect 26521 40533 26567 40571
rect 26521 40499 26527 40533
rect 26561 40499 26567 40533
rect 26521 40461 26567 40499
rect 26521 40427 26527 40461
rect 26561 40427 26567 40461
rect 26521 40389 26567 40427
rect 26521 40355 26527 40389
rect 26561 40355 26567 40389
rect 26521 40317 26567 40355
rect 26521 40283 26527 40317
rect 26561 40283 26567 40317
rect 26521 40245 26567 40283
rect 26521 40211 26527 40245
rect 26561 40211 26567 40245
rect 26521 40173 26567 40211
rect 26521 40139 26527 40173
rect 26561 40139 26567 40173
rect 26521 40101 26567 40139
rect 26521 40067 26527 40101
rect 26561 40067 26567 40101
rect 26521 40029 26567 40067
rect 26521 39995 26527 40029
rect 26561 39995 26567 40029
rect 26521 39957 26567 39995
rect 26521 39923 26527 39957
rect 26561 39923 26567 39957
rect 26521 39907 26567 39923
rect 26979 41188 27025 41197
rect 27338 41188 27344 41200
rect 26979 41181 27344 41188
rect 26979 41147 26985 41181
rect 27019 41160 27344 41181
rect 27019 41147 27025 41160
rect 27338 41148 27344 41160
rect 27396 41148 27402 41200
rect 27437 41181 27483 41197
rect 26979 41109 27025 41147
rect 26979 41075 26985 41109
rect 27019 41075 27025 41109
rect 26979 41037 27025 41075
rect 26979 41003 26985 41037
rect 27019 41003 27025 41037
rect 26979 40965 27025 41003
rect 26979 40931 26985 40965
rect 27019 40931 27025 40965
rect 26979 40893 27025 40931
rect 26979 40859 26985 40893
rect 27019 40859 27025 40893
rect 26979 40821 27025 40859
rect 26979 40787 26985 40821
rect 27019 40787 27025 40821
rect 26979 40749 27025 40787
rect 26979 40715 26985 40749
rect 27019 40715 27025 40749
rect 26979 40677 27025 40715
rect 26979 40643 26985 40677
rect 27019 40643 27025 40677
rect 26979 40605 27025 40643
rect 26979 40571 26985 40605
rect 27019 40571 27025 40605
rect 26979 40533 27025 40571
rect 26979 40499 26985 40533
rect 27019 40499 27025 40533
rect 26979 40461 27025 40499
rect 26979 40427 26985 40461
rect 27019 40427 27025 40461
rect 26979 40389 27025 40427
rect 26979 40355 26985 40389
rect 27019 40355 27025 40389
rect 26979 40317 27025 40355
rect 26979 40283 26985 40317
rect 27019 40283 27025 40317
rect 26979 40245 27025 40283
rect 26979 40211 26985 40245
rect 27019 40211 27025 40245
rect 26979 40173 27025 40211
rect 26979 40139 26985 40173
rect 27019 40139 27025 40173
rect 26979 40101 27025 40139
rect 26979 40067 26985 40101
rect 27019 40067 27025 40101
rect 26979 40029 27025 40067
rect 26979 39995 26985 40029
rect 27019 39995 27025 40029
rect 26979 39957 27025 39995
rect 26979 39923 26985 39957
rect 27019 39923 27025 39957
rect 26979 39907 27025 39923
rect 27437 41147 27443 41181
rect 27477 41147 27483 41181
rect 27437 41109 27483 41147
rect 27437 41075 27443 41109
rect 27477 41075 27483 41109
rect 27437 41037 27483 41075
rect 27437 41003 27443 41037
rect 27477 41003 27483 41037
rect 27437 40965 27483 41003
rect 27437 40931 27443 40965
rect 27477 40931 27483 40965
rect 27437 40893 27483 40931
rect 27437 40859 27443 40893
rect 27477 40859 27483 40893
rect 27437 40821 27483 40859
rect 27437 40787 27443 40821
rect 27477 40787 27483 40821
rect 27437 40749 27483 40787
rect 27437 40715 27443 40749
rect 27477 40715 27483 40749
rect 27437 40677 27483 40715
rect 27437 40643 27443 40677
rect 27477 40643 27483 40677
rect 27437 40605 27483 40643
rect 27437 40571 27443 40605
rect 27477 40571 27483 40605
rect 27437 40533 27483 40571
rect 27437 40499 27443 40533
rect 27477 40499 27483 40533
rect 27437 40461 27483 40499
rect 27437 40427 27443 40461
rect 27477 40427 27483 40461
rect 27437 40389 27483 40427
rect 27437 40355 27443 40389
rect 27477 40355 27483 40389
rect 27437 40317 27483 40355
rect 27437 40283 27443 40317
rect 27477 40283 27483 40317
rect 27437 40245 27483 40283
rect 27437 40211 27443 40245
rect 27477 40211 27483 40245
rect 27437 40173 27483 40211
rect 27437 40139 27443 40173
rect 27477 40139 27483 40173
rect 27437 40101 27483 40139
rect 27437 40067 27443 40101
rect 27477 40067 27483 40101
rect 27437 40029 27483 40067
rect 27437 39995 27443 40029
rect 27477 39995 27483 40029
rect 27437 39957 27483 39995
rect 27437 39923 27443 39957
rect 27477 39923 27483 39957
rect 27437 39907 27483 39923
rect 27895 41181 27941 41197
rect 27895 41147 27901 41181
rect 27935 41147 27941 41181
rect 27895 41109 27941 41147
rect 27895 41075 27901 41109
rect 27935 41075 27941 41109
rect 27895 41037 27941 41075
rect 27895 41003 27901 41037
rect 27935 41003 27941 41037
rect 27895 40965 27941 41003
rect 27895 40931 27901 40965
rect 27935 40931 27941 40965
rect 27895 40893 27941 40931
rect 27895 40859 27901 40893
rect 27935 40859 27941 40893
rect 27895 40821 27941 40859
rect 27895 40787 27901 40821
rect 27935 40787 27941 40821
rect 27895 40749 27941 40787
rect 27895 40715 27901 40749
rect 27935 40715 27941 40749
rect 27895 40677 27941 40715
rect 27895 40643 27901 40677
rect 27935 40643 27941 40677
rect 27895 40605 27941 40643
rect 27895 40571 27901 40605
rect 27935 40571 27941 40605
rect 27895 40533 27941 40571
rect 27895 40499 27901 40533
rect 27935 40499 27941 40533
rect 27895 40461 27941 40499
rect 27895 40427 27901 40461
rect 27935 40427 27941 40461
rect 27895 40389 27941 40427
rect 27895 40355 27901 40389
rect 27935 40355 27941 40389
rect 27895 40317 27941 40355
rect 27895 40283 27901 40317
rect 27935 40283 27941 40317
rect 27895 40245 27941 40283
rect 27895 40211 27901 40245
rect 27935 40211 27941 40245
rect 27895 40173 27941 40211
rect 27895 40139 27901 40173
rect 27935 40139 27941 40173
rect 27895 40101 27941 40139
rect 27895 40067 27901 40101
rect 27935 40067 27941 40101
rect 27895 40029 27941 40067
rect 27895 39995 27901 40029
rect 27935 39995 27941 40029
rect 27895 39957 27941 39995
rect 27895 39923 27901 39957
rect 27935 39923 27941 39957
rect 27895 39907 27941 39923
rect 28353 41181 28399 41197
rect 28353 41147 28359 41181
rect 28393 41147 28399 41181
rect 28353 41109 28399 41147
rect 28353 41075 28359 41109
rect 28393 41075 28399 41109
rect 28353 41037 28399 41075
rect 28353 41003 28359 41037
rect 28393 41003 28399 41037
rect 28353 40965 28399 41003
rect 28353 40931 28359 40965
rect 28393 40931 28399 40965
rect 28353 40893 28399 40931
rect 28353 40859 28359 40893
rect 28393 40859 28399 40893
rect 28353 40821 28399 40859
rect 28353 40787 28359 40821
rect 28393 40787 28399 40821
rect 28353 40749 28399 40787
rect 28353 40715 28359 40749
rect 28393 40715 28399 40749
rect 28353 40677 28399 40715
rect 28353 40643 28359 40677
rect 28393 40643 28399 40677
rect 28353 40605 28399 40643
rect 28353 40571 28359 40605
rect 28393 40571 28399 40605
rect 28353 40533 28399 40571
rect 28353 40499 28359 40533
rect 28393 40499 28399 40533
rect 28353 40461 28399 40499
rect 28353 40427 28359 40461
rect 28393 40427 28399 40461
rect 28353 40389 28399 40427
rect 28353 40355 28359 40389
rect 28393 40355 28399 40389
rect 28353 40317 28399 40355
rect 28353 40283 28359 40317
rect 28393 40283 28399 40317
rect 28353 40245 28399 40283
rect 28353 40211 28359 40245
rect 28393 40211 28399 40245
rect 28353 40173 28399 40211
rect 28353 40139 28359 40173
rect 28393 40139 28399 40173
rect 28353 40101 28399 40139
rect 28353 40067 28359 40101
rect 28393 40067 28399 40101
rect 28353 40029 28399 40067
rect 28353 39995 28359 40029
rect 28393 39995 28399 40029
rect 28353 39957 28399 39995
rect 28353 39923 28359 39957
rect 28393 39923 28399 39957
rect 28353 39907 28399 39923
rect 28811 41181 28857 41197
rect 28811 41147 28817 41181
rect 28851 41147 28857 41181
rect 28811 41109 28857 41147
rect 28811 41075 28817 41109
rect 28851 41075 28857 41109
rect 28811 41037 28857 41075
rect 28811 41003 28817 41037
rect 28851 41003 28857 41037
rect 28811 40965 28857 41003
rect 28811 40931 28817 40965
rect 28851 40931 28857 40965
rect 28811 40893 28857 40931
rect 28811 40859 28817 40893
rect 28851 40859 28857 40893
rect 28811 40821 28857 40859
rect 28811 40787 28817 40821
rect 28851 40787 28857 40821
rect 28811 40749 28857 40787
rect 28811 40715 28817 40749
rect 28851 40715 28857 40749
rect 28811 40677 28857 40715
rect 28811 40643 28817 40677
rect 28851 40643 28857 40677
rect 28811 40605 28857 40643
rect 28811 40571 28817 40605
rect 28851 40571 28857 40605
rect 28811 40533 28857 40571
rect 28811 40499 28817 40533
rect 28851 40499 28857 40533
rect 28811 40461 28857 40499
rect 28811 40427 28817 40461
rect 28851 40427 28857 40461
rect 28811 40389 28857 40427
rect 28811 40355 28817 40389
rect 28851 40355 28857 40389
rect 28811 40317 28857 40355
rect 28811 40283 28817 40317
rect 28851 40283 28857 40317
rect 28811 40245 28857 40283
rect 28811 40211 28817 40245
rect 28851 40211 28857 40245
rect 28811 40173 28857 40211
rect 28811 40139 28817 40173
rect 28851 40139 28857 40173
rect 28811 40101 28857 40139
rect 28811 40067 28817 40101
rect 28851 40067 28857 40101
rect 28811 40029 28857 40067
rect 28811 39995 28817 40029
rect 28851 39995 28857 40029
rect 28811 39957 28857 39995
rect 28811 39923 28817 39957
rect 28851 39923 28857 39957
rect 28811 39907 28857 39923
rect 29269 41181 29315 41197
rect 29269 41147 29275 41181
rect 29309 41147 29315 41181
rect 29269 41109 29315 41147
rect 29269 41075 29275 41109
rect 29309 41075 29315 41109
rect 29269 41037 29315 41075
rect 29269 41003 29275 41037
rect 29309 41003 29315 41037
rect 29269 40965 29315 41003
rect 29269 40931 29275 40965
rect 29309 40931 29315 40965
rect 29269 40893 29315 40931
rect 29269 40859 29275 40893
rect 29309 40859 29315 40893
rect 29269 40821 29315 40859
rect 29269 40787 29275 40821
rect 29309 40787 29315 40821
rect 29269 40749 29315 40787
rect 29269 40715 29275 40749
rect 29309 40715 29315 40749
rect 29269 40677 29315 40715
rect 29269 40643 29275 40677
rect 29309 40643 29315 40677
rect 29269 40605 29315 40643
rect 29269 40571 29275 40605
rect 29309 40571 29315 40605
rect 29269 40533 29315 40571
rect 29269 40499 29275 40533
rect 29309 40499 29315 40533
rect 29269 40461 29315 40499
rect 29269 40427 29275 40461
rect 29309 40427 29315 40461
rect 29269 40389 29315 40427
rect 29269 40355 29275 40389
rect 29309 40355 29315 40389
rect 29269 40317 29315 40355
rect 29269 40283 29275 40317
rect 29309 40283 29315 40317
rect 29269 40245 29315 40283
rect 29269 40211 29275 40245
rect 29309 40211 29315 40245
rect 29269 40173 29315 40211
rect 29269 40139 29275 40173
rect 29309 40139 29315 40173
rect 29269 40101 29315 40139
rect 29269 40067 29275 40101
rect 29309 40067 29315 40101
rect 29269 40029 29315 40067
rect 29269 39995 29275 40029
rect 29309 39995 29315 40029
rect 29269 39957 29315 39995
rect 29269 39923 29275 39957
rect 29309 39923 29315 39957
rect 29269 39907 29315 39923
rect 29727 41181 29773 41197
rect 29727 41147 29733 41181
rect 29767 41147 29773 41181
rect 29727 41109 29773 41147
rect 29727 41075 29733 41109
rect 29767 41075 29773 41109
rect 29727 41037 29773 41075
rect 29727 41003 29733 41037
rect 29767 41003 29773 41037
rect 29727 40965 29773 41003
rect 29727 40931 29733 40965
rect 29767 40931 29773 40965
rect 29727 40893 29773 40931
rect 29727 40859 29733 40893
rect 29767 40859 29773 40893
rect 29727 40821 29773 40859
rect 29727 40787 29733 40821
rect 29767 40787 29773 40821
rect 29727 40749 29773 40787
rect 29727 40715 29733 40749
rect 29767 40715 29773 40749
rect 29727 40677 29773 40715
rect 29727 40643 29733 40677
rect 29767 40643 29773 40677
rect 29727 40605 29773 40643
rect 29727 40571 29733 40605
rect 29767 40571 29773 40605
rect 29727 40533 29773 40571
rect 29727 40499 29733 40533
rect 29767 40499 29773 40533
rect 29727 40461 29773 40499
rect 29727 40427 29733 40461
rect 29767 40427 29773 40461
rect 29727 40389 29773 40427
rect 29727 40355 29733 40389
rect 29767 40355 29773 40389
rect 29727 40317 29773 40355
rect 29727 40283 29733 40317
rect 29767 40283 29773 40317
rect 29727 40245 29773 40283
rect 29727 40211 29733 40245
rect 29767 40211 29773 40245
rect 29727 40173 29773 40211
rect 29727 40139 29733 40173
rect 29767 40139 29773 40173
rect 29727 40101 29773 40139
rect 29727 40067 29733 40101
rect 29767 40067 29773 40101
rect 29727 40029 29773 40067
rect 29727 39995 29733 40029
rect 29767 39995 29773 40029
rect 29727 39957 29773 39995
rect 29727 39923 29733 39957
rect 29767 39923 29773 39957
rect 29727 39907 29773 39923
rect 30185 41181 30231 41197
rect 30185 41147 30191 41181
rect 30225 41147 30231 41181
rect 30185 41109 30231 41147
rect 30185 41075 30191 41109
rect 30225 41075 30231 41109
rect 30185 41037 30231 41075
rect 30185 41003 30191 41037
rect 30225 41003 30231 41037
rect 30185 40965 30231 41003
rect 30185 40931 30191 40965
rect 30225 40931 30231 40965
rect 30185 40893 30231 40931
rect 30185 40859 30191 40893
rect 30225 40859 30231 40893
rect 30185 40821 30231 40859
rect 30185 40787 30191 40821
rect 30225 40787 30231 40821
rect 30185 40749 30231 40787
rect 30185 40715 30191 40749
rect 30225 40715 30231 40749
rect 30185 40677 30231 40715
rect 30185 40643 30191 40677
rect 30225 40643 30231 40677
rect 30185 40605 30231 40643
rect 30185 40571 30191 40605
rect 30225 40571 30231 40605
rect 30185 40533 30231 40571
rect 30185 40499 30191 40533
rect 30225 40499 30231 40533
rect 30185 40461 30231 40499
rect 30185 40427 30191 40461
rect 30225 40427 30231 40461
rect 30185 40389 30231 40427
rect 30185 40355 30191 40389
rect 30225 40355 30231 40389
rect 30185 40317 30231 40355
rect 30185 40283 30191 40317
rect 30225 40283 30231 40317
rect 30185 40245 30231 40283
rect 30185 40211 30191 40245
rect 30225 40211 30231 40245
rect 30185 40173 30231 40211
rect 30185 40139 30191 40173
rect 30225 40139 30231 40173
rect 30185 40101 30231 40139
rect 30185 40067 30191 40101
rect 30225 40067 30231 40101
rect 30185 40029 30231 40067
rect 30185 39995 30191 40029
rect 30225 39995 30231 40029
rect 30185 39957 30231 39995
rect 30185 39923 30191 39957
rect 30225 39923 30231 39957
rect 30185 39907 30231 39923
rect 30643 41181 30689 41197
rect 30643 41147 30649 41181
rect 30683 41147 30689 41181
rect 30643 41109 30689 41147
rect 30643 41075 30649 41109
rect 30683 41075 30689 41109
rect 30643 41037 30689 41075
rect 30643 41003 30649 41037
rect 30683 41003 30689 41037
rect 30643 40965 30689 41003
rect 30643 40931 30649 40965
rect 30683 40931 30689 40965
rect 30643 40893 30689 40931
rect 30643 40859 30649 40893
rect 30683 40859 30689 40893
rect 30643 40821 30689 40859
rect 30643 40787 30649 40821
rect 30683 40787 30689 40821
rect 30643 40749 30689 40787
rect 30643 40715 30649 40749
rect 30683 40715 30689 40749
rect 30643 40677 30689 40715
rect 30643 40643 30649 40677
rect 30683 40643 30689 40677
rect 30643 40605 30689 40643
rect 30643 40571 30649 40605
rect 30683 40571 30689 40605
rect 30643 40533 30689 40571
rect 30643 40499 30649 40533
rect 30683 40499 30689 40533
rect 30643 40461 30689 40499
rect 30643 40427 30649 40461
rect 30683 40427 30689 40461
rect 30643 40389 30689 40427
rect 30643 40355 30649 40389
rect 30683 40355 30689 40389
rect 30643 40317 30689 40355
rect 30643 40283 30649 40317
rect 30683 40283 30689 40317
rect 30643 40245 30689 40283
rect 30643 40211 30649 40245
rect 30683 40211 30689 40245
rect 30643 40173 30689 40211
rect 30643 40139 30649 40173
rect 30683 40139 30689 40173
rect 30643 40101 30689 40139
rect 30643 40067 30649 40101
rect 30683 40067 30689 40101
rect 30643 40029 30689 40067
rect 30643 39995 30649 40029
rect 30683 39995 30689 40029
rect 30643 39957 30689 39995
rect 30643 39923 30649 39957
rect 30683 39923 30689 39957
rect 30643 39907 30689 39923
rect 31101 41181 31147 41197
rect 31101 41147 31107 41181
rect 31141 41147 31147 41181
rect 31101 41109 31147 41147
rect 31101 41075 31107 41109
rect 31141 41075 31147 41109
rect 31101 41037 31147 41075
rect 31101 41003 31107 41037
rect 31141 41003 31147 41037
rect 31101 40965 31147 41003
rect 31101 40931 31107 40965
rect 31141 40931 31147 40965
rect 31101 40893 31147 40931
rect 31101 40859 31107 40893
rect 31141 40859 31147 40893
rect 31101 40821 31147 40859
rect 31101 40787 31107 40821
rect 31141 40787 31147 40821
rect 31101 40749 31147 40787
rect 31101 40715 31107 40749
rect 31141 40715 31147 40749
rect 31101 40677 31147 40715
rect 31101 40643 31107 40677
rect 31141 40643 31147 40677
rect 31101 40605 31147 40643
rect 31101 40571 31107 40605
rect 31141 40571 31147 40605
rect 31101 40533 31147 40571
rect 31101 40499 31107 40533
rect 31141 40499 31147 40533
rect 31101 40461 31147 40499
rect 31101 40427 31107 40461
rect 31141 40427 31147 40461
rect 31101 40389 31147 40427
rect 31101 40355 31107 40389
rect 31141 40355 31147 40389
rect 31101 40317 31147 40355
rect 31101 40283 31107 40317
rect 31141 40283 31147 40317
rect 31101 40245 31147 40283
rect 31101 40211 31107 40245
rect 31141 40211 31147 40245
rect 31101 40173 31147 40211
rect 31101 40139 31107 40173
rect 31141 40139 31147 40173
rect 31101 40101 31147 40139
rect 31101 40067 31107 40101
rect 31141 40067 31147 40101
rect 31101 40029 31147 40067
rect 31101 39995 31107 40029
rect 31141 39995 31147 40029
rect 31101 39957 31147 39995
rect 31101 39923 31107 39957
rect 31141 39923 31147 39957
rect 31101 39907 31147 39923
rect 31559 41181 31605 41197
rect 31559 41147 31565 41181
rect 31599 41147 31605 41181
rect 31559 41109 31605 41147
rect 31559 41075 31565 41109
rect 31599 41075 31605 41109
rect 31559 41037 31605 41075
rect 31559 41003 31565 41037
rect 31599 41003 31605 41037
rect 31559 40965 31605 41003
rect 31559 40931 31565 40965
rect 31599 40931 31605 40965
rect 31559 40893 31605 40931
rect 31559 40859 31565 40893
rect 31599 40859 31605 40893
rect 31559 40821 31605 40859
rect 31559 40787 31565 40821
rect 31599 40787 31605 40821
rect 31559 40749 31605 40787
rect 31559 40715 31565 40749
rect 31599 40715 31605 40749
rect 31559 40677 31605 40715
rect 31559 40643 31565 40677
rect 31599 40643 31605 40677
rect 31559 40605 31605 40643
rect 31559 40571 31565 40605
rect 31599 40571 31605 40605
rect 31559 40533 31605 40571
rect 31559 40499 31565 40533
rect 31599 40499 31605 40533
rect 31559 40461 31605 40499
rect 31559 40427 31565 40461
rect 31599 40427 31605 40461
rect 31559 40389 31605 40427
rect 31559 40355 31565 40389
rect 31599 40355 31605 40389
rect 31559 40317 31605 40355
rect 31559 40283 31565 40317
rect 31599 40283 31605 40317
rect 31559 40245 31605 40283
rect 31559 40211 31565 40245
rect 31599 40211 31605 40245
rect 31559 40173 31605 40211
rect 31559 40139 31565 40173
rect 31599 40139 31605 40173
rect 31559 40101 31605 40139
rect 31559 40067 31565 40101
rect 31599 40067 31605 40101
rect 31559 40029 31605 40067
rect 31559 39995 31565 40029
rect 31599 39995 31605 40029
rect 31559 39957 31605 39995
rect 31559 39923 31565 39957
rect 31599 39923 31605 39957
rect 31559 39907 31605 39923
rect 32017 41181 32063 41197
rect 32017 41147 32023 41181
rect 32057 41147 32063 41181
rect 32017 41109 32063 41147
rect 32017 41075 32023 41109
rect 32057 41075 32063 41109
rect 32017 41037 32063 41075
rect 32017 41003 32023 41037
rect 32057 41003 32063 41037
rect 32017 40965 32063 41003
rect 32017 40931 32023 40965
rect 32057 40931 32063 40965
rect 32017 40893 32063 40931
rect 32017 40859 32023 40893
rect 32057 40859 32063 40893
rect 32017 40821 32063 40859
rect 32017 40787 32023 40821
rect 32057 40787 32063 40821
rect 32017 40749 32063 40787
rect 32017 40715 32023 40749
rect 32057 40715 32063 40749
rect 32017 40677 32063 40715
rect 32017 40643 32023 40677
rect 32057 40643 32063 40677
rect 32017 40605 32063 40643
rect 32017 40571 32023 40605
rect 32057 40571 32063 40605
rect 32017 40533 32063 40571
rect 32017 40499 32023 40533
rect 32057 40499 32063 40533
rect 32017 40461 32063 40499
rect 32017 40427 32023 40461
rect 32057 40427 32063 40461
rect 32017 40389 32063 40427
rect 32017 40355 32023 40389
rect 32057 40355 32063 40389
rect 32017 40317 32063 40355
rect 32017 40283 32023 40317
rect 32057 40283 32063 40317
rect 32017 40245 32063 40283
rect 32017 40211 32023 40245
rect 32057 40211 32063 40245
rect 32017 40173 32063 40211
rect 32017 40139 32023 40173
rect 32057 40139 32063 40173
rect 32017 40101 32063 40139
rect 32017 40067 32023 40101
rect 32057 40067 32063 40101
rect 32017 40029 32063 40067
rect 32017 39995 32023 40029
rect 32057 39995 32063 40029
rect 32017 39957 32063 39995
rect 32017 39923 32023 39957
rect 32057 39923 32063 39957
rect 32017 39907 32063 39923
rect 32475 41181 32521 41197
rect 32475 41147 32481 41181
rect 32515 41147 32521 41181
rect 32475 41109 32521 41147
rect 32475 41075 32481 41109
rect 32515 41075 32521 41109
rect 32475 41037 32521 41075
rect 32475 41003 32481 41037
rect 32515 41003 32521 41037
rect 32475 40965 32521 41003
rect 32475 40931 32481 40965
rect 32515 40931 32521 40965
rect 32475 40893 32521 40931
rect 32475 40859 32481 40893
rect 32515 40859 32521 40893
rect 32475 40821 32521 40859
rect 32475 40787 32481 40821
rect 32515 40787 32521 40821
rect 32475 40749 32521 40787
rect 32475 40715 32481 40749
rect 32515 40715 32521 40749
rect 32475 40677 32521 40715
rect 32475 40643 32481 40677
rect 32515 40643 32521 40677
rect 32475 40605 32521 40643
rect 32475 40571 32481 40605
rect 32515 40571 32521 40605
rect 32475 40533 32521 40571
rect 32475 40499 32481 40533
rect 32515 40499 32521 40533
rect 32475 40461 32521 40499
rect 32475 40427 32481 40461
rect 32515 40427 32521 40461
rect 32475 40389 32521 40427
rect 32475 40355 32481 40389
rect 32515 40355 32521 40389
rect 32475 40317 32521 40355
rect 32475 40283 32481 40317
rect 32515 40283 32521 40317
rect 32475 40245 32521 40283
rect 32475 40211 32481 40245
rect 32515 40211 32521 40245
rect 32475 40173 32521 40211
rect 32475 40139 32481 40173
rect 32515 40139 32521 40173
rect 32475 40101 32521 40139
rect 32475 40067 32481 40101
rect 32515 40067 32521 40101
rect 32475 40029 32521 40067
rect 32475 39995 32481 40029
rect 32515 39995 32521 40029
rect 32475 39957 32521 39995
rect 32475 39923 32481 39957
rect 32515 39923 32521 39957
rect 32475 39907 32521 39923
rect 32933 41181 32979 41197
rect 32933 41147 32939 41181
rect 32973 41147 32979 41181
rect 32933 41109 32979 41147
rect 32933 41075 32939 41109
rect 32973 41075 32979 41109
rect 32933 41037 32979 41075
rect 32933 41003 32939 41037
rect 32973 41003 32979 41037
rect 32933 40965 32979 41003
rect 32933 40931 32939 40965
rect 32973 40931 32979 40965
rect 32933 40893 32979 40931
rect 32933 40859 32939 40893
rect 32973 40859 32979 40893
rect 32933 40821 32979 40859
rect 32933 40787 32939 40821
rect 32973 40787 32979 40821
rect 32933 40749 32979 40787
rect 32933 40715 32939 40749
rect 32973 40715 32979 40749
rect 32933 40677 32979 40715
rect 32933 40643 32939 40677
rect 32973 40643 32979 40677
rect 32933 40605 32979 40643
rect 32933 40571 32939 40605
rect 32973 40571 32979 40605
rect 32933 40533 32979 40571
rect 32933 40499 32939 40533
rect 32973 40499 32979 40533
rect 32933 40461 32979 40499
rect 32933 40427 32939 40461
rect 32973 40427 32979 40461
rect 32933 40389 32979 40427
rect 32933 40355 32939 40389
rect 32973 40355 32979 40389
rect 32933 40317 32979 40355
rect 32933 40283 32939 40317
rect 32973 40283 32979 40317
rect 32933 40245 32979 40283
rect 32933 40211 32939 40245
rect 32973 40211 32979 40245
rect 32933 40173 32979 40211
rect 32933 40139 32939 40173
rect 32973 40139 32979 40173
rect 32933 40101 32979 40139
rect 32933 40067 32939 40101
rect 32973 40067 32979 40101
rect 32933 40029 32979 40067
rect 32933 39995 32939 40029
rect 32973 39995 32979 40029
rect 32933 39957 32979 39995
rect 32933 39923 32939 39957
rect 32973 39923 32979 39957
rect 32933 39907 32979 39923
rect 33391 41181 33437 41197
rect 33391 41147 33397 41181
rect 33431 41147 33437 41181
rect 33391 41109 33437 41147
rect 33391 41075 33397 41109
rect 33431 41075 33437 41109
rect 33391 41037 33437 41075
rect 33391 41003 33397 41037
rect 33431 41003 33437 41037
rect 33391 40965 33437 41003
rect 33391 40931 33397 40965
rect 33431 40931 33437 40965
rect 33391 40893 33437 40931
rect 33391 40859 33397 40893
rect 33431 40859 33437 40893
rect 33391 40821 33437 40859
rect 33391 40787 33397 40821
rect 33431 40787 33437 40821
rect 33391 40749 33437 40787
rect 33391 40715 33397 40749
rect 33431 40715 33437 40749
rect 33391 40677 33437 40715
rect 33391 40643 33397 40677
rect 33431 40643 33437 40677
rect 33391 40605 33437 40643
rect 33391 40571 33397 40605
rect 33431 40571 33437 40605
rect 33391 40533 33437 40571
rect 33391 40499 33397 40533
rect 33431 40499 33437 40533
rect 33391 40461 33437 40499
rect 33391 40427 33397 40461
rect 33431 40427 33437 40461
rect 33391 40389 33437 40427
rect 33391 40355 33397 40389
rect 33431 40355 33437 40389
rect 33391 40317 33437 40355
rect 33391 40283 33397 40317
rect 33431 40283 33437 40317
rect 33391 40245 33437 40283
rect 33391 40211 33397 40245
rect 33431 40211 33437 40245
rect 33391 40173 33437 40211
rect 33391 40139 33397 40173
rect 33431 40139 33437 40173
rect 33391 40101 33437 40139
rect 33391 40067 33397 40101
rect 33431 40067 33437 40101
rect 33391 40029 33437 40067
rect 33391 39995 33397 40029
rect 33431 39995 33437 40029
rect 33391 39957 33437 39995
rect 33391 39923 33397 39957
rect 33431 39923 33437 39957
rect 33391 39907 33437 39923
rect 33849 41181 33895 41197
rect 33849 41147 33855 41181
rect 33889 41147 33895 41181
rect 33849 41109 33895 41147
rect 33849 41075 33855 41109
rect 33889 41075 33895 41109
rect 33849 41037 33895 41075
rect 33849 41003 33855 41037
rect 33889 41003 33895 41037
rect 33849 40965 33895 41003
rect 33849 40931 33855 40965
rect 33889 40931 33895 40965
rect 33849 40893 33895 40931
rect 33849 40859 33855 40893
rect 33889 40859 33895 40893
rect 33849 40821 33895 40859
rect 33849 40787 33855 40821
rect 33889 40787 33895 40821
rect 33849 40749 33895 40787
rect 33849 40715 33855 40749
rect 33889 40715 33895 40749
rect 33849 40677 33895 40715
rect 33849 40643 33855 40677
rect 33889 40643 33895 40677
rect 33849 40605 33895 40643
rect 33849 40571 33855 40605
rect 33889 40571 33895 40605
rect 33849 40533 33895 40571
rect 33849 40499 33855 40533
rect 33889 40499 33895 40533
rect 33849 40461 33895 40499
rect 33849 40427 33855 40461
rect 33889 40427 33895 40461
rect 33849 40389 33895 40427
rect 33849 40355 33855 40389
rect 33889 40355 33895 40389
rect 33849 40317 33895 40355
rect 33849 40283 33855 40317
rect 33889 40283 33895 40317
rect 33849 40245 33895 40283
rect 33849 40211 33855 40245
rect 33889 40211 33895 40245
rect 33849 40173 33895 40211
rect 33849 40139 33855 40173
rect 33889 40139 33895 40173
rect 33849 40101 33895 40139
rect 33849 40067 33855 40101
rect 33889 40067 33895 40101
rect 33849 40029 33895 40067
rect 33849 39995 33855 40029
rect 33889 39995 33895 40029
rect 33849 39957 33895 39995
rect 33849 39923 33855 39957
rect 33889 39923 33895 39957
rect 33849 39907 33895 39923
rect 34307 41181 34353 41197
rect 34307 41147 34313 41181
rect 34347 41147 34353 41181
rect 34307 41109 34353 41147
rect 34307 41075 34313 41109
rect 34347 41075 34353 41109
rect 34307 41037 34353 41075
rect 34307 41003 34313 41037
rect 34347 41003 34353 41037
rect 34307 40965 34353 41003
rect 34307 40931 34313 40965
rect 34347 40931 34353 40965
rect 34307 40893 34353 40931
rect 34307 40859 34313 40893
rect 34347 40859 34353 40893
rect 34307 40821 34353 40859
rect 34307 40787 34313 40821
rect 34347 40787 34353 40821
rect 34307 40749 34353 40787
rect 34307 40715 34313 40749
rect 34347 40715 34353 40749
rect 34307 40677 34353 40715
rect 34307 40643 34313 40677
rect 34347 40643 34353 40677
rect 34307 40605 34353 40643
rect 34307 40571 34313 40605
rect 34347 40571 34353 40605
rect 34307 40533 34353 40571
rect 34307 40499 34313 40533
rect 34347 40499 34353 40533
rect 34307 40461 34353 40499
rect 34307 40427 34313 40461
rect 34347 40427 34353 40461
rect 34307 40389 34353 40427
rect 34307 40355 34313 40389
rect 34347 40355 34353 40389
rect 34307 40317 34353 40355
rect 34307 40283 34313 40317
rect 34347 40283 34353 40317
rect 34307 40245 34353 40283
rect 34307 40211 34313 40245
rect 34347 40211 34353 40245
rect 34307 40173 34353 40211
rect 34307 40139 34313 40173
rect 34347 40139 34353 40173
rect 34307 40101 34353 40139
rect 34307 40067 34313 40101
rect 34347 40067 34353 40101
rect 34307 40029 34353 40067
rect 34307 39995 34313 40029
rect 34347 39995 34353 40029
rect 34307 39957 34353 39995
rect 34307 39923 34313 39957
rect 34347 39923 34353 39957
rect 34307 39907 34353 39923
rect 34765 41181 34811 41197
rect 34765 41147 34771 41181
rect 34805 41147 34811 41181
rect 34765 41109 34811 41147
rect 34765 41075 34771 41109
rect 34805 41075 34811 41109
rect 34765 41037 34811 41075
rect 34765 41003 34771 41037
rect 34805 41003 34811 41037
rect 34765 40965 34811 41003
rect 34765 40931 34771 40965
rect 34805 40931 34811 40965
rect 34765 40893 34811 40931
rect 34765 40859 34771 40893
rect 34805 40859 34811 40893
rect 34765 40821 34811 40859
rect 34765 40787 34771 40821
rect 34805 40787 34811 40821
rect 34765 40749 34811 40787
rect 34765 40715 34771 40749
rect 34805 40715 34811 40749
rect 34765 40677 34811 40715
rect 34765 40643 34771 40677
rect 34805 40643 34811 40677
rect 34765 40605 34811 40643
rect 34765 40571 34771 40605
rect 34805 40571 34811 40605
rect 34765 40533 34811 40571
rect 34765 40499 34771 40533
rect 34805 40499 34811 40533
rect 34765 40461 34811 40499
rect 34765 40427 34771 40461
rect 34805 40427 34811 40461
rect 34765 40389 34811 40427
rect 34765 40355 34771 40389
rect 34805 40355 34811 40389
rect 34765 40317 34811 40355
rect 34765 40283 34771 40317
rect 34805 40283 34811 40317
rect 34765 40245 34811 40283
rect 34765 40211 34771 40245
rect 34805 40211 34811 40245
rect 34765 40173 34811 40211
rect 34765 40139 34771 40173
rect 34805 40139 34811 40173
rect 34765 40101 34811 40139
rect 34765 40067 34771 40101
rect 34805 40067 34811 40101
rect 34765 40029 34811 40067
rect 34765 39995 34771 40029
rect 34805 39995 34811 40029
rect 34765 39957 34811 39995
rect 34765 39923 34771 39957
rect 34805 39923 34811 39957
rect 34765 39907 34811 39923
rect 35223 41181 35269 41197
rect 35223 41147 35229 41181
rect 35263 41147 35269 41181
rect 35223 41109 35269 41147
rect 35223 41075 35229 41109
rect 35263 41075 35269 41109
rect 35223 41037 35269 41075
rect 35223 41003 35229 41037
rect 35263 41003 35269 41037
rect 35223 40965 35269 41003
rect 35223 40931 35229 40965
rect 35263 40931 35269 40965
rect 35223 40893 35269 40931
rect 35223 40859 35229 40893
rect 35263 40859 35269 40893
rect 35223 40821 35269 40859
rect 35223 40787 35229 40821
rect 35263 40787 35269 40821
rect 35223 40749 35269 40787
rect 35223 40715 35229 40749
rect 35263 40715 35269 40749
rect 35223 40677 35269 40715
rect 35223 40643 35229 40677
rect 35263 40643 35269 40677
rect 35223 40605 35269 40643
rect 35223 40571 35229 40605
rect 35263 40571 35269 40605
rect 35223 40533 35269 40571
rect 35223 40499 35229 40533
rect 35263 40499 35269 40533
rect 35223 40461 35269 40499
rect 35223 40427 35229 40461
rect 35263 40427 35269 40461
rect 35223 40389 35269 40427
rect 35223 40355 35229 40389
rect 35263 40355 35269 40389
rect 35223 40317 35269 40355
rect 35223 40283 35229 40317
rect 35263 40283 35269 40317
rect 35223 40245 35269 40283
rect 35223 40211 35229 40245
rect 35263 40211 35269 40245
rect 35223 40173 35269 40211
rect 35223 40139 35229 40173
rect 35263 40139 35269 40173
rect 35223 40101 35269 40139
rect 35223 40067 35229 40101
rect 35263 40067 35269 40101
rect 35223 40029 35269 40067
rect 35223 39995 35229 40029
rect 35263 39995 35269 40029
rect 35223 39957 35269 39995
rect 35223 39923 35229 39957
rect 35263 39923 35269 39957
rect 35223 39907 35269 39923
rect 35681 41181 35727 41197
rect 35681 41147 35687 41181
rect 35721 41147 35727 41181
rect 35681 41109 35727 41147
rect 35681 41075 35687 41109
rect 35721 41075 35727 41109
rect 35681 41037 35727 41075
rect 35681 41003 35687 41037
rect 35721 41003 35727 41037
rect 35681 40965 35727 41003
rect 35681 40931 35687 40965
rect 35721 40931 35727 40965
rect 35681 40893 35727 40931
rect 35681 40859 35687 40893
rect 35721 40859 35727 40893
rect 35681 40821 35727 40859
rect 35681 40787 35687 40821
rect 35721 40787 35727 40821
rect 35681 40749 35727 40787
rect 35681 40715 35687 40749
rect 35721 40715 35727 40749
rect 35681 40677 35727 40715
rect 35681 40643 35687 40677
rect 35721 40643 35727 40677
rect 35681 40605 35727 40643
rect 35681 40571 35687 40605
rect 35721 40571 35727 40605
rect 35681 40533 35727 40571
rect 35681 40499 35687 40533
rect 35721 40499 35727 40533
rect 35681 40461 35727 40499
rect 35681 40427 35687 40461
rect 35721 40427 35727 40461
rect 35681 40389 35727 40427
rect 35681 40355 35687 40389
rect 35721 40355 35727 40389
rect 35681 40317 35727 40355
rect 35681 40283 35687 40317
rect 35721 40283 35727 40317
rect 35681 40245 35727 40283
rect 35681 40211 35687 40245
rect 35721 40211 35727 40245
rect 35681 40173 35727 40211
rect 35681 40139 35687 40173
rect 35721 40139 35727 40173
rect 35681 40101 35727 40139
rect 35681 40067 35687 40101
rect 35721 40067 35727 40101
rect 35681 40029 35727 40067
rect 35681 39995 35687 40029
rect 35721 39995 35727 40029
rect 35681 39957 35727 39995
rect 35681 39923 35687 39957
rect 35721 39923 35727 39957
rect 35681 39907 35727 39923
rect 36139 41181 36185 41197
rect 36139 41147 36145 41181
rect 36179 41147 36185 41181
rect 36139 41109 36185 41147
rect 36139 41075 36145 41109
rect 36179 41075 36185 41109
rect 36139 41037 36185 41075
rect 36139 41003 36145 41037
rect 36179 41003 36185 41037
rect 36139 40965 36185 41003
rect 36139 40931 36145 40965
rect 36179 40931 36185 40965
rect 36139 40893 36185 40931
rect 36139 40859 36145 40893
rect 36179 40859 36185 40893
rect 36139 40821 36185 40859
rect 36139 40787 36145 40821
rect 36179 40787 36185 40821
rect 36139 40749 36185 40787
rect 36139 40715 36145 40749
rect 36179 40715 36185 40749
rect 36139 40677 36185 40715
rect 36139 40643 36145 40677
rect 36179 40643 36185 40677
rect 36139 40605 36185 40643
rect 36139 40571 36145 40605
rect 36179 40571 36185 40605
rect 36139 40533 36185 40571
rect 36139 40499 36145 40533
rect 36179 40499 36185 40533
rect 36139 40461 36185 40499
rect 36139 40427 36145 40461
rect 36179 40427 36185 40461
rect 36139 40389 36185 40427
rect 36139 40355 36145 40389
rect 36179 40355 36185 40389
rect 36139 40317 36185 40355
rect 36139 40283 36145 40317
rect 36179 40283 36185 40317
rect 36139 40245 36185 40283
rect 36139 40211 36145 40245
rect 36179 40211 36185 40245
rect 36139 40173 36185 40211
rect 36139 40139 36145 40173
rect 36179 40139 36185 40173
rect 36139 40101 36185 40139
rect 36139 40067 36145 40101
rect 36179 40067 36185 40101
rect 36139 40029 36185 40067
rect 36139 39995 36145 40029
rect 36179 39995 36185 40029
rect 36139 39957 36185 39995
rect 36139 39923 36145 39957
rect 36179 39923 36185 39957
rect 36139 39907 36185 39923
rect 36597 41181 36643 41197
rect 36597 41147 36603 41181
rect 36637 41147 36643 41181
rect 36597 41109 36643 41147
rect 36597 41075 36603 41109
rect 36637 41075 36643 41109
rect 36597 41037 36643 41075
rect 36597 41003 36603 41037
rect 36637 41003 36643 41037
rect 36597 40965 36643 41003
rect 36597 40931 36603 40965
rect 36637 40931 36643 40965
rect 36597 40893 36643 40931
rect 36597 40859 36603 40893
rect 36637 40859 36643 40893
rect 36597 40821 36643 40859
rect 36597 40787 36603 40821
rect 36637 40787 36643 40821
rect 36597 40749 36643 40787
rect 36597 40715 36603 40749
rect 36637 40715 36643 40749
rect 36597 40677 36643 40715
rect 36597 40643 36603 40677
rect 36637 40643 36643 40677
rect 36597 40605 36643 40643
rect 36597 40571 36603 40605
rect 36637 40571 36643 40605
rect 36597 40533 36643 40571
rect 36597 40499 36603 40533
rect 36637 40499 36643 40533
rect 36597 40461 36643 40499
rect 36597 40427 36603 40461
rect 36637 40427 36643 40461
rect 36597 40389 36643 40427
rect 36597 40355 36603 40389
rect 36637 40355 36643 40389
rect 36597 40317 36643 40355
rect 36597 40283 36603 40317
rect 36637 40283 36643 40317
rect 36597 40245 36643 40283
rect 36597 40211 36603 40245
rect 36637 40211 36643 40245
rect 36597 40173 36643 40211
rect 36597 40139 36603 40173
rect 36637 40139 36643 40173
rect 36597 40101 36643 40139
rect 36597 40067 36603 40101
rect 36637 40067 36643 40101
rect 36597 40029 36643 40067
rect 36597 39995 36603 40029
rect 36637 39995 36643 40029
rect 36597 39957 36643 39995
rect 36597 39923 36603 39957
rect 36637 39923 36643 39957
rect 36597 39907 36643 39923
rect 37055 41181 37101 41197
rect 37055 41147 37061 41181
rect 37095 41147 37101 41181
rect 37055 41109 37101 41147
rect 37055 41075 37061 41109
rect 37095 41075 37101 41109
rect 37055 41037 37101 41075
rect 37055 41003 37061 41037
rect 37095 41003 37101 41037
rect 37055 40965 37101 41003
rect 37055 40931 37061 40965
rect 37095 40931 37101 40965
rect 37055 40893 37101 40931
rect 37055 40859 37061 40893
rect 37095 40859 37101 40893
rect 37055 40821 37101 40859
rect 37055 40787 37061 40821
rect 37095 40787 37101 40821
rect 37055 40749 37101 40787
rect 37055 40715 37061 40749
rect 37095 40715 37101 40749
rect 37055 40677 37101 40715
rect 37055 40643 37061 40677
rect 37095 40643 37101 40677
rect 37055 40605 37101 40643
rect 37055 40571 37061 40605
rect 37095 40571 37101 40605
rect 37055 40533 37101 40571
rect 37055 40499 37061 40533
rect 37095 40499 37101 40533
rect 37055 40461 37101 40499
rect 37055 40427 37061 40461
rect 37095 40427 37101 40461
rect 37055 40389 37101 40427
rect 37055 40355 37061 40389
rect 37095 40355 37101 40389
rect 37055 40317 37101 40355
rect 37055 40283 37061 40317
rect 37095 40283 37101 40317
rect 37055 40245 37101 40283
rect 37055 40211 37061 40245
rect 37095 40211 37101 40245
rect 37055 40173 37101 40211
rect 37055 40139 37061 40173
rect 37095 40139 37101 40173
rect 37055 40101 37101 40139
rect 37055 40067 37061 40101
rect 37095 40067 37101 40101
rect 37055 40029 37101 40067
rect 37055 39995 37061 40029
rect 37095 39995 37101 40029
rect 37055 39957 37101 39995
rect 37055 39923 37061 39957
rect 37095 39923 37101 39957
rect 37055 39907 37101 39923
rect 37513 41181 37559 41197
rect 37513 41147 37519 41181
rect 37553 41147 37559 41181
rect 37513 41109 37559 41147
rect 37513 41075 37519 41109
rect 37553 41075 37559 41109
rect 37513 41037 37559 41075
rect 37513 41003 37519 41037
rect 37553 41003 37559 41037
rect 37513 40965 37559 41003
rect 37513 40931 37519 40965
rect 37553 40931 37559 40965
rect 37513 40893 37559 40931
rect 37513 40859 37519 40893
rect 37553 40859 37559 40893
rect 37513 40821 37559 40859
rect 37513 40787 37519 40821
rect 37553 40787 37559 40821
rect 37513 40749 37559 40787
rect 37513 40715 37519 40749
rect 37553 40715 37559 40749
rect 37513 40677 37559 40715
rect 37513 40643 37519 40677
rect 37553 40643 37559 40677
rect 37513 40605 37559 40643
rect 37513 40571 37519 40605
rect 37553 40571 37559 40605
rect 37513 40533 37559 40571
rect 37513 40499 37519 40533
rect 37553 40499 37559 40533
rect 37513 40461 37559 40499
rect 37513 40427 37519 40461
rect 37553 40427 37559 40461
rect 37513 40389 37559 40427
rect 37513 40355 37519 40389
rect 37553 40355 37559 40389
rect 37513 40317 37559 40355
rect 37513 40283 37519 40317
rect 37553 40283 37559 40317
rect 37513 40245 37559 40283
rect 37513 40211 37519 40245
rect 37553 40211 37559 40245
rect 37513 40173 37559 40211
rect 37513 40139 37519 40173
rect 37553 40139 37559 40173
rect 37513 40101 37559 40139
rect 37513 40067 37519 40101
rect 37553 40067 37559 40101
rect 37513 40029 37559 40067
rect 37513 39995 37519 40029
rect 37553 39995 37559 40029
rect 37513 39957 37559 39995
rect 37513 39923 37519 39957
rect 37553 39923 37559 39957
rect 37513 39907 37559 39923
rect 37971 41181 38017 41197
rect 37971 41147 37977 41181
rect 38011 41147 38017 41181
rect 37971 41109 38017 41147
rect 37971 41075 37977 41109
rect 38011 41075 38017 41109
rect 37971 41037 38017 41075
rect 37971 41003 37977 41037
rect 38011 41003 38017 41037
rect 37971 40965 38017 41003
rect 37971 40931 37977 40965
rect 38011 40931 38017 40965
rect 37971 40893 38017 40931
rect 37971 40859 37977 40893
rect 38011 40859 38017 40893
rect 37971 40821 38017 40859
rect 37971 40787 37977 40821
rect 38011 40787 38017 40821
rect 37971 40749 38017 40787
rect 37971 40715 37977 40749
rect 38011 40715 38017 40749
rect 37971 40677 38017 40715
rect 37971 40643 37977 40677
rect 38011 40643 38017 40677
rect 37971 40605 38017 40643
rect 37971 40571 37977 40605
rect 38011 40571 38017 40605
rect 37971 40533 38017 40571
rect 37971 40499 37977 40533
rect 38011 40499 38017 40533
rect 37971 40461 38017 40499
rect 37971 40427 37977 40461
rect 38011 40427 38017 40461
rect 37971 40389 38017 40427
rect 37971 40355 37977 40389
rect 38011 40355 38017 40389
rect 37971 40317 38017 40355
rect 37971 40283 37977 40317
rect 38011 40283 38017 40317
rect 37971 40245 38017 40283
rect 37971 40211 37977 40245
rect 38011 40211 38017 40245
rect 37971 40173 38017 40211
rect 37971 40139 37977 40173
rect 38011 40139 38017 40173
rect 37971 40101 38017 40139
rect 37971 40067 37977 40101
rect 38011 40067 38017 40101
rect 37971 40029 38017 40067
rect 37971 39995 37977 40029
rect 38011 39995 38017 40029
rect 37971 39957 38017 39995
rect 37971 39923 37977 39957
rect 38011 39923 38017 39957
rect 37971 39907 38017 39923
rect 38429 41181 38475 41197
rect 38429 41147 38435 41181
rect 38469 41147 38475 41181
rect 38429 41109 38475 41147
rect 38429 41075 38435 41109
rect 38469 41075 38475 41109
rect 38429 41037 38475 41075
rect 38429 41003 38435 41037
rect 38469 41003 38475 41037
rect 38429 40965 38475 41003
rect 38429 40931 38435 40965
rect 38469 40931 38475 40965
rect 38429 40893 38475 40931
rect 38429 40859 38435 40893
rect 38469 40859 38475 40893
rect 38429 40821 38475 40859
rect 38429 40787 38435 40821
rect 38469 40787 38475 40821
rect 38429 40749 38475 40787
rect 38429 40715 38435 40749
rect 38469 40715 38475 40749
rect 38429 40677 38475 40715
rect 38429 40643 38435 40677
rect 38469 40643 38475 40677
rect 38429 40605 38475 40643
rect 38429 40571 38435 40605
rect 38469 40571 38475 40605
rect 38429 40533 38475 40571
rect 38429 40499 38435 40533
rect 38469 40499 38475 40533
rect 38429 40461 38475 40499
rect 38429 40427 38435 40461
rect 38469 40427 38475 40461
rect 38429 40389 38475 40427
rect 38429 40355 38435 40389
rect 38469 40355 38475 40389
rect 38429 40317 38475 40355
rect 38429 40283 38435 40317
rect 38469 40283 38475 40317
rect 38429 40245 38475 40283
rect 38429 40211 38435 40245
rect 38469 40211 38475 40245
rect 38429 40173 38475 40211
rect 38429 40139 38435 40173
rect 38469 40139 38475 40173
rect 38429 40101 38475 40139
rect 38429 40067 38435 40101
rect 38469 40067 38475 40101
rect 38429 40029 38475 40067
rect 38429 39995 38435 40029
rect 38469 39995 38475 40029
rect 38429 39957 38475 39995
rect 38429 39923 38435 39957
rect 38469 39923 38475 39957
rect 38429 39907 38475 39923
rect 38887 41181 38933 41197
rect 38887 41147 38893 41181
rect 38927 41147 38933 41181
rect 38887 41109 38933 41147
rect 38887 41075 38893 41109
rect 38927 41075 38933 41109
rect 38887 41037 38933 41075
rect 38887 41003 38893 41037
rect 38927 41003 38933 41037
rect 38887 40965 38933 41003
rect 38887 40931 38893 40965
rect 38927 40931 38933 40965
rect 38887 40893 38933 40931
rect 38887 40859 38893 40893
rect 38927 40859 38933 40893
rect 38887 40821 38933 40859
rect 38887 40787 38893 40821
rect 38927 40787 38933 40821
rect 38887 40749 38933 40787
rect 38887 40715 38893 40749
rect 38927 40715 38933 40749
rect 38887 40677 38933 40715
rect 38887 40643 38893 40677
rect 38927 40643 38933 40677
rect 38887 40605 38933 40643
rect 38887 40571 38893 40605
rect 38927 40571 38933 40605
rect 38887 40533 38933 40571
rect 38887 40499 38893 40533
rect 38927 40499 38933 40533
rect 38887 40461 38933 40499
rect 38887 40427 38893 40461
rect 38927 40427 38933 40461
rect 38887 40389 38933 40427
rect 38887 40355 38893 40389
rect 38927 40355 38933 40389
rect 38887 40317 38933 40355
rect 38887 40283 38893 40317
rect 38927 40283 38933 40317
rect 38887 40245 38933 40283
rect 38887 40211 38893 40245
rect 38927 40211 38933 40245
rect 38887 40173 38933 40211
rect 38887 40139 38893 40173
rect 38927 40139 38933 40173
rect 38887 40101 38933 40139
rect 38887 40067 38893 40101
rect 38927 40067 38933 40101
rect 38887 40029 38933 40067
rect 38887 39995 38893 40029
rect 38927 39995 38933 40029
rect 38887 39957 38933 39995
rect 38887 39923 38893 39957
rect 38927 39923 38933 39957
rect 38887 39907 38933 39923
rect 39345 41181 39391 41197
rect 39345 41147 39351 41181
rect 39385 41147 39391 41181
rect 39345 41109 39391 41147
rect 39345 41075 39351 41109
rect 39385 41075 39391 41109
rect 39345 41037 39391 41075
rect 39345 41003 39351 41037
rect 39385 41003 39391 41037
rect 39345 40965 39391 41003
rect 39345 40931 39351 40965
rect 39385 40931 39391 40965
rect 39345 40893 39391 40931
rect 39345 40859 39351 40893
rect 39385 40859 39391 40893
rect 39345 40821 39391 40859
rect 39345 40787 39351 40821
rect 39385 40787 39391 40821
rect 39345 40749 39391 40787
rect 39345 40715 39351 40749
rect 39385 40715 39391 40749
rect 39345 40677 39391 40715
rect 39345 40643 39351 40677
rect 39385 40643 39391 40677
rect 39345 40605 39391 40643
rect 39345 40571 39351 40605
rect 39385 40571 39391 40605
rect 39345 40533 39391 40571
rect 39345 40499 39351 40533
rect 39385 40499 39391 40533
rect 39345 40461 39391 40499
rect 39345 40427 39351 40461
rect 39385 40427 39391 40461
rect 39345 40389 39391 40427
rect 39345 40355 39351 40389
rect 39385 40355 39391 40389
rect 39345 40317 39391 40355
rect 39345 40283 39351 40317
rect 39385 40283 39391 40317
rect 39345 40245 39391 40283
rect 39345 40211 39351 40245
rect 39385 40211 39391 40245
rect 39345 40173 39391 40211
rect 39345 40139 39351 40173
rect 39385 40139 39391 40173
rect 39345 40101 39391 40139
rect 39345 40067 39351 40101
rect 39385 40067 39391 40101
rect 39345 40029 39391 40067
rect 39345 39995 39351 40029
rect 39385 39995 39391 40029
rect 39345 39957 39391 39995
rect 39345 39923 39351 39957
rect 39385 39923 39391 39957
rect 39345 39907 39391 39923
rect 39803 41181 39849 41197
rect 39803 41147 39809 41181
rect 39843 41147 39849 41181
rect 39803 41109 39849 41147
rect 39803 41075 39809 41109
rect 39843 41075 39849 41109
rect 39803 41037 39849 41075
rect 39803 41003 39809 41037
rect 39843 41003 39849 41037
rect 39803 40965 39849 41003
rect 39803 40931 39809 40965
rect 39843 40931 39849 40965
rect 39803 40893 39849 40931
rect 39803 40859 39809 40893
rect 39843 40859 39849 40893
rect 39803 40821 39849 40859
rect 39803 40787 39809 40821
rect 39843 40787 39849 40821
rect 39803 40749 39849 40787
rect 39803 40715 39809 40749
rect 39843 40715 39849 40749
rect 39803 40677 39849 40715
rect 39803 40643 39809 40677
rect 39843 40643 39849 40677
rect 39803 40605 39849 40643
rect 39803 40571 39809 40605
rect 39843 40571 39849 40605
rect 39803 40533 39849 40571
rect 39803 40499 39809 40533
rect 39843 40499 39849 40533
rect 39803 40461 39849 40499
rect 39803 40427 39809 40461
rect 39843 40427 39849 40461
rect 39803 40389 39849 40427
rect 39803 40355 39809 40389
rect 39843 40355 39849 40389
rect 39803 40317 39849 40355
rect 39803 40283 39809 40317
rect 39843 40283 39849 40317
rect 39803 40245 39849 40283
rect 39803 40211 39809 40245
rect 39843 40211 39849 40245
rect 39803 40173 39849 40211
rect 39803 40139 39809 40173
rect 39843 40139 39849 40173
rect 39803 40101 39849 40139
rect 39803 40067 39809 40101
rect 39843 40067 39849 40101
rect 39803 40029 39849 40067
rect 39803 39995 39809 40029
rect 39843 39995 39849 40029
rect 39803 39957 39849 39995
rect 39803 39923 39809 39957
rect 39843 39923 39849 39957
rect 39803 39907 39849 39923
rect 40261 41181 40307 41197
rect 40261 41147 40267 41181
rect 40301 41147 40307 41181
rect 40261 41109 40307 41147
rect 40261 41075 40267 41109
rect 40301 41075 40307 41109
rect 40261 41037 40307 41075
rect 40261 41003 40267 41037
rect 40301 41003 40307 41037
rect 40261 40965 40307 41003
rect 40261 40931 40267 40965
rect 40301 40931 40307 40965
rect 40261 40893 40307 40931
rect 40261 40859 40267 40893
rect 40301 40859 40307 40893
rect 40261 40821 40307 40859
rect 40261 40787 40267 40821
rect 40301 40787 40307 40821
rect 40261 40749 40307 40787
rect 40261 40715 40267 40749
rect 40301 40715 40307 40749
rect 40261 40677 40307 40715
rect 40261 40643 40267 40677
rect 40301 40643 40307 40677
rect 40261 40605 40307 40643
rect 40261 40571 40267 40605
rect 40301 40571 40307 40605
rect 40261 40533 40307 40571
rect 40261 40499 40267 40533
rect 40301 40499 40307 40533
rect 40261 40461 40307 40499
rect 40261 40427 40267 40461
rect 40301 40427 40307 40461
rect 40261 40389 40307 40427
rect 40261 40355 40267 40389
rect 40301 40355 40307 40389
rect 40261 40317 40307 40355
rect 40261 40283 40267 40317
rect 40301 40283 40307 40317
rect 40261 40245 40307 40283
rect 40261 40211 40267 40245
rect 40301 40211 40307 40245
rect 40261 40173 40307 40211
rect 40261 40139 40267 40173
rect 40301 40139 40307 40173
rect 40261 40101 40307 40139
rect 40261 40067 40267 40101
rect 40301 40067 40307 40101
rect 40261 40029 40307 40067
rect 40261 39995 40267 40029
rect 40301 39995 40307 40029
rect 40261 39957 40307 39995
rect 40261 39923 40267 39957
rect 40301 39923 40307 39957
rect 40261 39907 40307 39923
rect 40719 41181 40765 41197
rect 40719 41147 40725 41181
rect 40759 41147 40765 41181
rect 40719 41109 40765 41147
rect 40719 41075 40725 41109
rect 40759 41075 40765 41109
rect 40719 41037 40765 41075
rect 40719 41003 40725 41037
rect 40759 41003 40765 41037
rect 40719 40965 40765 41003
rect 40719 40931 40725 40965
rect 40759 40931 40765 40965
rect 40719 40893 40765 40931
rect 40719 40859 40725 40893
rect 40759 40859 40765 40893
rect 40719 40821 40765 40859
rect 40719 40787 40725 40821
rect 40759 40787 40765 40821
rect 40719 40749 40765 40787
rect 40719 40715 40725 40749
rect 40759 40715 40765 40749
rect 40719 40677 40765 40715
rect 40719 40643 40725 40677
rect 40759 40643 40765 40677
rect 40719 40605 40765 40643
rect 40719 40571 40725 40605
rect 40759 40571 40765 40605
rect 40719 40533 40765 40571
rect 40719 40499 40725 40533
rect 40759 40499 40765 40533
rect 40719 40461 40765 40499
rect 40719 40427 40725 40461
rect 40759 40427 40765 40461
rect 40719 40389 40765 40427
rect 40719 40355 40725 40389
rect 40759 40355 40765 40389
rect 40719 40317 40765 40355
rect 40719 40283 40725 40317
rect 40759 40283 40765 40317
rect 40719 40245 40765 40283
rect 40719 40211 40725 40245
rect 40759 40211 40765 40245
rect 40719 40173 40765 40211
rect 40719 40139 40725 40173
rect 40759 40139 40765 40173
rect 40719 40101 40765 40139
rect 40719 40067 40725 40101
rect 40759 40067 40765 40101
rect 40719 40029 40765 40067
rect 40719 39995 40725 40029
rect 40759 39995 40765 40029
rect 40719 39957 40765 39995
rect 40719 39923 40725 39957
rect 40759 39923 40765 39957
rect 40719 39907 40765 39923
rect 41177 41181 41223 41197
rect 41177 41147 41183 41181
rect 41217 41147 41223 41181
rect 41177 41109 41223 41147
rect 41177 41075 41183 41109
rect 41217 41075 41223 41109
rect 41177 41037 41223 41075
rect 41177 41003 41183 41037
rect 41217 41003 41223 41037
rect 41177 40965 41223 41003
rect 41177 40931 41183 40965
rect 41217 40931 41223 40965
rect 41177 40893 41223 40931
rect 41177 40859 41183 40893
rect 41217 40859 41223 40893
rect 41177 40821 41223 40859
rect 41177 40787 41183 40821
rect 41217 40787 41223 40821
rect 41177 40749 41223 40787
rect 41177 40715 41183 40749
rect 41217 40715 41223 40749
rect 41177 40677 41223 40715
rect 41177 40643 41183 40677
rect 41217 40643 41223 40677
rect 41177 40605 41223 40643
rect 41177 40571 41183 40605
rect 41217 40571 41223 40605
rect 41177 40533 41223 40571
rect 41177 40499 41183 40533
rect 41217 40499 41223 40533
rect 41177 40461 41223 40499
rect 41177 40427 41183 40461
rect 41217 40427 41223 40461
rect 41177 40389 41223 40427
rect 41177 40355 41183 40389
rect 41217 40355 41223 40389
rect 41177 40317 41223 40355
rect 41177 40283 41183 40317
rect 41217 40283 41223 40317
rect 41177 40245 41223 40283
rect 41177 40211 41183 40245
rect 41217 40211 41223 40245
rect 41177 40173 41223 40211
rect 41177 40139 41183 40173
rect 41217 40139 41223 40173
rect 41177 40101 41223 40139
rect 41177 40067 41183 40101
rect 41217 40067 41223 40101
rect 41177 40029 41223 40067
rect 41177 39995 41183 40029
rect 41217 39995 41223 40029
rect 41177 39957 41223 39995
rect 41177 39923 41183 39957
rect 41217 39923 41223 39957
rect 41177 39907 41223 39923
rect 41635 41181 41681 41197
rect 41635 41147 41641 41181
rect 41675 41147 41681 41181
rect 41635 41109 41681 41147
rect 41635 41075 41641 41109
rect 41675 41075 41681 41109
rect 41635 41037 41681 41075
rect 41635 41003 41641 41037
rect 41675 41003 41681 41037
rect 41635 40965 41681 41003
rect 41635 40931 41641 40965
rect 41675 40931 41681 40965
rect 41635 40893 41681 40931
rect 41635 40859 41641 40893
rect 41675 40859 41681 40893
rect 41635 40821 41681 40859
rect 41635 40787 41641 40821
rect 41675 40787 41681 40821
rect 41635 40749 41681 40787
rect 41635 40715 41641 40749
rect 41675 40715 41681 40749
rect 41635 40677 41681 40715
rect 41635 40643 41641 40677
rect 41675 40643 41681 40677
rect 41635 40605 41681 40643
rect 41635 40571 41641 40605
rect 41675 40571 41681 40605
rect 41635 40533 41681 40571
rect 41635 40499 41641 40533
rect 41675 40499 41681 40533
rect 41635 40461 41681 40499
rect 41635 40427 41641 40461
rect 41675 40427 41681 40461
rect 41635 40389 41681 40427
rect 41635 40355 41641 40389
rect 41675 40355 41681 40389
rect 41635 40317 41681 40355
rect 41635 40283 41641 40317
rect 41675 40283 41681 40317
rect 41635 40245 41681 40283
rect 41635 40211 41641 40245
rect 41675 40211 41681 40245
rect 41635 40173 41681 40211
rect 41635 40139 41641 40173
rect 41675 40139 41681 40173
rect 41635 40101 41681 40139
rect 41635 40067 41641 40101
rect 41675 40067 41681 40101
rect 41635 40029 41681 40067
rect 41635 39995 41641 40029
rect 41675 39995 41681 40029
rect 41635 39957 41681 39995
rect 41635 39923 41641 39957
rect 41675 39923 41681 39957
rect 41635 39907 41681 39923
rect 42093 41181 42139 41197
rect 42093 41147 42099 41181
rect 42133 41147 42139 41181
rect 42093 41109 42139 41147
rect 42093 41075 42099 41109
rect 42133 41075 42139 41109
rect 42093 41037 42139 41075
rect 42093 41003 42099 41037
rect 42133 41003 42139 41037
rect 42093 40965 42139 41003
rect 42093 40931 42099 40965
rect 42133 40931 42139 40965
rect 42093 40893 42139 40931
rect 42093 40859 42099 40893
rect 42133 40859 42139 40893
rect 42093 40821 42139 40859
rect 42093 40787 42099 40821
rect 42133 40787 42139 40821
rect 42093 40749 42139 40787
rect 42093 40715 42099 40749
rect 42133 40715 42139 40749
rect 42093 40677 42139 40715
rect 42093 40643 42099 40677
rect 42133 40643 42139 40677
rect 42093 40605 42139 40643
rect 42093 40571 42099 40605
rect 42133 40571 42139 40605
rect 42093 40533 42139 40571
rect 42093 40499 42099 40533
rect 42133 40499 42139 40533
rect 42093 40461 42139 40499
rect 42093 40427 42099 40461
rect 42133 40427 42139 40461
rect 42093 40389 42139 40427
rect 42093 40355 42099 40389
rect 42133 40355 42139 40389
rect 42093 40317 42139 40355
rect 42093 40283 42099 40317
rect 42133 40283 42139 40317
rect 42093 40245 42139 40283
rect 42093 40211 42099 40245
rect 42133 40211 42139 40245
rect 42093 40173 42139 40211
rect 42093 40139 42099 40173
rect 42133 40139 42139 40173
rect 42093 40101 42139 40139
rect 42093 40067 42099 40101
rect 42133 40067 42139 40101
rect 42093 40029 42139 40067
rect 42093 39995 42099 40029
rect 42133 39995 42139 40029
rect 42093 39957 42139 39995
rect 42093 39923 42099 39957
rect 42133 39923 42139 39957
rect 42093 39907 42139 39923
rect 42551 41181 42597 41197
rect 42551 41147 42557 41181
rect 42591 41147 42597 41181
rect 42551 41109 42597 41147
rect 42551 41075 42557 41109
rect 42591 41075 42597 41109
rect 42551 41037 42597 41075
rect 42551 41003 42557 41037
rect 42591 41003 42597 41037
rect 42551 40965 42597 41003
rect 42551 40931 42557 40965
rect 42591 40931 42597 40965
rect 42551 40893 42597 40931
rect 42551 40859 42557 40893
rect 42591 40859 42597 40893
rect 42551 40821 42597 40859
rect 42551 40787 42557 40821
rect 42591 40787 42597 40821
rect 42551 40749 42597 40787
rect 42551 40715 42557 40749
rect 42591 40715 42597 40749
rect 42551 40677 42597 40715
rect 42551 40643 42557 40677
rect 42591 40643 42597 40677
rect 42551 40605 42597 40643
rect 42551 40571 42557 40605
rect 42591 40571 42597 40605
rect 42551 40533 42597 40571
rect 42551 40499 42557 40533
rect 42591 40499 42597 40533
rect 42551 40461 42597 40499
rect 42551 40427 42557 40461
rect 42591 40427 42597 40461
rect 42551 40389 42597 40427
rect 42551 40355 42557 40389
rect 42591 40355 42597 40389
rect 42551 40317 42597 40355
rect 42551 40283 42557 40317
rect 42591 40283 42597 40317
rect 42551 40245 42597 40283
rect 42551 40211 42557 40245
rect 42591 40211 42597 40245
rect 42551 40173 42597 40211
rect 42551 40139 42557 40173
rect 42591 40139 42597 40173
rect 42551 40101 42597 40139
rect 42551 40067 42557 40101
rect 42591 40067 42597 40101
rect 42551 40029 42597 40067
rect 42551 39995 42557 40029
rect 42591 39995 42597 40029
rect 42551 39957 42597 39995
rect 42551 39923 42557 39957
rect 42591 39923 42597 39957
rect 42551 39907 42597 39923
rect 38654 39828 38660 39840
rect 38599 39800 38660 39828
rect 38654 39788 38660 39800
rect 38712 39788 38718 39840
rect 6457 39763 6515 39769
rect 6457 39729 6469 39763
rect 6503 39760 6515 39763
rect 6503 39732 9628 39760
rect 6503 39729 6515 39732
rect 6457 39723 6515 39729
rect 9600 39704 9628 39732
rect 9582 39652 9588 39704
rect 9640 39652 9646 39704
rect 15010 39692 15016 39704
rect 14955 39664 15016 39692
rect 15010 39652 15016 39664
rect 15068 39652 15074 39704
rect 27614 39692 27620 39704
rect 27559 39664 27620 39692
rect 27614 39652 27620 39664
rect 27672 39652 27678 39704
rect 900 39610 47736 39612
rect 900 39494 922 39610
rect 2510 39569 46126 39610
rect 2510 39535 6167 39569
rect 6201 39535 6983 39569
rect 7017 39535 7383 39569
rect 7417 39535 7783 39569
rect 7817 39535 8183 39569
rect 8217 39535 8583 39569
rect 8617 39535 8983 39569
rect 9017 39535 9383 39569
rect 9417 39535 9783 39569
rect 9817 39535 10183 39569
rect 10217 39535 10583 39569
rect 10617 39535 10983 39569
rect 11017 39535 11383 39569
rect 11417 39535 11783 39569
rect 11817 39535 12183 39569
rect 12217 39535 12583 39569
rect 12617 39535 12983 39569
rect 13017 39535 13383 39569
rect 13417 39535 13783 39569
rect 13817 39535 15213 39569
rect 15247 39535 15613 39569
rect 15647 39535 16013 39569
rect 16047 39535 16413 39569
rect 16447 39535 16813 39569
rect 16847 39535 17213 39569
rect 17247 39535 17613 39569
rect 17647 39535 18013 39569
rect 18047 39535 18413 39569
rect 18447 39535 18813 39569
rect 18847 39535 19213 39569
rect 19247 39535 19613 39569
rect 19647 39535 20013 39569
rect 20047 39535 20413 39569
rect 20447 39535 20813 39569
rect 20847 39535 21213 39569
rect 21247 39535 21613 39569
rect 21647 39535 22013 39569
rect 22047 39535 22413 39569
rect 22447 39535 22813 39569
rect 22847 39535 23213 39569
rect 23247 39535 23613 39569
rect 23647 39535 24013 39569
rect 24047 39535 24413 39569
rect 24447 39535 24813 39569
rect 24847 39535 25213 39569
rect 25247 39535 25613 39569
rect 25647 39535 26013 39569
rect 26047 39535 26413 39569
rect 26447 39535 26813 39569
rect 26847 39535 27213 39569
rect 27247 39535 27613 39569
rect 27647 39535 28013 39569
rect 28047 39535 28413 39569
rect 28447 39535 28813 39569
rect 28847 39535 29213 39569
rect 29247 39535 29613 39569
rect 29647 39535 30013 39569
rect 30047 39535 30413 39569
rect 30447 39535 30813 39569
rect 30847 39535 31213 39569
rect 31247 39535 31613 39569
rect 31647 39535 32013 39569
rect 32047 39535 32413 39569
rect 32447 39535 32813 39569
rect 32847 39535 33213 39569
rect 33247 39535 33613 39569
rect 33647 39535 34013 39569
rect 34047 39535 34413 39569
rect 34447 39535 34813 39569
rect 34847 39535 35213 39569
rect 35247 39535 35613 39569
rect 35647 39535 36013 39569
rect 36047 39535 36413 39569
rect 36447 39535 36813 39569
rect 36847 39535 37213 39569
rect 37247 39535 37613 39569
rect 37647 39535 38013 39569
rect 38047 39535 38413 39569
rect 38447 39535 38813 39569
rect 38847 39535 39213 39569
rect 39247 39535 39613 39569
rect 39647 39535 40013 39569
rect 40047 39535 40413 39569
rect 40447 39535 40813 39569
rect 40847 39535 41213 39569
rect 41247 39535 41613 39569
rect 41647 39535 42013 39569
rect 42047 39535 42413 39569
rect 42447 39535 46126 39569
rect 2510 39494 46126 39535
rect 47714 39494 47736 39610
rect 900 39492 47736 39494
rect 3348 37730 45288 37732
rect 3348 37614 3370 37730
rect 4958 37689 43678 37730
rect 4958 37655 6101 37689
rect 6135 37655 6501 37689
rect 6535 37655 6901 37689
rect 6935 37655 7301 37689
rect 7335 37655 7701 37689
rect 7735 37655 8101 37689
rect 8135 37655 8501 37689
rect 8535 37655 8901 37689
rect 8935 37655 9301 37689
rect 9335 37655 9701 37689
rect 9735 37655 10101 37689
rect 10135 37655 10501 37689
rect 10535 37655 10901 37689
rect 10935 37655 11301 37689
rect 11335 37655 11701 37689
rect 11735 37655 12101 37689
rect 12135 37655 12501 37689
rect 12535 37655 12901 37689
rect 12935 37664 13549 37689
rect 12935 37655 12992 37664
rect 4958 37614 12992 37655
rect 3348 37612 12992 37614
rect 13044 37655 13549 37664
rect 13583 37655 13949 37689
rect 13983 37655 14349 37689
rect 14383 37655 14749 37689
rect 14783 37655 15149 37689
rect 15183 37655 15549 37689
rect 15583 37655 15949 37689
rect 15983 37655 16349 37689
rect 16383 37655 16749 37689
rect 16783 37664 17149 37689
rect 16783 37655 16856 37664
rect 13044 37612 16856 37655
rect 16908 37655 17149 37664
rect 17183 37655 17549 37689
rect 17583 37655 17949 37689
rect 17983 37655 18349 37689
rect 18383 37655 18749 37689
rect 18783 37655 19149 37689
rect 19183 37655 19549 37689
rect 19583 37655 19949 37689
rect 19983 37655 20349 37689
rect 20383 37655 20997 37689
rect 21031 37655 21397 37689
rect 21431 37655 21797 37689
rect 21831 37655 22197 37689
rect 22231 37655 22597 37689
rect 22631 37655 22997 37689
rect 23031 37655 23397 37689
rect 23431 37655 23797 37689
rect 23831 37655 24197 37689
rect 24231 37655 24597 37689
rect 24631 37655 24997 37689
rect 25031 37655 25397 37689
rect 25431 37655 25797 37689
rect 25831 37655 26197 37689
rect 26231 37655 26597 37689
rect 26631 37655 26997 37689
rect 27031 37655 27397 37689
rect 27431 37655 27797 37689
rect 27831 37664 28511 37689
rect 27831 37655 27896 37664
rect 16908 37612 27896 37655
rect 27948 37655 28511 37664
rect 28545 37655 30207 37689
rect 30241 37655 30407 37689
rect 30441 37655 30607 37689
rect 30641 37655 30807 37689
rect 30841 37655 31007 37689
rect 31041 37655 31207 37689
rect 31241 37655 31407 37689
rect 31441 37655 31607 37689
rect 31641 37655 31807 37689
rect 31841 37655 32007 37689
rect 32041 37655 32207 37689
rect 32241 37655 32407 37689
rect 32441 37655 32607 37689
rect 32641 37655 32807 37689
rect 32841 37655 33007 37689
rect 33041 37655 33207 37689
rect 33241 37655 33407 37689
rect 33441 37655 33607 37689
rect 33641 37655 33807 37689
rect 33841 37655 34007 37689
rect 34041 37655 34207 37689
rect 34241 37655 34407 37689
rect 34441 37655 34607 37689
rect 34641 37655 34807 37689
rect 34841 37655 35007 37689
rect 35041 37655 35207 37689
rect 35241 37655 35407 37689
rect 35441 37655 35607 37689
rect 35641 37655 35807 37689
rect 35841 37655 36007 37689
rect 36041 37655 36207 37689
rect 36241 37655 36407 37689
rect 36441 37655 36607 37689
rect 36641 37655 36807 37689
rect 36841 37655 37007 37689
rect 37041 37655 37207 37689
rect 37241 37655 37407 37689
rect 37441 37655 37607 37689
rect 37641 37655 37807 37689
rect 37841 37655 38007 37689
rect 38041 37655 38207 37689
rect 38241 37655 38407 37689
rect 38441 37655 38607 37689
rect 38641 37655 38807 37689
rect 38841 37655 39007 37689
rect 39041 37655 39207 37689
rect 39241 37655 39929 37689
rect 39963 37655 40129 37689
rect 40163 37655 40329 37689
rect 40363 37655 40529 37689
rect 40563 37655 40729 37689
rect 40763 37655 40929 37689
rect 40963 37655 41129 37689
rect 41163 37655 41329 37689
rect 41363 37655 41529 37689
rect 41563 37655 41729 37689
rect 41763 37655 41929 37689
rect 41963 37655 43678 37689
rect 27948 37614 43678 37655
rect 45266 37614 45288 37730
rect 27948 37612 45288 37614
rect 28813 37519 28871 37525
rect 28813 37485 28825 37519
rect 28859 37485 28871 37519
rect 28813 37479 28871 37485
rect 28828 37380 28856 37479
rect 39757 37421 40167 37433
rect 28828 37362 30144 37380
rect 28828 37356 39378 37362
rect 28828 37352 30070 37356
rect 30050 37322 30070 37352
rect 30104 37322 30160 37356
rect 30194 37322 30250 37356
rect 30284 37322 30340 37356
rect 30374 37322 30430 37356
rect 30464 37322 30520 37356
rect 30554 37322 30610 37356
rect 30644 37322 30700 37356
rect 30734 37322 30790 37356
rect 30824 37322 30880 37356
rect 30914 37322 30970 37356
rect 31004 37322 31060 37356
rect 31094 37322 31150 37356
rect 31184 37322 31240 37356
rect 31274 37322 31410 37356
rect 31444 37322 31500 37356
rect 31534 37322 31590 37356
rect 31624 37322 31680 37356
rect 31714 37322 31770 37356
rect 31804 37322 31860 37356
rect 31894 37322 31950 37356
rect 31984 37322 32040 37356
rect 32074 37322 32130 37356
rect 32164 37322 32220 37356
rect 32254 37322 32310 37356
rect 32344 37322 32400 37356
rect 32434 37322 32490 37356
rect 32524 37322 32580 37356
rect 32614 37322 32750 37356
rect 32784 37322 32840 37356
rect 32874 37322 32930 37356
rect 32964 37322 33020 37356
rect 33054 37322 33110 37356
rect 33144 37322 33200 37356
rect 33234 37322 33290 37356
rect 33324 37322 33380 37356
rect 33414 37322 33470 37356
rect 33504 37322 33560 37356
rect 33594 37322 33650 37356
rect 33684 37322 33740 37356
rect 33774 37322 33830 37356
rect 33864 37322 33920 37356
rect 33954 37322 34090 37356
rect 34124 37322 34180 37356
rect 34214 37322 34270 37356
rect 34304 37322 34360 37356
rect 34394 37322 34450 37356
rect 34484 37322 34540 37356
rect 34574 37322 34630 37356
rect 34664 37322 34720 37356
rect 34754 37322 34810 37356
rect 34844 37322 34900 37356
rect 34934 37322 34990 37356
rect 35024 37322 35080 37356
rect 35114 37322 35170 37356
rect 35204 37322 35260 37356
rect 35294 37322 35430 37356
rect 35464 37322 35520 37356
rect 35554 37322 35610 37356
rect 35644 37322 35700 37356
rect 35734 37322 35790 37356
rect 35824 37322 35880 37356
rect 35914 37322 35970 37356
rect 36004 37322 36060 37356
rect 36094 37322 36150 37356
rect 36184 37322 36240 37356
rect 36274 37322 36330 37356
rect 36364 37322 36420 37356
rect 36454 37322 36510 37356
rect 36544 37322 36600 37356
rect 36634 37322 36770 37356
rect 36804 37322 36860 37356
rect 36894 37322 36950 37356
rect 36984 37322 37040 37356
rect 37074 37322 37130 37356
rect 37164 37322 37220 37356
rect 37254 37322 37310 37356
rect 37344 37322 37400 37356
rect 37434 37322 37490 37356
rect 37524 37322 37580 37356
rect 37614 37322 37670 37356
rect 37704 37322 37760 37356
rect 37794 37322 37850 37356
rect 37884 37322 37940 37356
rect 37974 37322 38110 37356
rect 38144 37322 38200 37356
rect 38234 37322 38290 37356
rect 38324 37322 38380 37356
rect 38414 37322 38470 37356
rect 38504 37322 38560 37356
rect 38594 37322 38650 37356
rect 38684 37322 38740 37356
rect 38774 37322 38830 37356
rect 38864 37322 38920 37356
rect 38954 37322 39010 37356
rect 39044 37322 39100 37356
rect 39134 37322 39190 37356
rect 39224 37322 39280 37356
rect 39314 37322 39378 37356
rect 30050 37292 39378 37322
rect 28334 37169 28380 37192
rect 28334 37135 28340 37169
rect 28374 37135 28380 37169
rect 28334 37097 28380 37135
rect 28334 37063 28340 37097
rect 28374 37063 28380 37097
rect 28334 37025 28380 37063
rect 28334 36991 28340 37025
rect 28374 36991 28380 37025
rect 28334 36953 28380 36991
rect 28334 36919 28340 36953
rect 28374 36919 28380 36953
rect 28334 36881 28380 36919
rect 28334 36847 28340 36881
rect 28374 36847 28380 36881
rect 28334 36809 28380 36847
rect 28334 36775 28340 36809
rect 28374 36775 28380 36809
rect 28334 36737 28380 36775
rect 28334 36703 28340 36737
rect 28374 36703 28380 36737
rect 28334 36665 28380 36703
rect 28334 36631 28340 36665
rect 28374 36631 28380 36665
rect 28334 36593 28380 36631
rect 28334 36559 28340 36593
rect 28374 36559 28380 36593
rect 28334 36521 28380 36559
rect 28334 36487 28340 36521
rect 28374 36487 28380 36521
rect 28334 36449 28380 36487
rect 28334 36415 28340 36449
rect 28374 36415 28380 36449
rect 28334 36392 28380 36415
rect 28792 37169 28838 37192
rect 28792 37135 28798 37169
rect 28832 37135 28838 37169
rect 30116 37176 30144 37292
rect 30214 37196 39214 37212
rect 30214 37188 30234 37196
rect 30190 37176 30196 37188
rect 30116 37148 30196 37176
rect 30268 37162 30324 37196
rect 30358 37162 30414 37196
rect 30448 37162 30504 37196
rect 30538 37162 30594 37196
rect 30628 37162 30684 37196
rect 30718 37162 30774 37196
rect 30808 37162 30864 37196
rect 30898 37162 30954 37196
rect 30988 37162 31044 37196
rect 31078 37162 31134 37196
rect 31168 37162 31574 37196
rect 31608 37162 31664 37196
rect 31698 37162 31754 37196
rect 31788 37162 31844 37196
rect 31878 37162 31934 37196
rect 31968 37162 32024 37196
rect 32058 37162 32114 37196
rect 32148 37162 32204 37196
rect 32238 37162 32294 37196
rect 32328 37162 32384 37196
rect 32418 37162 32474 37196
rect 32508 37162 32914 37196
rect 32948 37162 33004 37196
rect 33038 37162 33094 37196
rect 33128 37162 33184 37196
rect 33218 37162 33274 37196
rect 33308 37162 33364 37196
rect 33398 37162 33454 37196
rect 33488 37162 33544 37196
rect 33578 37162 33634 37196
rect 33668 37162 33724 37196
rect 33758 37162 33814 37196
rect 33848 37162 34254 37196
rect 34288 37162 34344 37196
rect 34378 37162 34434 37196
rect 34468 37162 34524 37196
rect 34558 37162 34614 37196
rect 34648 37162 34704 37196
rect 34738 37162 34794 37196
rect 34828 37162 34884 37196
rect 34918 37162 34974 37196
rect 35008 37162 35064 37196
rect 35098 37162 35154 37196
rect 35188 37162 35594 37196
rect 35628 37162 35684 37196
rect 35718 37162 35774 37196
rect 35808 37162 35864 37196
rect 35898 37162 35954 37196
rect 35988 37162 36044 37196
rect 36078 37162 36134 37196
rect 36168 37162 36224 37196
rect 36258 37162 36314 37196
rect 36348 37162 36404 37196
rect 36438 37162 36494 37196
rect 36528 37162 36934 37196
rect 36968 37162 37024 37196
rect 37058 37162 37114 37196
rect 37148 37162 37204 37196
rect 37238 37162 37294 37196
rect 37328 37162 37384 37196
rect 37418 37162 37474 37196
rect 37508 37162 37564 37196
rect 37598 37162 37654 37196
rect 37688 37162 37744 37196
rect 37778 37162 37834 37196
rect 37868 37162 38274 37196
rect 38308 37162 38364 37196
rect 38398 37162 38454 37196
rect 38488 37162 38544 37196
rect 38578 37162 38634 37196
rect 38668 37162 38724 37196
rect 38758 37162 38814 37196
rect 38848 37162 38904 37196
rect 38938 37162 38994 37196
rect 39028 37162 39084 37196
rect 39118 37162 39174 37196
rect 39208 37162 39214 37196
rect 30190 37136 30196 37148
rect 30248 37142 39214 37162
rect 30248 37136 30254 37142
rect 28792 37097 28838 37135
rect 28792 37063 28798 37097
rect 28832 37063 28838 37097
rect 28792 37025 28838 37063
rect 28792 36991 28798 37025
rect 28832 36991 28838 37025
rect 28792 36953 28838 36991
rect 28792 36919 28798 36953
rect 28832 36919 28838 36953
rect 28792 36881 28838 36919
rect 28792 36847 28798 36881
rect 28832 36847 28838 36881
rect 28792 36809 28838 36847
rect 28792 36775 28798 36809
rect 28832 36775 28838 36809
rect 28792 36737 28838 36775
rect 28792 36703 28798 36737
rect 28832 36703 28838 36737
rect 28792 36665 28838 36703
rect 28792 36631 28798 36665
rect 28832 36631 28838 36665
rect 28792 36593 28838 36631
rect 28792 36559 28798 36593
rect 28832 36559 28838 36593
rect 28792 36521 28838 36559
rect 28792 36487 28798 36521
rect 28832 36487 28838 36521
rect 28792 36449 28838 36487
rect 28792 36415 28798 36449
rect 28832 36415 28838 36449
rect 30388 36992 39040 37038
rect 30388 36958 30420 36992
rect 30454 36958 30520 36992
rect 30554 36958 30620 36992
rect 30654 36958 30720 36992
rect 30754 36958 30820 36992
rect 30854 36958 30920 36992
rect 30954 36958 31760 36992
rect 31794 36958 31860 36992
rect 31894 36958 31960 36992
rect 31994 36958 32060 36992
rect 32094 36958 32160 36992
rect 32194 36958 32260 36992
rect 32294 36958 33100 36992
rect 33134 36958 33200 36992
rect 33234 36958 33300 36992
rect 33334 36958 33400 36992
rect 33434 36958 33500 36992
rect 33534 36958 33600 36992
rect 33634 36958 34440 36992
rect 34474 36958 34540 36992
rect 34574 36958 34640 36992
rect 34674 36958 34740 36992
rect 34774 36958 34840 36992
rect 34874 36958 34940 36992
rect 34974 36958 35780 36992
rect 35814 36958 35880 36992
rect 35914 36958 35980 36992
rect 36014 36958 36080 36992
rect 36114 36958 36180 36992
rect 36214 36958 36280 36992
rect 36314 36958 37120 36992
rect 37154 36958 37220 36992
rect 37254 36958 37320 36992
rect 37354 36958 37420 36992
rect 37454 36958 37520 36992
rect 37554 36958 37620 36992
rect 37654 36958 38460 36992
rect 38494 36958 38560 36992
rect 38594 36958 38660 36992
rect 38694 36958 38760 36992
rect 38794 36958 38860 36992
rect 38894 36958 38960 36992
rect 38994 36958 39040 36992
rect 30388 36892 39040 36958
rect 30388 36858 30420 36892
rect 30454 36858 30520 36892
rect 30554 36858 30620 36892
rect 30654 36858 30720 36892
rect 30754 36858 30820 36892
rect 30854 36858 30920 36892
rect 30954 36858 31760 36892
rect 31794 36858 31860 36892
rect 31894 36858 31960 36892
rect 31994 36858 32060 36892
rect 32094 36858 32160 36892
rect 32194 36858 32260 36892
rect 32294 36858 33100 36892
rect 33134 36858 33200 36892
rect 33234 36858 33300 36892
rect 33334 36858 33400 36892
rect 33434 36858 33500 36892
rect 33534 36858 33600 36892
rect 33634 36858 34440 36892
rect 34474 36858 34540 36892
rect 34574 36858 34640 36892
rect 34674 36858 34740 36892
rect 34774 36858 34840 36892
rect 34874 36858 34940 36892
rect 34974 36858 35780 36892
rect 35814 36858 35880 36892
rect 35914 36858 35980 36892
rect 36014 36858 36080 36892
rect 36114 36858 36180 36892
rect 36214 36858 36280 36892
rect 36314 36858 37120 36892
rect 37154 36858 37220 36892
rect 37254 36858 37320 36892
rect 37354 36858 37420 36892
rect 37454 36858 37520 36892
rect 37554 36858 37620 36892
rect 37654 36858 38460 36892
rect 38494 36858 38560 36892
rect 38594 36858 38660 36892
rect 38694 36858 38760 36892
rect 38794 36858 38860 36892
rect 38894 36858 38960 36892
rect 38994 36858 39040 36892
rect 39757 36883 39765 37421
rect 40159 36883 40167 37421
rect 39757 36871 40167 36883
rect 41765 37421 42175 37433
rect 41765 36883 41772 37421
rect 42166 36883 42175 37421
rect 41765 36871 42175 36883
rect 30388 36792 39040 36858
rect 30388 36758 30420 36792
rect 30454 36758 30520 36792
rect 30554 36758 30620 36792
rect 30654 36758 30720 36792
rect 30754 36758 30820 36792
rect 30854 36758 30920 36792
rect 30954 36758 31760 36792
rect 31794 36758 31860 36792
rect 31894 36758 31960 36792
rect 31994 36758 32060 36792
rect 32094 36758 32160 36792
rect 32194 36758 32260 36792
rect 32294 36758 33100 36792
rect 33134 36758 33200 36792
rect 33234 36758 33300 36792
rect 33334 36758 33400 36792
rect 33434 36758 33500 36792
rect 33534 36758 33600 36792
rect 33634 36758 34440 36792
rect 34474 36758 34540 36792
rect 34574 36758 34640 36792
rect 34674 36758 34740 36792
rect 34774 36758 34840 36792
rect 34874 36758 34940 36792
rect 34974 36758 35780 36792
rect 35814 36758 35880 36792
rect 35914 36758 35980 36792
rect 36014 36758 36080 36792
rect 36114 36758 36180 36792
rect 36214 36758 36280 36792
rect 36314 36758 37120 36792
rect 37154 36758 37220 36792
rect 37254 36758 37320 36792
rect 37354 36758 37420 36792
rect 37454 36758 37520 36792
rect 37554 36758 37620 36792
rect 37654 36758 38460 36792
rect 38494 36758 38560 36792
rect 38594 36758 38660 36792
rect 38694 36758 38760 36792
rect 38794 36758 38860 36792
rect 38894 36758 38960 36792
rect 38994 36758 39040 36792
rect 39960 36780 39988 36871
rect 30388 36692 39040 36758
rect 39942 36728 39948 36780
rect 40000 36728 40006 36780
rect 30388 36658 30420 36692
rect 30454 36658 30520 36692
rect 30554 36658 30620 36692
rect 30654 36658 30720 36692
rect 30754 36658 30820 36692
rect 30854 36658 30920 36692
rect 30954 36658 31760 36692
rect 31794 36658 31860 36692
rect 31894 36658 31960 36692
rect 31994 36658 32060 36692
rect 32094 36658 32160 36692
rect 32194 36658 32260 36692
rect 32294 36658 33100 36692
rect 33134 36658 33200 36692
rect 33234 36658 33300 36692
rect 33334 36658 33400 36692
rect 33434 36658 33500 36692
rect 33534 36658 33600 36692
rect 33634 36658 34440 36692
rect 34474 36658 34540 36692
rect 34574 36658 34640 36692
rect 34674 36658 34740 36692
rect 34774 36658 34840 36692
rect 34874 36658 34940 36692
rect 34974 36658 35780 36692
rect 35814 36658 35880 36692
rect 35914 36658 35980 36692
rect 36014 36658 36080 36692
rect 36114 36658 36180 36692
rect 36214 36658 36280 36692
rect 36314 36658 37120 36692
rect 37154 36658 37220 36692
rect 37254 36658 37320 36692
rect 37354 36658 37420 36692
rect 37454 36658 37520 36692
rect 37554 36658 37620 36692
rect 37654 36658 38460 36692
rect 38494 36658 38560 36692
rect 38594 36658 38660 36692
rect 38694 36658 38760 36692
rect 38794 36658 38860 36692
rect 38894 36658 38960 36692
rect 38994 36658 39040 36692
rect 30388 36592 39040 36658
rect 30388 36558 30420 36592
rect 30454 36558 30520 36592
rect 30554 36558 30620 36592
rect 30654 36558 30720 36592
rect 30754 36558 30820 36592
rect 30854 36558 30920 36592
rect 30954 36558 31760 36592
rect 31794 36558 31860 36592
rect 31894 36558 31960 36592
rect 31994 36558 32060 36592
rect 32094 36558 32160 36592
rect 32194 36558 32260 36592
rect 32294 36558 33100 36592
rect 33134 36558 33200 36592
rect 33234 36558 33300 36592
rect 33334 36558 33400 36592
rect 33434 36558 33500 36592
rect 33534 36558 33600 36592
rect 33634 36558 34440 36592
rect 34474 36558 34540 36592
rect 34574 36558 34640 36592
rect 34674 36558 34740 36592
rect 34774 36558 34840 36592
rect 34874 36558 34940 36592
rect 34974 36558 35780 36592
rect 35814 36558 35880 36592
rect 35914 36558 35980 36592
rect 36014 36558 36080 36592
rect 36114 36558 36180 36592
rect 36214 36558 36280 36592
rect 36314 36558 37120 36592
rect 37154 36558 37220 36592
rect 37254 36558 37320 36592
rect 37354 36558 37420 36592
rect 37454 36558 37520 36592
rect 37554 36558 37620 36592
rect 37654 36558 38460 36592
rect 38494 36558 38560 36592
rect 38594 36558 38660 36592
rect 38694 36558 38760 36592
rect 38794 36558 38860 36592
rect 38894 36558 38960 36592
rect 38994 36558 39040 36592
rect 30388 36508 39040 36558
rect 30388 36492 31668 36508
rect 30388 36458 30420 36492
rect 30454 36458 30520 36492
rect 30554 36458 30620 36492
rect 30654 36458 30720 36492
rect 30754 36458 30820 36492
rect 30854 36458 30920 36492
rect 30954 36458 31668 36492
rect 30388 36456 31668 36458
rect 31720 36496 39040 36508
rect 31720 36492 39344 36496
rect 31720 36458 31760 36492
rect 31794 36458 31860 36492
rect 31894 36458 31960 36492
rect 31994 36458 32060 36492
rect 32094 36458 32160 36492
rect 32194 36458 32260 36492
rect 32294 36458 33100 36492
rect 33134 36458 33200 36492
rect 33234 36458 33300 36492
rect 33334 36458 33400 36492
rect 33434 36458 33500 36492
rect 33534 36458 33600 36492
rect 33634 36458 34440 36492
rect 34474 36458 34540 36492
rect 34574 36458 34640 36492
rect 34674 36458 34740 36492
rect 34774 36458 34840 36492
rect 34874 36458 34940 36492
rect 34974 36458 35780 36492
rect 35814 36458 35880 36492
rect 35914 36458 35980 36492
rect 36014 36458 36080 36492
rect 36114 36458 36180 36492
rect 36214 36458 36280 36492
rect 36314 36458 37120 36492
rect 37154 36458 37220 36492
rect 37254 36458 37320 36492
rect 37354 36458 37420 36492
rect 37454 36458 37520 36492
rect 37554 36458 37620 36492
rect 37654 36458 38460 36492
rect 38494 36458 38560 36492
rect 38594 36458 38660 36492
rect 38694 36458 38760 36492
rect 38794 36458 38860 36492
rect 38894 36458 38960 36492
rect 38994 36468 39344 36492
rect 38994 36458 39040 36468
rect 31720 36456 39040 36458
rect 30388 36426 39040 36456
rect 39316 36428 39344 36468
rect 39757 36461 40167 36473
rect 39757 36428 39765 36461
rect 28792 36392 28838 36415
rect 39316 36400 39765 36428
rect 28353 36227 28411 36233
rect 28353 36224 28365 36227
rect 26252 36196 28365 36224
rect 26252 36168 26280 36196
rect 28353 36193 28365 36196
rect 28399 36193 28411 36227
rect 28353 36187 28411 36193
rect 26234 36116 26240 36168
rect 26292 36116 26298 36168
rect 9582 36048 9588 36100
rect 9640 36088 9646 36100
rect 9640 36060 28488 36088
rect 9640 36048 9646 36060
rect 28460 35961 28488 36060
rect 28445 35955 28503 35961
rect 28445 35921 28457 35955
rect 28491 35921 28503 35955
rect 28445 35915 28503 35921
rect 39757 35923 39765 36400
rect 40159 35923 40167 36461
rect 39757 35911 40167 35923
rect 41754 36461 42186 36871
rect 41754 35923 41772 36461
rect 42166 35923 42186 36461
rect 41754 35907 42186 35923
rect 900 35850 47736 35852
rect 900 35734 922 35850
rect 2510 35828 46126 35850
rect 2510 35809 30196 35828
rect 30248 35809 46126 35828
rect 2510 35775 6101 35809
rect 6135 35775 6501 35809
rect 6535 35775 6901 35809
rect 6935 35775 7301 35809
rect 7335 35775 7701 35809
rect 7735 35775 8101 35809
rect 8135 35775 8501 35809
rect 8535 35775 8901 35809
rect 8935 35775 9301 35809
rect 9335 35775 9701 35809
rect 9735 35775 10101 35809
rect 10135 35775 10501 35809
rect 10535 35775 10901 35809
rect 10935 35775 11301 35809
rect 11335 35775 11701 35809
rect 11735 35775 12101 35809
rect 12135 35775 12501 35809
rect 12535 35775 12901 35809
rect 12935 35775 13549 35809
rect 13583 35775 13949 35809
rect 13983 35775 14349 35809
rect 14383 35775 14749 35809
rect 14783 35775 15149 35809
rect 15183 35775 15549 35809
rect 15583 35775 15949 35809
rect 15983 35775 16349 35809
rect 16383 35775 16749 35809
rect 16783 35775 17149 35809
rect 17183 35775 17549 35809
rect 17583 35775 17949 35809
rect 17983 35775 18349 35809
rect 18383 35775 18749 35809
rect 18783 35775 19149 35809
rect 19183 35775 19549 35809
rect 19583 35775 19949 35809
rect 19983 35775 20349 35809
rect 20383 35775 20997 35809
rect 21031 35775 21397 35809
rect 21431 35775 21797 35809
rect 21831 35775 22197 35809
rect 22231 35775 22597 35809
rect 22631 35775 22997 35809
rect 23031 35775 23397 35809
rect 23431 35775 23797 35809
rect 23831 35775 24197 35809
rect 24231 35775 24597 35809
rect 24631 35775 24997 35809
rect 25031 35775 25397 35809
rect 25431 35775 25797 35809
rect 25831 35775 26197 35809
rect 26231 35775 26597 35809
rect 26631 35775 26997 35809
rect 27031 35775 27397 35809
rect 27431 35775 27797 35809
rect 27831 35775 28511 35809
rect 28545 35776 30196 35809
rect 30248 35776 30407 35809
rect 28545 35775 30207 35776
rect 30241 35775 30407 35776
rect 30441 35775 30607 35809
rect 30641 35775 30807 35809
rect 30841 35775 31007 35809
rect 31041 35775 31207 35809
rect 31241 35775 31407 35809
rect 31441 35775 31607 35809
rect 31641 35775 31807 35809
rect 31841 35775 32007 35809
rect 32041 35775 32207 35809
rect 32241 35775 32407 35809
rect 32441 35775 32607 35809
rect 32641 35775 32807 35809
rect 32841 35775 33007 35809
rect 33041 35775 33207 35809
rect 33241 35775 33407 35809
rect 33441 35775 33607 35809
rect 33641 35775 33807 35809
rect 33841 35775 34007 35809
rect 34041 35775 34207 35809
rect 34241 35775 34407 35809
rect 34441 35775 34607 35809
rect 34641 35775 34807 35809
rect 34841 35775 35007 35809
rect 35041 35775 35207 35809
rect 35241 35775 35407 35809
rect 35441 35775 35607 35809
rect 35641 35775 35807 35809
rect 35841 35775 36007 35809
rect 36041 35775 36207 35809
rect 36241 35775 36407 35809
rect 36441 35775 36607 35809
rect 36641 35775 36807 35809
rect 36841 35775 37007 35809
rect 37041 35775 37207 35809
rect 37241 35775 37407 35809
rect 37441 35775 37607 35809
rect 37641 35775 37807 35809
rect 37841 35775 38007 35809
rect 38041 35775 38207 35809
rect 38241 35775 38407 35809
rect 38441 35775 38607 35809
rect 38641 35775 38807 35809
rect 38841 35775 39007 35809
rect 39041 35775 39207 35809
rect 39241 35775 39929 35809
rect 39963 35775 40129 35809
rect 40163 35775 40329 35809
rect 40363 35775 40529 35809
rect 40563 35775 40729 35809
rect 40763 35775 40929 35809
rect 40963 35775 41129 35809
rect 41163 35775 41329 35809
rect 41363 35775 41529 35809
rect 41563 35775 41729 35809
rect 41763 35775 41929 35809
rect 41963 35775 46126 35809
rect 2510 35734 46126 35775
rect 47714 35734 47736 35850
rect 900 35732 47736 35734
rect 3348 33970 45288 33972
rect 3348 33854 3370 33970
rect 4958 33929 43678 33970
rect 4958 33895 6787 33929
rect 6821 33895 7187 33929
rect 7221 33895 7587 33929
rect 7621 33895 7987 33929
rect 8021 33895 8387 33929
rect 8421 33895 8787 33929
rect 8821 33895 9187 33929
rect 9221 33895 9587 33929
rect 9621 33924 9987 33929
rect 9621 33895 9956 33924
rect 10021 33895 10387 33929
rect 10421 33895 10787 33929
rect 10821 33895 11187 33929
rect 11221 33895 11587 33929
rect 11621 33895 11987 33929
rect 12021 33895 12387 33929
rect 12421 33895 12787 33929
rect 12821 33895 13187 33929
rect 13221 33895 13587 33929
rect 13621 33895 14331 33929
rect 14365 33895 14731 33929
rect 14765 33895 15131 33929
rect 15165 33895 15531 33929
rect 15565 33895 15931 33929
rect 15965 33895 16331 33929
rect 16365 33895 16731 33929
rect 16765 33895 17131 33929
rect 17165 33895 17531 33929
rect 17565 33895 17931 33929
rect 17965 33895 18331 33929
rect 18365 33895 18731 33929
rect 18765 33895 19131 33929
rect 19165 33895 19531 33929
rect 19565 33895 19931 33929
rect 19965 33895 20331 33929
rect 20365 33895 20731 33929
rect 20765 33895 21131 33929
rect 21165 33895 21531 33929
rect 21565 33895 21931 33929
rect 21965 33895 22331 33929
rect 22365 33895 22731 33929
rect 22765 33895 23131 33929
rect 23165 33895 23531 33929
rect 23565 33895 23931 33929
rect 23965 33895 24331 33929
rect 24365 33895 24731 33929
rect 24765 33895 25131 33929
rect 25165 33895 25531 33929
rect 25565 33895 25931 33929
rect 25965 33895 26331 33929
rect 26365 33895 26731 33929
rect 26765 33895 27131 33929
rect 27165 33895 27531 33929
rect 27565 33895 27931 33929
rect 27965 33895 28331 33929
rect 28365 33895 28731 33929
rect 28765 33895 29131 33929
rect 29165 33895 29531 33929
rect 29565 33895 29931 33929
rect 29965 33895 30331 33929
rect 30365 33895 30731 33929
rect 30765 33895 31131 33929
rect 31165 33895 31531 33929
rect 31565 33895 31931 33929
rect 31965 33895 32331 33929
rect 32365 33895 32731 33929
rect 32765 33895 33131 33929
rect 33165 33895 33531 33929
rect 33565 33895 33931 33929
rect 33965 33895 34331 33929
rect 34365 33895 34731 33929
rect 34765 33895 35131 33929
rect 35165 33895 35531 33929
rect 35565 33895 35931 33929
rect 35965 33895 36331 33929
rect 36365 33895 36731 33929
rect 36765 33895 37131 33929
rect 37165 33895 37531 33929
rect 37565 33895 37931 33929
rect 37965 33895 38331 33929
rect 38365 33895 38731 33929
rect 38765 33895 39131 33929
rect 39165 33895 39531 33929
rect 39565 33895 39931 33929
rect 39965 33895 40331 33929
rect 40365 33895 40731 33929
rect 40765 33895 41131 33929
rect 41165 33895 41531 33929
rect 41565 33895 43678 33929
rect 4958 33872 9956 33895
rect 10008 33872 43678 33895
rect 4958 33854 43678 33872
rect 45266 33854 45288 33970
rect 3348 33852 45288 33854
rect 14660 33677 14688 33852
rect 14189 33661 14235 33677
rect 14189 33627 14195 33661
rect 14229 33627 14235 33661
rect 14189 33589 14235 33627
rect 14189 33555 14195 33589
rect 14229 33555 14235 33589
rect 14189 33517 14235 33555
rect 14189 33483 14195 33517
rect 14229 33483 14235 33517
rect 14189 33445 14235 33483
rect 14189 33411 14195 33445
rect 14229 33411 14235 33445
rect 14189 33373 14235 33411
rect 14189 33339 14195 33373
rect 14229 33339 14235 33373
rect 14189 33301 14235 33339
rect 14189 33267 14195 33301
rect 14229 33267 14235 33301
rect 14189 33229 14235 33267
rect 14189 33195 14195 33229
rect 14229 33195 14235 33229
rect 14189 33157 14235 33195
rect 14189 33123 14195 33157
rect 14229 33123 14235 33157
rect 14189 33085 14235 33123
rect 14189 33051 14195 33085
rect 14229 33051 14235 33085
rect 14189 33013 14235 33051
rect 14189 32979 14195 33013
rect 14229 32979 14235 33013
rect 14189 32941 14235 32979
rect 14189 32907 14195 32941
rect 14229 32907 14235 32941
rect 14189 32869 14235 32907
rect 14189 32835 14195 32869
rect 14229 32835 14235 32869
rect 14189 32797 14235 32835
rect 14189 32763 14195 32797
rect 14229 32763 14235 32797
rect 14189 32725 14235 32763
rect 14189 32691 14195 32725
rect 14229 32691 14235 32725
rect 14189 32653 14235 32691
rect 14189 32619 14195 32653
rect 14229 32619 14235 32653
rect 14189 32581 14235 32619
rect 14189 32547 14195 32581
rect 14229 32547 14235 32581
rect 14189 32509 14235 32547
rect 14189 32475 14195 32509
rect 14229 32475 14235 32509
rect 14189 32437 14235 32475
rect 14189 32403 14195 32437
rect 14229 32403 14235 32437
rect 14189 32387 14235 32403
rect 14647 33661 14693 33677
rect 14647 33627 14653 33661
rect 14687 33627 14693 33661
rect 14647 33589 14693 33627
rect 14647 33555 14653 33589
rect 14687 33555 14693 33589
rect 14647 33517 14693 33555
rect 14647 33483 14653 33517
rect 14687 33483 14693 33517
rect 14647 33445 14693 33483
rect 14647 33411 14653 33445
rect 14687 33411 14693 33445
rect 14647 33373 14693 33411
rect 14647 33339 14653 33373
rect 14687 33339 14693 33373
rect 14647 33301 14693 33339
rect 14647 33267 14653 33301
rect 14687 33267 14693 33301
rect 14647 33229 14693 33267
rect 14647 33195 14653 33229
rect 14687 33195 14693 33229
rect 14647 33157 14693 33195
rect 14647 33123 14653 33157
rect 14687 33123 14693 33157
rect 14647 33085 14693 33123
rect 14647 33051 14653 33085
rect 14687 33051 14693 33085
rect 14647 33013 14693 33051
rect 14647 32979 14653 33013
rect 14687 32979 14693 33013
rect 14647 32941 14693 32979
rect 14647 32907 14653 32941
rect 14687 32907 14693 32941
rect 14647 32869 14693 32907
rect 14647 32835 14653 32869
rect 14687 32835 14693 32869
rect 14647 32797 14693 32835
rect 14647 32763 14653 32797
rect 14687 32763 14693 32797
rect 14647 32725 14693 32763
rect 14647 32691 14653 32725
rect 14687 32691 14693 32725
rect 14647 32653 14693 32691
rect 14647 32619 14653 32653
rect 14687 32619 14693 32653
rect 14647 32581 14693 32619
rect 14647 32547 14653 32581
rect 14687 32547 14693 32581
rect 14647 32509 14693 32547
rect 14647 32475 14653 32509
rect 14687 32475 14693 32509
rect 14647 32437 14693 32475
rect 14647 32403 14653 32437
rect 14687 32403 14693 32437
rect 14647 32387 14693 32403
rect 15105 33661 15151 33677
rect 15105 33627 15111 33661
rect 15145 33627 15151 33661
rect 15105 33589 15151 33627
rect 15105 33555 15111 33589
rect 15145 33555 15151 33589
rect 15105 33517 15151 33555
rect 15105 33483 15111 33517
rect 15145 33483 15151 33517
rect 15105 33445 15151 33483
rect 15105 33411 15111 33445
rect 15145 33411 15151 33445
rect 15105 33373 15151 33411
rect 15105 33339 15111 33373
rect 15145 33339 15151 33373
rect 15105 33301 15151 33339
rect 15105 33267 15111 33301
rect 15145 33267 15151 33301
rect 15105 33229 15151 33267
rect 15105 33195 15111 33229
rect 15145 33195 15151 33229
rect 15105 33157 15151 33195
rect 15105 33123 15111 33157
rect 15145 33123 15151 33157
rect 15105 33085 15151 33123
rect 15105 33051 15111 33085
rect 15145 33051 15151 33085
rect 15105 33013 15151 33051
rect 15105 32979 15111 33013
rect 15145 32979 15151 33013
rect 15105 32941 15151 32979
rect 15105 32907 15111 32941
rect 15145 32907 15151 32941
rect 15105 32869 15151 32907
rect 15105 32835 15111 32869
rect 15145 32835 15151 32869
rect 15105 32797 15151 32835
rect 15105 32763 15111 32797
rect 15145 32763 15151 32797
rect 15105 32725 15151 32763
rect 15105 32691 15111 32725
rect 15145 32691 15151 32725
rect 15105 32653 15151 32691
rect 15105 32619 15111 32653
rect 15145 32619 15151 32653
rect 15105 32581 15151 32619
rect 15105 32547 15111 32581
rect 15145 32547 15151 32581
rect 15105 32509 15151 32547
rect 15105 32475 15111 32509
rect 15145 32475 15151 32509
rect 15105 32437 15151 32475
rect 15105 32403 15111 32437
rect 15145 32403 15151 32437
rect 15105 32387 15151 32403
rect 15563 33661 15609 33677
rect 15563 33627 15569 33661
rect 15603 33627 15609 33661
rect 15563 33589 15609 33627
rect 15563 33555 15569 33589
rect 15603 33555 15609 33589
rect 15563 33517 15609 33555
rect 15563 33483 15569 33517
rect 15603 33483 15609 33517
rect 15563 33445 15609 33483
rect 15563 33411 15569 33445
rect 15603 33411 15609 33445
rect 15563 33373 15609 33411
rect 15563 33339 15569 33373
rect 15603 33339 15609 33373
rect 15563 33301 15609 33339
rect 15563 33267 15569 33301
rect 15603 33267 15609 33301
rect 15563 33229 15609 33267
rect 15563 33195 15569 33229
rect 15603 33195 15609 33229
rect 15563 33157 15609 33195
rect 15563 33123 15569 33157
rect 15603 33123 15609 33157
rect 15563 33085 15609 33123
rect 15563 33051 15569 33085
rect 15603 33051 15609 33085
rect 15563 33013 15609 33051
rect 15563 32979 15569 33013
rect 15603 32979 15609 33013
rect 15563 32941 15609 32979
rect 15563 32907 15569 32941
rect 15603 32907 15609 32941
rect 15563 32869 15609 32907
rect 15563 32835 15569 32869
rect 15603 32835 15609 32869
rect 15563 32797 15609 32835
rect 15563 32763 15569 32797
rect 15603 32763 15609 32797
rect 15563 32725 15609 32763
rect 15563 32691 15569 32725
rect 15603 32691 15609 32725
rect 15563 32653 15609 32691
rect 15563 32619 15569 32653
rect 15603 32619 15609 32653
rect 15563 32581 15609 32619
rect 15563 32547 15569 32581
rect 15603 32547 15609 32581
rect 15563 32509 15609 32547
rect 15563 32475 15569 32509
rect 15603 32475 15609 32509
rect 15563 32437 15609 32475
rect 15563 32403 15569 32437
rect 15603 32403 15609 32437
rect 15563 32387 15609 32403
rect 16021 33661 16067 33677
rect 16021 33627 16027 33661
rect 16061 33627 16067 33661
rect 16021 33589 16067 33627
rect 16021 33555 16027 33589
rect 16061 33555 16067 33589
rect 16021 33517 16067 33555
rect 16021 33483 16027 33517
rect 16061 33483 16067 33517
rect 16021 33445 16067 33483
rect 16021 33411 16027 33445
rect 16061 33411 16067 33445
rect 16021 33373 16067 33411
rect 16021 33339 16027 33373
rect 16061 33339 16067 33373
rect 16021 33301 16067 33339
rect 16021 33267 16027 33301
rect 16061 33267 16067 33301
rect 16021 33229 16067 33267
rect 16021 33195 16027 33229
rect 16061 33195 16067 33229
rect 16021 33157 16067 33195
rect 16021 33123 16027 33157
rect 16061 33123 16067 33157
rect 16021 33085 16067 33123
rect 16021 33051 16027 33085
rect 16061 33051 16067 33085
rect 16021 33013 16067 33051
rect 16021 32979 16027 33013
rect 16061 32979 16067 33013
rect 16021 32941 16067 32979
rect 16021 32907 16027 32941
rect 16061 32907 16067 32941
rect 16021 32869 16067 32907
rect 16021 32835 16027 32869
rect 16061 32835 16067 32869
rect 16021 32797 16067 32835
rect 16021 32763 16027 32797
rect 16061 32763 16067 32797
rect 16021 32725 16067 32763
rect 16021 32691 16027 32725
rect 16061 32691 16067 32725
rect 16021 32653 16067 32691
rect 16021 32619 16027 32653
rect 16061 32619 16067 32653
rect 16021 32581 16067 32619
rect 16021 32547 16027 32581
rect 16061 32547 16067 32581
rect 16021 32509 16067 32547
rect 16021 32475 16027 32509
rect 16061 32475 16067 32509
rect 16021 32437 16067 32475
rect 16021 32403 16027 32437
rect 16061 32403 16067 32437
rect 16021 32387 16067 32403
rect 16479 33661 16525 33677
rect 16479 33627 16485 33661
rect 16519 33627 16525 33661
rect 16479 33589 16525 33627
rect 16479 33555 16485 33589
rect 16519 33555 16525 33589
rect 16479 33517 16525 33555
rect 16479 33483 16485 33517
rect 16519 33483 16525 33517
rect 16479 33445 16525 33483
rect 16479 33411 16485 33445
rect 16519 33411 16525 33445
rect 16479 33373 16525 33411
rect 16479 33339 16485 33373
rect 16519 33339 16525 33373
rect 16479 33301 16525 33339
rect 16479 33267 16485 33301
rect 16519 33267 16525 33301
rect 16479 33229 16525 33267
rect 16479 33195 16485 33229
rect 16519 33195 16525 33229
rect 16479 33157 16525 33195
rect 16479 33123 16485 33157
rect 16519 33123 16525 33157
rect 16479 33085 16525 33123
rect 16479 33051 16485 33085
rect 16519 33051 16525 33085
rect 16479 33013 16525 33051
rect 16479 32979 16485 33013
rect 16519 32979 16525 33013
rect 16479 32941 16525 32979
rect 16479 32907 16485 32941
rect 16519 32907 16525 32941
rect 16479 32869 16525 32907
rect 16479 32835 16485 32869
rect 16519 32835 16525 32869
rect 16479 32797 16525 32835
rect 16479 32763 16485 32797
rect 16519 32763 16525 32797
rect 16479 32725 16525 32763
rect 16479 32691 16485 32725
rect 16519 32691 16525 32725
rect 16479 32653 16525 32691
rect 16479 32619 16485 32653
rect 16519 32619 16525 32653
rect 16479 32581 16525 32619
rect 16479 32547 16485 32581
rect 16519 32547 16525 32581
rect 16479 32509 16525 32547
rect 16479 32475 16485 32509
rect 16519 32475 16525 32509
rect 16479 32437 16525 32475
rect 16479 32403 16485 32437
rect 16519 32403 16525 32437
rect 16479 32387 16525 32403
rect 16937 33661 16983 33677
rect 16937 33627 16943 33661
rect 16977 33627 16983 33661
rect 16937 33589 16983 33627
rect 16937 33555 16943 33589
rect 16977 33555 16983 33589
rect 16937 33517 16983 33555
rect 16937 33483 16943 33517
rect 16977 33483 16983 33517
rect 16937 33445 16983 33483
rect 16937 33411 16943 33445
rect 16977 33411 16983 33445
rect 16937 33373 16983 33411
rect 16937 33339 16943 33373
rect 16977 33339 16983 33373
rect 16937 33301 16983 33339
rect 16937 33267 16943 33301
rect 16977 33267 16983 33301
rect 16937 33229 16983 33267
rect 16937 33195 16943 33229
rect 16977 33195 16983 33229
rect 16937 33157 16983 33195
rect 16937 33123 16943 33157
rect 16977 33123 16983 33157
rect 16937 33085 16983 33123
rect 16937 33051 16943 33085
rect 16977 33051 16983 33085
rect 16937 33013 16983 33051
rect 16937 32979 16943 33013
rect 16977 32979 16983 33013
rect 16937 32941 16983 32979
rect 16937 32907 16943 32941
rect 16977 32907 16983 32941
rect 16937 32869 16983 32907
rect 16937 32835 16943 32869
rect 16977 32835 16983 32869
rect 16937 32797 16983 32835
rect 16937 32763 16943 32797
rect 16977 32763 16983 32797
rect 16937 32725 16983 32763
rect 16937 32691 16943 32725
rect 16977 32691 16983 32725
rect 16937 32653 16983 32691
rect 16937 32619 16943 32653
rect 16977 32619 16983 32653
rect 16937 32581 16983 32619
rect 16937 32547 16943 32581
rect 16977 32547 16983 32581
rect 16937 32509 16983 32547
rect 16937 32475 16943 32509
rect 16977 32475 16983 32509
rect 16937 32437 16983 32475
rect 16937 32403 16943 32437
rect 16977 32403 16983 32437
rect 16937 32387 16983 32403
rect 17395 33661 17441 33677
rect 17395 33627 17401 33661
rect 17435 33627 17441 33661
rect 17395 33589 17441 33627
rect 17395 33555 17401 33589
rect 17435 33555 17441 33589
rect 17395 33517 17441 33555
rect 17395 33483 17401 33517
rect 17435 33483 17441 33517
rect 17395 33445 17441 33483
rect 17395 33411 17401 33445
rect 17435 33411 17441 33445
rect 17395 33373 17441 33411
rect 17395 33339 17401 33373
rect 17435 33339 17441 33373
rect 17395 33301 17441 33339
rect 17395 33267 17401 33301
rect 17435 33267 17441 33301
rect 17395 33229 17441 33267
rect 17395 33195 17401 33229
rect 17435 33195 17441 33229
rect 17395 33157 17441 33195
rect 17395 33123 17401 33157
rect 17435 33123 17441 33157
rect 17395 33085 17441 33123
rect 17395 33051 17401 33085
rect 17435 33051 17441 33085
rect 17395 33013 17441 33051
rect 17395 32979 17401 33013
rect 17435 32979 17441 33013
rect 17395 32941 17441 32979
rect 17395 32907 17401 32941
rect 17435 32907 17441 32941
rect 17395 32869 17441 32907
rect 17395 32835 17401 32869
rect 17435 32835 17441 32869
rect 17395 32797 17441 32835
rect 17395 32763 17401 32797
rect 17435 32763 17441 32797
rect 17395 32725 17441 32763
rect 17395 32691 17401 32725
rect 17435 32691 17441 32725
rect 17395 32653 17441 32691
rect 17395 32619 17401 32653
rect 17435 32619 17441 32653
rect 17395 32581 17441 32619
rect 17395 32547 17401 32581
rect 17435 32547 17441 32581
rect 17395 32509 17441 32547
rect 17395 32475 17401 32509
rect 17435 32475 17441 32509
rect 17395 32437 17441 32475
rect 17395 32403 17401 32437
rect 17435 32403 17441 32437
rect 17395 32387 17441 32403
rect 17853 33661 17899 33677
rect 17853 33627 17859 33661
rect 17893 33627 17899 33661
rect 17853 33589 17899 33627
rect 17853 33555 17859 33589
rect 17893 33555 17899 33589
rect 17853 33517 17899 33555
rect 17853 33483 17859 33517
rect 17893 33483 17899 33517
rect 17853 33445 17899 33483
rect 17853 33411 17859 33445
rect 17893 33411 17899 33445
rect 17853 33373 17899 33411
rect 17853 33339 17859 33373
rect 17893 33339 17899 33373
rect 17853 33301 17899 33339
rect 17853 33267 17859 33301
rect 17893 33267 17899 33301
rect 17853 33229 17899 33267
rect 17853 33195 17859 33229
rect 17893 33195 17899 33229
rect 17853 33157 17899 33195
rect 17853 33123 17859 33157
rect 17893 33123 17899 33157
rect 17853 33085 17899 33123
rect 17853 33051 17859 33085
rect 17893 33051 17899 33085
rect 17853 33013 17899 33051
rect 17853 32979 17859 33013
rect 17893 32979 17899 33013
rect 17853 32941 17899 32979
rect 17853 32907 17859 32941
rect 17893 32907 17899 32941
rect 17853 32869 17899 32907
rect 17853 32835 17859 32869
rect 17893 32835 17899 32869
rect 17853 32797 17899 32835
rect 17853 32763 17859 32797
rect 17893 32763 17899 32797
rect 17853 32725 17899 32763
rect 17853 32691 17859 32725
rect 17893 32691 17899 32725
rect 17853 32653 17899 32691
rect 17853 32619 17859 32653
rect 17893 32619 17899 32653
rect 17853 32581 17899 32619
rect 17853 32547 17859 32581
rect 17893 32547 17899 32581
rect 17853 32509 17899 32547
rect 17853 32475 17859 32509
rect 17893 32475 17899 32509
rect 17853 32437 17899 32475
rect 17853 32403 17859 32437
rect 17893 32403 17899 32437
rect 17853 32387 17899 32403
rect 18311 33661 18357 33677
rect 18311 33627 18317 33661
rect 18351 33627 18357 33661
rect 18311 33589 18357 33627
rect 18311 33555 18317 33589
rect 18351 33555 18357 33589
rect 18311 33517 18357 33555
rect 18311 33483 18317 33517
rect 18351 33483 18357 33517
rect 18311 33445 18357 33483
rect 18311 33411 18317 33445
rect 18351 33411 18357 33445
rect 18311 33373 18357 33411
rect 18311 33339 18317 33373
rect 18351 33339 18357 33373
rect 18311 33301 18357 33339
rect 18311 33267 18317 33301
rect 18351 33267 18357 33301
rect 18311 33229 18357 33267
rect 18311 33195 18317 33229
rect 18351 33195 18357 33229
rect 18311 33157 18357 33195
rect 18311 33123 18317 33157
rect 18351 33123 18357 33157
rect 18311 33085 18357 33123
rect 18311 33051 18317 33085
rect 18351 33051 18357 33085
rect 18311 33013 18357 33051
rect 18311 32979 18317 33013
rect 18351 32979 18357 33013
rect 18311 32941 18357 32979
rect 18311 32907 18317 32941
rect 18351 32907 18357 32941
rect 18311 32869 18357 32907
rect 18311 32835 18317 32869
rect 18351 32835 18357 32869
rect 18311 32797 18357 32835
rect 18311 32763 18317 32797
rect 18351 32763 18357 32797
rect 18311 32725 18357 32763
rect 18311 32691 18317 32725
rect 18351 32691 18357 32725
rect 18311 32653 18357 32691
rect 18311 32619 18317 32653
rect 18351 32619 18357 32653
rect 18311 32581 18357 32619
rect 18311 32547 18317 32581
rect 18351 32547 18357 32581
rect 18311 32509 18357 32547
rect 18311 32475 18317 32509
rect 18351 32475 18357 32509
rect 18311 32437 18357 32475
rect 18311 32403 18317 32437
rect 18351 32403 18357 32437
rect 18311 32387 18357 32403
rect 18769 33661 18815 33677
rect 18769 33627 18775 33661
rect 18809 33627 18815 33661
rect 18769 33589 18815 33627
rect 18769 33555 18775 33589
rect 18809 33555 18815 33589
rect 18769 33517 18815 33555
rect 18769 33483 18775 33517
rect 18809 33483 18815 33517
rect 18769 33445 18815 33483
rect 18769 33411 18775 33445
rect 18809 33411 18815 33445
rect 18769 33373 18815 33411
rect 18769 33339 18775 33373
rect 18809 33339 18815 33373
rect 18769 33301 18815 33339
rect 18769 33267 18775 33301
rect 18809 33267 18815 33301
rect 18769 33229 18815 33267
rect 18769 33195 18775 33229
rect 18809 33195 18815 33229
rect 18769 33157 18815 33195
rect 18769 33123 18775 33157
rect 18809 33123 18815 33157
rect 18769 33085 18815 33123
rect 18769 33051 18775 33085
rect 18809 33051 18815 33085
rect 18769 33013 18815 33051
rect 18769 32979 18775 33013
rect 18809 32979 18815 33013
rect 18769 32941 18815 32979
rect 18769 32907 18775 32941
rect 18809 32907 18815 32941
rect 18769 32869 18815 32907
rect 18769 32835 18775 32869
rect 18809 32835 18815 32869
rect 18769 32797 18815 32835
rect 18769 32763 18775 32797
rect 18809 32763 18815 32797
rect 18769 32725 18815 32763
rect 18769 32691 18775 32725
rect 18809 32691 18815 32725
rect 18769 32653 18815 32691
rect 18769 32619 18775 32653
rect 18809 32619 18815 32653
rect 18769 32581 18815 32619
rect 18769 32547 18775 32581
rect 18809 32547 18815 32581
rect 18769 32509 18815 32547
rect 18769 32475 18775 32509
rect 18809 32475 18815 32509
rect 18769 32437 18815 32475
rect 18769 32403 18775 32437
rect 18809 32403 18815 32437
rect 18769 32387 18815 32403
rect 19227 33661 19273 33677
rect 19227 33627 19233 33661
rect 19267 33627 19273 33661
rect 19227 33589 19273 33627
rect 19227 33555 19233 33589
rect 19267 33555 19273 33589
rect 19227 33517 19273 33555
rect 19227 33483 19233 33517
rect 19267 33483 19273 33517
rect 19227 33445 19273 33483
rect 19227 33411 19233 33445
rect 19267 33411 19273 33445
rect 19227 33373 19273 33411
rect 19227 33339 19233 33373
rect 19267 33339 19273 33373
rect 19227 33301 19273 33339
rect 19227 33267 19233 33301
rect 19267 33267 19273 33301
rect 19227 33229 19273 33267
rect 19227 33195 19233 33229
rect 19267 33195 19273 33229
rect 19227 33157 19273 33195
rect 19227 33123 19233 33157
rect 19267 33123 19273 33157
rect 19227 33085 19273 33123
rect 19227 33051 19233 33085
rect 19267 33051 19273 33085
rect 19227 33013 19273 33051
rect 19227 32979 19233 33013
rect 19267 32979 19273 33013
rect 19227 32941 19273 32979
rect 19227 32907 19233 32941
rect 19267 32907 19273 32941
rect 19227 32869 19273 32907
rect 19227 32835 19233 32869
rect 19267 32835 19273 32869
rect 19227 32797 19273 32835
rect 19227 32763 19233 32797
rect 19267 32763 19273 32797
rect 19227 32725 19273 32763
rect 19227 32691 19233 32725
rect 19267 32691 19273 32725
rect 19227 32653 19273 32691
rect 19227 32619 19233 32653
rect 19267 32619 19273 32653
rect 19227 32581 19273 32619
rect 19227 32547 19233 32581
rect 19267 32547 19273 32581
rect 19227 32509 19273 32547
rect 19227 32475 19233 32509
rect 19267 32475 19273 32509
rect 19227 32437 19273 32475
rect 19227 32403 19233 32437
rect 19267 32403 19273 32437
rect 19227 32387 19273 32403
rect 19685 33661 19731 33677
rect 19685 33627 19691 33661
rect 19725 33627 19731 33661
rect 19685 33589 19731 33627
rect 19685 33555 19691 33589
rect 19725 33555 19731 33589
rect 19685 33517 19731 33555
rect 19685 33483 19691 33517
rect 19725 33483 19731 33517
rect 19685 33445 19731 33483
rect 19685 33411 19691 33445
rect 19725 33411 19731 33445
rect 19685 33373 19731 33411
rect 19685 33339 19691 33373
rect 19725 33339 19731 33373
rect 19685 33301 19731 33339
rect 19685 33267 19691 33301
rect 19725 33267 19731 33301
rect 19685 33229 19731 33267
rect 19685 33195 19691 33229
rect 19725 33195 19731 33229
rect 19685 33157 19731 33195
rect 19685 33123 19691 33157
rect 19725 33123 19731 33157
rect 19685 33085 19731 33123
rect 19685 33051 19691 33085
rect 19725 33051 19731 33085
rect 19685 33013 19731 33051
rect 19685 32979 19691 33013
rect 19725 32979 19731 33013
rect 19685 32941 19731 32979
rect 19685 32907 19691 32941
rect 19725 32907 19731 32941
rect 19685 32869 19731 32907
rect 19685 32835 19691 32869
rect 19725 32835 19731 32869
rect 19685 32797 19731 32835
rect 19685 32763 19691 32797
rect 19725 32763 19731 32797
rect 19685 32725 19731 32763
rect 19685 32691 19691 32725
rect 19725 32691 19731 32725
rect 19685 32653 19731 32691
rect 19685 32619 19691 32653
rect 19725 32619 19731 32653
rect 19685 32581 19731 32619
rect 19685 32547 19691 32581
rect 19725 32547 19731 32581
rect 19685 32509 19731 32547
rect 19685 32475 19691 32509
rect 19725 32475 19731 32509
rect 19685 32437 19731 32475
rect 19685 32403 19691 32437
rect 19725 32403 19731 32437
rect 19685 32387 19731 32403
rect 20143 33661 20189 33677
rect 20143 33627 20149 33661
rect 20183 33627 20189 33661
rect 20143 33589 20189 33627
rect 20143 33555 20149 33589
rect 20183 33555 20189 33589
rect 20143 33517 20189 33555
rect 20143 33483 20149 33517
rect 20183 33483 20189 33517
rect 20143 33445 20189 33483
rect 20143 33411 20149 33445
rect 20183 33411 20189 33445
rect 20143 33373 20189 33411
rect 20143 33339 20149 33373
rect 20183 33339 20189 33373
rect 20143 33301 20189 33339
rect 20143 33267 20149 33301
rect 20183 33267 20189 33301
rect 20143 33229 20189 33267
rect 20143 33195 20149 33229
rect 20183 33195 20189 33229
rect 20143 33157 20189 33195
rect 20143 33123 20149 33157
rect 20183 33123 20189 33157
rect 20143 33085 20189 33123
rect 20143 33051 20149 33085
rect 20183 33051 20189 33085
rect 20143 33013 20189 33051
rect 20143 32979 20149 33013
rect 20183 32979 20189 33013
rect 20143 32941 20189 32979
rect 20143 32907 20149 32941
rect 20183 32907 20189 32941
rect 20143 32869 20189 32907
rect 20143 32835 20149 32869
rect 20183 32835 20189 32869
rect 20143 32797 20189 32835
rect 20143 32763 20149 32797
rect 20183 32763 20189 32797
rect 20143 32725 20189 32763
rect 20143 32691 20149 32725
rect 20183 32691 20189 32725
rect 20143 32653 20189 32691
rect 20143 32619 20149 32653
rect 20183 32619 20189 32653
rect 20143 32581 20189 32619
rect 20143 32547 20149 32581
rect 20183 32547 20189 32581
rect 20143 32509 20189 32547
rect 20143 32475 20149 32509
rect 20183 32475 20189 32509
rect 20143 32437 20189 32475
rect 20143 32403 20149 32437
rect 20183 32403 20189 32437
rect 20143 32387 20189 32403
rect 20601 33661 20647 33677
rect 20601 33627 20607 33661
rect 20641 33627 20647 33661
rect 20601 33589 20647 33627
rect 20601 33555 20607 33589
rect 20641 33555 20647 33589
rect 20601 33517 20647 33555
rect 20601 33483 20607 33517
rect 20641 33483 20647 33517
rect 20601 33445 20647 33483
rect 20601 33411 20607 33445
rect 20641 33411 20647 33445
rect 20601 33373 20647 33411
rect 20601 33339 20607 33373
rect 20641 33339 20647 33373
rect 20601 33301 20647 33339
rect 20601 33267 20607 33301
rect 20641 33267 20647 33301
rect 20601 33229 20647 33267
rect 20601 33195 20607 33229
rect 20641 33195 20647 33229
rect 20601 33157 20647 33195
rect 20601 33123 20607 33157
rect 20641 33123 20647 33157
rect 20601 33085 20647 33123
rect 20601 33051 20607 33085
rect 20641 33051 20647 33085
rect 20601 33013 20647 33051
rect 20601 32979 20607 33013
rect 20641 32979 20647 33013
rect 20601 32941 20647 32979
rect 20601 32907 20607 32941
rect 20641 32907 20647 32941
rect 20601 32869 20647 32907
rect 20601 32835 20607 32869
rect 20641 32835 20647 32869
rect 20601 32797 20647 32835
rect 20601 32763 20607 32797
rect 20641 32763 20647 32797
rect 20601 32725 20647 32763
rect 20601 32691 20607 32725
rect 20641 32691 20647 32725
rect 20601 32653 20647 32691
rect 20601 32619 20607 32653
rect 20641 32619 20647 32653
rect 20601 32581 20647 32619
rect 20601 32547 20607 32581
rect 20641 32547 20647 32581
rect 20601 32509 20647 32547
rect 20601 32475 20607 32509
rect 20641 32475 20647 32509
rect 20601 32437 20647 32475
rect 20601 32403 20607 32437
rect 20641 32403 20647 32437
rect 20601 32387 20647 32403
rect 21059 33661 21105 33677
rect 21059 33627 21065 33661
rect 21099 33627 21105 33661
rect 21059 33589 21105 33627
rect 21059 33555 21065 33589
rect 21099 33555 21105 33589
rect 21059 33517 21105 33555
rect 21059 33483 21065 33517
rect 21099 33483 21105 33517
rect 21059 33445 21105 33483
rect 21059 33411 21065 33445
rect 21099 33411 21105 33445
rect 21059 33373 21105 33411
rect 21059 33339 21065 33373
rect 21099 33339 21105 33373
rect 21059 33301 21105 33339
rect 21059 33267 21065 33301
rect 21099 33267 21105 33301
rect 21059 33229 21105 33267
rect 21059 33195 21065 33229
rect 21099 33195 21105 33229
rect 21059 33157 21105 33195
rect 21059 33123 21065 33157
rect 21099 33123 21105 33157
rect 21059 33085 21105 33123
rect 21059 33051 21065 33085
rect 21099 33051 21105 33085
rect 21059 33013 21105 33051
rect 21059 32979 21065 33013
rect 21099 32979 21105 33013
rect 21059 32941 21105 32979
rect 21059 32907 21065 32941
rect 21099 32907 21105 32941
rect 21059 32869 21105 32907
rect 21059 32835 21065 32869
rect 21099 32835 21105 32869
rect 21059 32797 21105 32835
rect 21059 32763 21065 32797
rect 21099 32763 21105 32797
rect 21059 32725 21105 32763
rect 21059 32691 21065 32725
rect 21099 32691 21105 32725
rect 21059 32653 21105 32691
rect 21059 32619 21065 32653
rect 21099 32619 21105 32653
rect 21059 32581 21105 32619
rect 21059 32547 21065 32581
rect 21099 32547 21105 32581
rect 21059 32509 21105 32547
rect 21059 32475 21065 32509
rect 21099 32475 21105 32509
rect 21059 32437 21105 32475
rect 21059 32403 21065 32437
rect 21099 32403 21105 32437
rect 21059 32387 21105 32403
rect 21517 33661 21563 33677
rect 21517 33627 21523 33661
rect 21557 33627 21563 33661
rect 21517 33589 21563 33627
rect 21517 33555 21523 33589
rect 21557 33555 21563 33589
rect 21517 33517 21563 33555
rect 21517 33483 21523 33517
rect 21557 33483 21563 33517
rect 21517 33445 21563 33483
rect 21517 33411 21523 33445
rect 21557 33411 21563 33445
rect 21517 33373 21563 33411
rect 21517 33339 21523 33373
rect 21557 33339 21563 33373
rect 21517 33301 21563 33339
rect 21517 33267 21523 33301
rect 21557 33267 21563 33301
rect 21517 33229 21563 33267
rect 21517 33195 21523 33229
rect 21557 33195 21563 33229
rect 21517 33157 21563 33195
rect 21517 33123 21523 33157
rect 21557 33123 21563 33157
rect 21517 33085 21563 33123
rect 21517 33051 21523 33085
rect 21557 33051 21563 33085
rect 21517 33013 21563 33051
rect 21517 32979 21523 33013
rect 21557 32979 21563 33013
rect 21517 32941 21563 32979
rect 21517 32907 21523 32941
rect 21557 32907 21563 32941
rect 21517 32869 21563 32907
rect 21517 32835 21523 32869
rect 21557 32835 21563 32869
rect 21517 32797 21563 32835
rect 21517 32763 21523 32797
rect 21557 32763 21563 32797
rect 21517 32725 21563 32763
rect 21517 32691 21523 32725
rect 21557 32691 21563 32725
rect 21517 32653 21563 32691
rect 21517 32619 21523 32653
rect 21557 32619 21563 32653
rect 21517 32581 21563 32619
rect 21517 32547 21523 32581
rect 21557 32547 21563 32581
rect 21517 32509 21563 32547
rect 21517 32475 21523 32509
rect 21557 32475 21563 32509
rect 21517 32437 21563 32475
rect 21517 32403 21523 32437
rect 21557 32403 21563 32437
rect 21517 32387 21563 32403
rect 21975 33661 22021 33677
rect 21975 33627 21981 33661
rect 22015 33627 22021 33661
rect 21975 33589 22021 33627
rect 21975 33555 21981 33589
rect 22015 33555 22021 33589
rect 21975 33517 22021 33555
rect 21975 33483 21981 33517
rect 22015 33483 22021 33517
rect 21975 33445 22021 33483
rect 21975 33411 21981 33445
rect 22015 33411 22021 33445
rect 21975 33373 22021 33411
rect 21975 33339 21981 33373
rect 22015 33339 22021 33373
rect 21975 33301 22021 33339
rect 21975 33267 21981 33301
rect 22015 33267 22021 33301
rect 21975 33229 22021 33267
rect 21975 33195 21981 33229
rect 22015 33195 22021 33229
rect 21975 33157 22021 33195
rect 21975 33123 21981 33157
rect 22015 33123 22021 33157
rect 21975 33085 22021 33123
rect 21975 33051 21981 33085
rect 22015 33051 22021 33085
rect 21975 33013 22021 33051
rect 21975 32979 21981 33013
rect 22015 32979 22021 33013
rect 21975 32941 22021 32979
rect 21975 32907 21981 32941
rect 22015 32907 22021 32941
rect 21975 32869 22021 32907
rect 21975 32835 21981 32869
rect 22015 32835 22021 32869
rect 21975 32797 22021 32835
rect 21975 32763 21981 32797
rect 22015 32763 22021 32797
rect 21975 32725 22021 32763
rect 21975 32691 21981 32725
rect 22015 32691 22021 32725
rect 21975 32653 22021 32691
rect 21975 32619 21981 32653
rect 22015 32619 22021 32653
rect 21975 32581 22021 32619
rect 21975 32547 21981 32581
rect 22015 32547 22021 32581
rect 21975 32509 22021 32547
rect 21975 32475 21981 32509
rect 22015 32475 22021 32509
rect 21975 32437 22021 32475
rect 21975 32403 21981 32437
rect 22015 32403 22021 32437
rect 21975 32387 22021 32403
rect 22433 33661 22479 33677
rect 22433 33627 22439 33661
rect 22473 33627 22479 33661
rect 22433 33589 22479 33627
rect 22433 33555 22439 33589
rect 22473 33555 22479 33589
rect 22433 33517 22479 33555
rect 22433 33483 22439 33517
rect 22473 33483 22479 33517
rect 22433 33445 22479 33483
rect 22433 33411 22439 33445
rect 22473 33411 22479 33445
rect 22433 33373 22479 33411
rect 22433 33339 22439 33373
rect 22473 33339 22479 33373
rect 22433 33301 22479 33339
rect 22433 33267 22439 33301
rect 22473 33267 22479 33301
rect 22433 33229 22479 33267
rect 22433 33195 22439 33229
rect 22473 33195 22479 33229
rect 22433 33157 22479 33195
rect 22433 33123 22439 33157
rect 22473 33123 22479 33157
rect 22433 33085 22479 33123
rect 22433 33051 22439 33085
rect 22473 33051 22479 33085
rect 22433 33013 22479 33051
rect 22433 32979 22439 33013
rect 22473 32979 22479 33013
rect 22433 32941 22479 32979
rect 22433 32907 22439 32941
rect 22473 32907 22479 32941
rect 22433 32869 22479 32907
rect 22433 32835 22439 32869
rect 22473 32835 22479 32869
rect 22433 32797 22479 32835
rect 22433 32763 22439 32797
rect 22473 32763 22479 32797
rect 22433 32725 22479 32763
rect 22433 32691 22439 32725
rect 22473 32691 22479 32725
rect 22433 32653 22479 32691
rect 22433 32619 22439 32653
rect 22473 32619 22479 32653
rect 22433 32581 22479 32619
rect 22433 32547 22439 32581
rect 22473 32547 22479 32581
rect 22433 32509 22479 32547
rect 22433 32475 22439 32509
rect 22473 32475 22479 32509
rect 22433 32437 22479 32475
rect 22433 32403 22439 32437
rect 22473 32403 22479 32437
rect 22433 32387 22479 32403
rect 22891 33661 22937 33677
rect 22891 33627 22897 33661
rect 22931 33627 22937 33661
rect 22891 33589 22937 33627
rect 22891 33555 22897 33589
rect 22931 33555 22937 33589
rect 22891 33517 22937 33555
rect 22891 33483 22897 33517
rect 22931 33483 22937 33517
rect 22891 33445 22937 33483
rect 22891 33411 22897 33445
rect 22931 33411 22937 33445
rect 22891 33373 22937 33411
rect 22891 33339 22897 33373
rect 22931 33339 22937 33373
rect 22891 33301 22937 33339
rect 22891 33267 22897 33301
rect 22931 33267 22937 33301
rect 22891 33229 22937 33267
rect 22891 33195 22897 33229
rect 22931 33195 22937 33229
rect 22891 33157 22937 33195
rect 22891 33123 22897 33157
rect 22931 33123 22937 33157
rect 22891 33085 22937 33123
rect 22891 33051 22897 33085
rect 22931 33051 22937 33085
rect 22891 33013 22937 33051
rect 22891 32979 22897 33013
rect 22931 32979 22937 33013
rect 22891 32941 22937 32979
rect 22891 32907 22897 32941
rect 22931 32907 22937 32941
rect 22891 32869 22937 32907
rect 22891 32835 22897 32869
rect 22931 32835 22937 32869
rect 22891 32797 22937 32835
rect 22891 32763 22897 32797
rect 22931 32763 22937 32797
rect 22891 32725 22937 32763
rect 22891 32691 22897 32725
rect 22931 32691 22937 32725
rect 22891 32653 22937 32691
rect 22891 32619 22897 32653
rect 22931 32619 22937 32653
rect 22891 32581 22937 32619
rect 22891 32547 22897 32581
rect 22931 32547 22937 32581
rect 22891 32509 22937 32547
rect 22891 32475 22897 32509
rect 22931 32475 22937 32509
rect 22891 32437 22937 32475
rect 22891 32403 22897 32437
rect 22931 32403 22937 32437
rect 22891 32387 22937 32403
rect 23349 33661 23395 33677
rect 23349 33627 23355 33661
rect 23389 33627 23395 33661
rect 23349 33589 23395 33627
rect 23349 33555 23355 33589
rect 23389 33555 23395 33589
rect 23349 33517 23395 33555
rect 23349 33483 23355 33517
rect 23389 33483 23395 33517
rect 23349 33445 23395 33483
rect 23349 33411 23355 33445
rect 23389 33411 23395 33445
rect 23349 33373 23395 33411
rect 23349 33339 23355 33373
rect 23389 33339 23395 33373
rect 23349 33301 23395 33339
rect 23349 33267 23355 33301
rect 23389 33267 23395 33301
rect 23349 33229 23395 33267
rect 23349 33195 23355 33229
rect 23389 33195 23395 33229
rect 23349 33157 23395 33195
rect 23349 33123 23355 33157
rect 23389 33123 23395 33157
rect 23349 33085 23395 33123
rect 23349 33051 23355 33085
rect 23389 33051 23395 33085
rect 23349 33013 23395 33051
rect 23349 32979 23355 33013
rect 23389 32979 23395 33013
rect 23349 32941 23395 32979
rect 23349 32907 23355 32941
rect 23389 32907 23395 32941
rect 23349 32869 23395 32907
rect 23349 32835 23355 32869
rect 23389 32835 23395 32869
rect 23349 32797 23395 32835
rect 23349 32763 23355 32797
rect 23389 32763 23395 32797
rect 23349 32725 23395 32763
rect 23349 32691 23355 32725
rect 23389 32691 23395 32725
rect 23349 32653 23395 32691
rect 23349 32619 23355 32653
rect 23389 32619 23395 32653
rect 23349 32581 23395 32619
rect 23349 32547 23355 32581
rect 23389 32547 23395 32581
rect 23349 32509 23395 32547
rect 23349 32475 23355 32509
rect 23389 32475 23395 32509
rect 23349 32437 23395 32475
rect 23349 32403 23355 32437
rect 23389 32403 23395 32437
rect 23349 32387 23395 32403
rect 23807 33661 23853 33677
rect 23807 33627 23813 33661
rect 23847 33627 23853 33661
rect 23807 33589 23853 33627
rect 23807 33555 23813 33589
rect 23847 33555 23853 33589
rect 23807 33517 23853 33555
rect 23807 33483 23813 33517
rect 23847 33483 23853 33517
rect 23807 33445 23853 33483
rect 23807 33411 23813 33445
rect 23847 33411 23853 33445
rect 23807 33373 23853 33411
rect 23807 33339 23813 33373
rect 23847 33339 23853 33373
rect 23807 33301 23853 33339
rect 23807 33267 23813 33301
rect 23847 33267 23853 33301
rect 23807 33229 23853 33267
rect 23807 33195 23813 33229
rect 23847 33195 23853 33229
rect 23807 33157 23853 33195
rect 23807 33123 23813 33157
rect 23847 33123 23853 33157
rect 23807 33085 23853 33123
rect 23807 33051 23813 33085
rect 23847 33051 23853 33085
rect 23807 33013 23853 33051
rect 23807 32979 23813 33013
rect 23847 32979 23853 33013
rect 23807 32941 23853 32979
rect 23807 32907 23813 32941
rect 23847 32907 23853 32941
rect 23807 32869 23853 32907
rect 23807 32835 23813 32869
rect 23847 32835 23853 32869
rect 23807 32797 23853 32835
rect 23807 32763 23813 32797
rect 23847 32763 23853 32797
rect 23807 32725 23853 32763
rect 23807 32691 23813 32725
rect 23847 32691 23853 32725
rect 23807 32653 23853 32691
rect 23807 32619 23813 32653
rect 23847 32619 23853 32653
rect 23807 32581 23853 32619
rect 23807 32547 23813 32581
rect 23847 32547 23853 32581
rect 23807 32509 23853 32547
rect 23807 32475 23813 32509
rect 23847 32475 23853 32509
rect 23807 32437 23853 32475
rect 23807 32403 23813 32437
rect 23847 32403 23853 32437
rect 23807 32387 23853 32403
rect 24265 33661 24311 33677
rect 24265 33627 24271 33661
rect 24305 33627 24311 33661
rect 24265 33589 24311 33627
rect 24265 33555 24271 33589
rect 24305 33555 24311 33589
rect 24265 33517 24311 33555
rect 24265 33483 24271 33517
rect 24305 33483 24311 33517
rect 24265 33445 24311 33483
rect 24265 33411 24271 33445
rect 24305 33411 24311 33445
rect 24265 33373 24311 33411
rect 24265 33339 24271 33373
rect 24305 33339 24311 33373
rect 24265 33301 24311 33339
rect 24265 33267 24271 33301
rect 24305 33267 24311 33301
rect 24265 33229 24311 33267
rect 24265 33195 24271 33229
rect 24305 33195 24311 33229
rect 24265 33157 24311 33195
rect 24265 33123 24271 33157
rect 24305 33123 24311 33157
rect 24265 33085 24311 33123
rect 24265 33051 24271 33085
rect 24305 33051 24311 33085
rect 24265 33013 24311 33051
rect 24265 32979 24271 33013
rect 24305 32979 24311 33013
rect 24265 32941 24311 32979
rect 24265 32907 24271 32941
rect 24305 32907 24311 32941
rect 24265 32869 24311 32907
rect 24265 32835 24271 32869
rect 24305 32835 24311 32869
rect 24265 32797 24311 32835
rect 24265 32763 24271 32797
rect 24305 32763 24311 32797
rect 24265 32725 24311 32763
rect 24265 32691 24271 32725
rect 24305 32691 24311 32725
rect 24265 32653 24311 32691
rect 24265 32619 24271 32653
rect 24305 32619 24311 32653
rect 24265 32581 24311 32619
rect 24265 32547 24271 32581
rect 24305 32547 24311 32581
rect 24265 32509 24311 32547
rect 24265 32475 24271 32509
rect 24305 32475 24311 32509
rect 24265 32437 24311 32475
rect 24265 32403 24271 32437
rect 24305 32403 24311 32437
rect 24265 32387 24311 32403
rect 24723 33661 24769 33677
rect 24723 33627 24729 33661
rect 24763 33627 24769 33661
rect 24723 33589 24769 33627
rect 24723 33555 24729 33589
rect 24763 33555 24769 33589
rect 24723 33517 24769 33555
rect 24723 33483 24729 33517
rect 24763 33483 24769 33517
rect 24723 33445 24769 33483
rect 24723 33411 24729 33445
rect 24763 33411 24769 33445
rect 24723 33373 24769 33411
rect 24723 33339 24729 33373
rect 24763 33339 24769 33373
rect 24723 33301 24769 33339
rect 24723 33267 24729 33301
rect 24763 33267 24769 33301
rect 24723 33229 24769 33267
rect 24723 33195 24729 33229
rect 24763 33195 24769 33229
rect 24723 33157 24769 33195
rect 24723 33123 24729 33157
rect 24763 33123 24769 33157
rect 24723 33085 24769 33123
rect 24723 33051 24729 33085
rect 24763 33051 24769 33085
rect 24723 33013 24769 33051
rect 24723 32979 24729 33013
rect 24763 32979 24769 33013
rect 24723 32941 24769 32979
rect 24723 32907 24729 32941
rect 24763 32907 24769 32941
rect 24723 32869 24769 32907
rect 24723 32835 24729 32869
rect 24763 32835 24769 32869
rect 24723 32797 24769 32835
rect 24723 32763 24729 32797
rect 24763 32763 24769 32797
rect 24723 32725 24769 32763
rect 24723 32691 24729 32725
rect 24763 32691 24769 32725
rect 24723 32653 24769 32691
rect 24723 32619 24729 32653
rect 24763 32619 24769 32653
rect 24723 32581 24769 32619
rect 24723 32547 24729 32581
rect 24763 32547 24769 32581
rect 24723 32509 24769 32547
rect 24723 32475 24729 32509
rect 24763 32475 24769 32509
rect 24723 32437 24769 32475
rect 24723 32403 24729 32437
rect 24763 32403 24769 32437
rect 24723 32387 24769 32403
rect 25181 33661 25227 33677
rect 25181 33627 25187 33661
rect 25221 33627 25227 33661
rect 25181 33589 25227 33627
rect 25181 33555 25187 33589
rect 25221 33555 25227 33589
rect 25181 33517 25227 33555
rect 25181 33483 25187 33517
rect 25221 33483 25227 33517
rect 25181 33445 25227 33483
rect 25181 33411 25187 33445
rect 25221 33411 25227 33445
rect 25181 33373 25227 33411
rect 25181 33339 25187 33373
rect 25221 33339 25227 33373
rect 25181 33301 25227 33339
rect 25181 33267 25187 33301
rect 25221 33267 25227 33301
rect 25181 33229 25227 33267
rect 25181 33195 25187 33229
rect 25221 33195 25227 33229
rect 25181 33157 25227 33195
rect 25181 33123 25187 33157
rect 25221 33123 25227 33157
rect 25181 33085 25227 33123
rect 25181 33051 25187 33085
rect 25221 33051 25227 33085
rect 25181 33013 25227 33051
rect 25181 32979 25187 33013
rect 25221 32979 25227 33013
rect 25181 32941 25227 32979
rect 25181 32907 25187 32941
rect 25221 32907 25227 32941
rect 25181 32869 25227 32907
rect 25181 32835 25187 32869
rect 25221 32835 25227 32869
rect 25181 32797 25227 32835
rect 25181 32763 25187 32797
rect 25221 32763 25227 32797
rect 25181 32725 25227 32763
rect 25181 32691 25187 32725
rect 25221 32691 25227 32725
rect 25181 32653 25227 32691
rect 25181 32619 25187 32653
rect 25221 32619 25227 32653
rect 25181 32581 25227 32619
rect 25181 32547 25187 32581
rect 25221 32547 25227 32581
rect 25181 32509 25227 32547
rect 25181 32475 25187 32509
rect 25221 32475 25227 32509
rect 25181 32437 25227 32475
rect 25181 32403 25187 32437
rect 25221 32403 25227 32437
rect 25181 32387 25227 32403
rect 25639 33661 25685 33677
rect 25639 33627 25645 33661
rect 25679 33627 25685 33661
rect 25639 33589 25685 33627
rect 25639 33555 25645 33589
rect 25679 33555 25685 33589
rect 25639 33517 25685 33555
rect 25639 33483 25645 33517
rect 25679 33483 25685 33517
rect 25639 33445 25685 33483
rect 25639 33411 25645 33445
rect 25679 33411 25685 33445
rect 25639 33373 25685 33411
rect 25639 33339 25645 33373
rect 25679 33339 25685 33373
rect 25639 33301 25685 33339
rect 25639 33267 25645 33301
rect 25679 33267 25685 33301
rect 25639 33229 25685 33267
rect 25639 33195 25645 33229
rect 25679 33195 25685 33229
rect 25639 33157 25685 33195
rect 25639 33123 25645 33157
rect 25679 33123 25685 33157
rect 25639 33085 25685 33123
rect 25639 33051 25645 33085
rect 25679 33051 25685 33085
rect 25639 33013 25685 33051
rect 25639 32979 25645 33013
rect 25679 32979 25685 33013
rect 25639 32941 25685 32979
rect 25639 32907 25645 32941
rect 25679 32907 25685 32941
rect 25639 32869 25685 32907
rect 25639 32835 25645 32869
rect 25679 32835 25685 32869
rect 25639 32797 25685 32835
rect 25639 32763 25645 32797
rect 25679 32763 25685 32797
rect 25639 32725 25685 32763
rect 25639 32691 25645 32725
rect 25679 32691 25685 32725
rect 25639 32653 25685 32691
rect 25639 32619 25645 32653
rect 25679 32619 25685 32653
rect 25639 32581 25685 32619
rect 25639 32547 25645 32581
rect 25679 32547 25685 32581
rect 25639 32509 25685 32547
rect 25639 32475 25645 32509
rect 25679 32475 25685 32509
rect 25639 32437 25685 32475
rect 25639 32403 25645 32437
rect 25679 32403 25685 32437
rect 25639 32387 25685 32403
rect 26097 33661 26143 33677
rect 26097 33627 26103 33661
rect 26137 33627 26143 33661
rect 26097 33589 26143 33627
rect 26097 33555 26103 33589
rect 26137 33555 26143 33589
rect 26097 33517 26143 33555
rect 26097 33483 26103 33517
rect 26137 33483 26143 33517
rect 26097 33445 26143 33483
rect 26097 33411 26103 33445
rect 26137 33411 26143 33445
rect 26097 33373 26143 33411
rect 26097 33339 26103 33373
rect 26137 33339 26143 33373
rect 26097 33301 26143 33339
rect 26097 33267 26103 33301
rect 26137 33267 26143 33301
rect 26097 33229 26143 33267
rect 26097 33195 26103 33229
rect 26137 33195 26143 33229
rect 26097 33157 26143 33195
rect 26097 33123 26103 33157
rect 26137 33123 26143 33157
rect 26097 33085 26143 33123
rect 26097 33051 26103 33085
rect 26137 33051 26143 33085
rect 26097 33013 26143 33051
rect 26097 32979 26103 33013
rect 26137 32979 26143 33013
rect 26097 32941 26143 32979
rect 26097 32907 26103 32941
rect 26137 32907 26143 32941
rect 26097 32869 26143 32907
rect 26097 32835 26103 32869
rect 26137 32835 26143 32869
rect 26097 32797 26143 32835
rect 26097 32763 26103 32797
rect 26137 32763 26143 32797
rect 26097 32725 26143 32763
rect 26097 32691 26103 32725
rect 26137 32691 26143 32725
rect 26097 32653 26143 32691
rect 26097 32619 26103 32653
rect 26137 32619 26143 32653
rect 26097 32581 26143 32619
rect 26097 32547 26103 32581
rect 26137 32547 26143 32581
rect 26097 32509 26143 32547
rect 26097 32475 26103 32509
rect 26137 32475 26143 32509
rect 26097 32437 26143 32475
rect 26097 32403 26103 32437
rect 26137 32403 26143 32437
rect 26097 32387 26143 32403
rect 26555 33661 26601 33677
rect 26555 33627 26561 33661
rect 26595 33627 26601 33661
rect 26555 33589 26601 33627
rect 26555 33555 26561 33589
rect 26595 33555 26601 33589
rect 26555 33517 26601 33555
rect 26555 33483 26561 33517
rect 26595 33483 26601 33517
rect 26555 33445 26601 33483
rect 26555 33411 26561 33445
rect 26595 33411 26601 33445
rect 26555 33373 26601 33411
rect 26555 33339 26561 33373
rect 26595 33339 26601 33373
rect 26555 33301 26601 33339
rect 26555 33267 26561 33301
rect 26595 33267 26601 33301
rect 26555 33229 26601 33267
rect 26555 33195 26561 33229
rect 26595 33195 26601 33229
rect 26555 33157 26601 33195
rect 26555 33123 26561 33157
rect 26595 33123 26601 33157
rect 26555 33085 26601 33123
rect 26555 33051 26561 33085
rect 26595 33051 26601 33085
rect 26555 33013 26601 33051
rect 26555 32979 26561 33013
rect 26595 32979 26601 33013
rect 26555 32941 26601 32979
rect 26555 32907 26561 32941
rect 26595 32907 26601 32941
rect 26555 32869 26601 32907
rect 26555 32835 26561 32869
rect 26595 32835 26601 32869
rect 26555 32797 26601 32835
rect 26555 32763 26561 32797
rect 26595 32763 26601 32797
rect 26555 32725 26601 32763
rect 26555 32691 26561 32725
rect 26595 32691 26601 32725
rect 26555 32653 26601 32691
rect 26555 32619 26561 32653
rect 26595 32619 26601 32653
rect 26555 32581 26601 32619
rect 26555 32547 26561 32581
rect 26595 32547 26601 32581
rect 26555 32509 26601 32547
rect 26555 32475 26561 32509
rect 26595 32475 26601 32509
rect 26555 32437 26601 32475
rect 26555 32403 26561 32437
rect 26595 32403 26601 32437
rect 26555 32387 26601 32403
rect 27013 33661 27059 33677
rect 27013 33627 27019 33661
rect 27053 33627 27059 33661
rect 27013 33589 27059 33627
rect 27013 33555 27019 33589
rect 27053 33555 27059 33589
rect 27013 33517 27059 33555
rect 27013 33483 27019 33517
rect 27053 33483 27059 33517
rect 27013 33445 27059 33483
rect 27013 33411 27019 33445
rect 27053 33411 27059 33445
rect 27013 33373 27059 33411
rect 27013 33339 27019 33373
rect 27053 33339 27059 33373
rect 27013 33301 27059 33339
rect 27013 33267 27019 33301
rect 27053 33267 27059 33301
rect 27013 33229 27059 33267
rect 27013 33195 27019 33229
rect 27053 33195 27059 33229
rect 27013 33157 27059 33195
rect 27013 33123 27019 33157
rect 27053 33123 27059 33157
rect 27013 33085 27059 33123
rect 27013 33051 27019 33085
rect 27053 33051 27059 33085
rect 27013 33013 27059 33051
rect 27013 32979 27019 33013
rect 27053 32979 27059 33013
rect 27013 32941 27059 32979
rect 27013 32907 27019 32941
rect 27053 32907 27059 32941
rect 27013 32869 27059 32907
rect 27013 32835 27019 32869
rect 27053 32835 27059 32869
rect 27013 32797 27059 32835
rect 27013 32763 27019 32797
rect 27053 32763 27059 32797
rect 27013 32725 27059 32763
rect 27013 32691 27019 32725
rect 27053 32691 27059 32725
rect 27013 32653 27059 32691
rect 27013 32619 27019 32653
rect 27053 32619 27059 32653
rect 27013 32581 27059 32619
rect 27013 32547 27019 32581
rect 27053 32547 27059 32581
rect 27013 32509 27059 32547
rect 27013 32475 27019 32509
rect 27053 32475 27059 32509
rect 27013 32437 27059 32475
rect 27013 32403 27019 32437
rect 27053 32403 27059 32437
rect 27013 32387 27059 32403
rect 27471 33661 27517 33677
rect 27471 33627 27477 33661
rect 27511 33627 27517 33661
rect 27471 33589 27517 33627
rect 27471 33555 27477 33589
rect 27511 33555 27517 33589
rect 27471 33517 27517 33555
rect 27471 33483 27477 33517
rect 27511 33483 27517 33517
rect 27471 33445 27517 33483
rect 27471 33411 27477 33445
rect 27511 33411 27517 33445
rect 27471 33373 27517 33411
rect 27471 33339 27477 33373
rect 27511 33339 27517 33373
rect 27471 33301 27517 33339
rect 27471 33267 27477 33301
rect 27511 33267 27517 33301
rect 27471 33229 27517 33267
rect 27471 33195 27477 33229
rect 27511 33195 27517 33229
rect 27471 33157 27517 33195
rect 27471 33123 27477 33157
rect 27511 33123 27517 33157
rect 27471 33085 27517 33123
rect 27471 33051 27477 33085
rect 27511 33051 27517 33085
rect 27471 33013 27517 33051
rect 27471 32979 27477 33013
rect 27511 32979 27517 33013
rect 27471 32941 27517 32979
rect 27471 32907 27477 32941
rect 27511 32907 27517 32941
rect 27471 32869 27517 32907
rect 27471 32835 27477 32869
rect 27511 32835 27517 32869
rect 27471 32797 27517 32835
rect 27471 32763 27477 32797
rect 27511 32763 27517 32797
rect 27471 32725 27517 32763
rect 27471 32691 27477 32725
rect 27511 32691 27517 32725
rect 27471 32653 27517 32691
rect 27471 32619 27477 32653
rect 27511 32619 27517 32653
rect 27471 32581 27517 32619
rect 27471 32547 27477 32581
rect 27511 32547 27517 32581
rect 27471 32509 27517 32547
rect 27471 32475 27477 32509
rect 27511 32475 27517 32509
rect 27471 32437 27517 32475
rect 27471 32403 27477 32437
rect 27511 32403 27517 32437
rect 27471 32387 27517 32403
rect 27929 33661 27975 33677
rect 27929 33627 27935 33661
rect 27969 33627 27975 33661
rect 27929 33589 27975 33627
rect 27929 33555 27935 33589
rect 27969 33555 27975 33589
rect 27929 33517 27975 33555
rect 27929 33483 27935 33517
rect 27969 33483 27975 33517
rect 27929 33445 27975 33483
rect 27929 33411 27935 33445
rect 27969 33411 27975 33445
rect 27929 33373 27975 33411
rect 27929 33339 27935 33373
rect 27969 33339 27975 33373
rect 27929 33301 27975 33339
rect 27929 33267 27935 33301
rect 27969 33267 27975 33301
rect 27929 33229 27975 33267
rect 27929 33195 27935 33229
rect 27969 33195 27975 33229
rect 27929 33157 27975 33195
rect 27929 33123 27935 33157
rect 27969 33123 27975 33157
rect 27929 33085 27975 33123
rect 27929 33051 27935 33085
rect 27969 33051 27975 33085
rect 27929 33013 27975 33051
rect 27929 32979 27935 33013
rect 27969 32979 27975 33013
rect 27929 32941 27975 32979
rect 27929 32907 27935 32941
rect 27969 32907 27975 32941
rect 27929 32869 27975 32907
rect 27929 32835 27935 32869
rect 27969 32835 27975 32869
rect 27929 32797 27975 32835
rect 27929 32763 27935 32797
rect 27969 32763 27975 32797
rect 27929 32725 27975 32763
rect 27929 32691 27935 32725
rect 27969 32691 27975 32725
rect 27929 32653 27975 32691
rect 27929 32619 27935 32653
rect 27969 32619 27975 32653
rect 27929 32581 27975 32619
rect 27929 32547 27935 32581
rect 27969 32547 27975 32581
rect 27929 32509 27975 32547
rect 27929 32475 27935 32509
rect 27969 32475 27975 32509
rect 27929 32437 27975 32475
rect 27929 32403 27935 32437
rect 27969 32403 27975 32437
rect 27929 32387 27975 32403
rect 28387 33661 28433 33677
rect 28387 33627 28393 33661
rect 28427 33627 28433 33661
rect 28387 33589 28433 33627
rect 28387 33555 28393 33589
rect 28427 33555 28433 33589
rect 28387 33517 28433 33555
rect 28387 33483 28393 33517
rect 28427 33483 28433 33517
rect 28387 33445 28433 33483
rect 28387 33411 28393 33445
rect 28427 33411 28433 33445
rect 28387 33373 28433 33411
rect 28387 33339 28393 33373
rect 28427 33339 28433 33373
rect 28387 33301 28433 33339
rect 28387 33267 28393 33301
rect 28427 33267 28433 33301
rect 28387 33229 28433 33267
rect 28387 33195 28393 33229
rect 28427 33195 28433 33229
rect 28387 33157 28433 33195
rect 28387 33123 28393 33157
rect 28427 33123 28433 33157
rect 28387 33085 28433 33123
rect 28387 33051 28393 33085
rect 28427 33051 28433 33085
rect 28387 33013 28433 33051
rect 28387 32979 28393 33013
rect 28427 32979 28433 33013
rect 28387 32941 28433 32979
rect 28387 32907 28393 32941
rect 28427 32907 28433 32941
rect 28387 32869 28433 32907
rect 28387 32835 28393 32869
rect 28427 32835 28433 32869
rect 28387 32797 28433 32835
rect 28387 32763 28393 32797
rect 28427 32763 28433 32797
rect 28387 32725 28433 32763
rect 28387 32691 28393 32725
rect 28427 32691 28433 32725
rect 28387 32653 28433 32691
rect 28387 32619 28393 32653
rect 28427 32619 28433 32653
rect 28387 32581 28433 32619
rect 28387 32547 28393 32581
rect 28427 32547 28433 32581
rect 28387 32509 28433 32547
rect 28387 32475 28393 32509
rect 28427 32475 28433 32509
rect 28387 32437 28433 32475
rect 28387 32403 28393 32437
rect 28427 32403 28433 32437
rect 28387 32387 28433 32403
rect 28845 33661 28891 33677
rect 28845 33627 28851 33661
rect 28885 33627 28891 33661
rect 28845 33589 28891 33627
rect 28845 33555 28851 33589
rect 28885 33555 28891 33589
rect 28845 33517 28891 33555
rect 28845 33483 28851 33517
rect 28885 33483 28891 33517
rect 28845 33445 28891 33483
rect 28845 33411 28851 33445
rect 28885 33411 28891 33445
rect 28845 33373 28891 33411
rect 28845 33339 28851 33373
rect 28885 33339 28891 33373
rect 28845 33301 28891 33339
rect 28845 33267 28851 33301
rect 28885 33267 28891 33301
rect 28845 33229 28891 33267
rect 28845 33195 28851 33229
rect 28885 33195 28891 33229
rect 28845 33157 28891 33195
rect 28845 33123 28851 33157
rect 28885 33123 28891 33157
rect 28845 33085 28891 33123
rect 28845 33051 28851 33085
rect 28885 33051 28891 33085
rect 28845 33013 28891 33051
rect 28845 32979 28851 33013
rect 28885 32979 28891 33013
rect 28845 32941 28891 32979
rect 28845 32907 28851 32941
rect 28885 32907 28891 32941
rect 28845 32869 28891 32907
rect 28845 32835 28851 32869
rect 28885 32835 28891 32869
rect 28845 32797 28891 32835
rect 28845 32763 28851 32797
rect 28885 32763 28891 32797
rect 28845 32725 28891 32763
rect 28845 32691 28851 32725
rect 28885 32691 28891 32725
rect 28845 32653 28891 32691
rect 28845 32619 28851 32653
rect 28885 32619 28891 32653
rect 28845 32581 28891 32619
rect 28845 32547 28851 32581
rect 28885 32547 28891 32581
rect 28845 32509 28891 32547
rect 28845 32475 28851 32509
rect 28885 32475 28891 32509
rect 28845 32437 28891 32475
rect 28845 32403 28851 32437
rect 28885 32403 28891 32437
rect 28845 32387 28891 32403
rect 29303 33661 29349 33677
rect 29303 33627 29309 33661
rect 29343 33627 29349 33661
rect 29303 33589 29349 33627
rect 29303 33555 29309 33589
rect 29343 33555 29349 33589
rect 29303 33517 29349 33555
rect 29303 33483 29309 33517
rect 29343 33483 29349 33517
rect 29303 33445 29349 33483
rect 29303 33411 29309 33445
rect 29343 33411 29349 33445
rect 29303 33373 29349 33411
rect 29303 33339 29309 33373
rect 29343 33339 29349 33373
rect 29303 33301 29349 33339
rect 29303 33267 29309 33301
rect 29343 33267 29349 33301
rect 29303 33229 29349 33267
rect 29303 33195 29309 33229
rect 29343 33195 29349 33229
rect 29303 33157 29349 33195
rect 29303 33123 29309 33157
rect 29343 33123 29349 33157
rect 29303 33085 29349 33123
rect 29303 33051 29309 33085
rect 29343 33051 29349 33085
rect 29303 33013 29349 33051
rect 29303 32979 29309 33013
rect 29343 32979 29349 33013
rect 29303 32941 29349 32979
rect 29303 32907 29309 32941
rect 29343 32907 29349 32941
rect 29303 32869 29349 32907
rect 29303 32835 29309 32869
rect 29343 32835 29349 32869
rect 29303 32797 29349 32835
rect 29303 32763 29309 32797
rect 29343 32763 29349 32797
rect 29303 32725 29349 32763
rect 29303 32691 29309 32725
rect 29343 32691 29349 32725
rect 29303 32653 29349 32691
rect 29303 32619 29309 32653
rect 29343 32619 29349 32653
rect 29303 32581 29349 32619
rect 29303 32547 29309 32581
rect 29343 32547 29349 32581
rect 29303 32509 29349 32547
rect 29303 32475 29309 32509
rect 29343 32475 29349 32509
rect 29303 32437 29349 32475
rect 29303 32403 29309 32437
rect 29343 32403 29349 32437
rect 29303 32387 29349 32403
rect 29761 33661 29807 33677
rect 29761 33627 29767 33661
rect 29801 33627 29807 33661
rect 29761 33589 29807 33627
rect 29761 33555 29767 33589
rect 29801 33555 29807 33589
rect 29761 33517 29807 33555
rect 29761 33483 29767 33517
rect 29801 33483 29807 33517
rect 29761 33445 29807 33483
rect 29761 33411 29767 33445
rect 29801 33411 29807 33445
rect 29761 33373 29807 33411
rect 29761 33339 29767 33373
rect 29801 33339 29807 33373
rect 29761 33301 29807 33339
rect 29761 33267 29767 33301
rect 29801 33267 29807 33301
rect 29761 33229 29807 33267
rect 29761 33195 29767 33229
rect 29801 33195 29807 33229
rect 29761 33157 29807 33195
rect 29761 33123 29767 33157
rect 29801 33123 29807 33157
rect 29761 33085 29807 33123
rect 29761 33051 29767 33085
rect 29801 33051 29807 33085
rect 29761 33013 29807 33051
rect 29761 32979 29767 33013
rect 29801 32979 29807 33013
rect 29761 32941 29807 32979
rect 29761 32907 29767 32941
rect 29801 32907 29807 32941
rect 29761 32869 29807 32907
rect 29761 32835 29767 32869
rect 29801 32835 29807 32869
rect 29761 32797 29807 32835
rect 29761 32763 29767 32797
rect 29801 32763 29807 32797
rect 29761 32725 29807 32763
rect 29761 32691 29767 32725
rect 29801 32691 29807 32725
rect 29761 32653 29807 32691
rect 29761 32619 29767 32653
rect 29801 32619 29807 32653
rect 29761 32581 29807 32619
rect 29761 32547 29767 32581
rect 29801 32547 29807 32581
rect 29761 32509 29807 32547
rect 29761 32475 29767 32509
rect 29801 32475 29807 32509
rect 29761 32437 29807 32475
rect 29761 32403 29767 32437
rect 29801 32403 29807 32437
rect 29761 32387 29807 32403
rect 30219 33661 30265 33677
rect 30219 33627 30225 33661
rect 30259 33627 30265 33661
rect 30219 33589 30265 33627
rect 30219 33555 30225 33589
rect 30259 33555 30265 33589
rect 30219 33517 30265 33555
rect 30219 33483 30225 33517
rect 30259 33483 30265 33517
rect 30219 33445 30265 33483
rect 30219 33411 30225 33445
rect 30259 33411 30265 33445
rect 30219 33373 30265 33411
rect 30219 33339 30225 33373
rect 30259 33339 30265 33373
rect 30219 33301 30265 33339
rect 30219 33267 30225 33301
rect 30259 33267 30265 33301
rect 30219 33229 30265 33267
rect 30219 33195 30225 33229
rect 30259 33195 30265 33229
rect 30219 33157 30265 33195
rect 30219 33123 30225 33157
rect 30259 33123 30265 33157
rect 30219 33085 30265 33123
rect 30219 33051 30225 33085
rect 30259 33051 30265 33085
rect 30219 33013 30265 33051
rect 30219 32979 30225 33013
rect 30259 32979 30265 33013
rect 30219 32941 30265 32979
rect 30219 32907 30225 32941
rect 30259 32907 30265 32941
rect 30219 32869 30265 32907
rect 30219 32835 30225 32869
rect 30259 32835 30265 32869
rect 30219 32797 30265 32835
rect 30219 32763 30225 32797
rect 30259 32763 30265 32797
rect 30219 32725 30265 32763
rect 30219 32691 30225 32725
rect 30259 32691 30265 32725
rect 30219 32653 30265 32691
rect 30219 32619 30225 32653
rect 30259 32619 30265 32653
rect 30219 32581 30265 32619
rect 30219 32547 30225 32581
rect 30259 32547 30265 32581
rect 30219 32509 30265 32547
rect 30219 32475 30225 32509
rect 30259 32475 30265 32509
rect 30219 32437 30265 32475
rect 30219 32403 30225 32437
rect 30259 32403 30265 32437
rect 30219 32387 30265 32403
rect 30677 33661 30723 33677
rect 30677 33627 30683 33661
rect 30717 33627 30723 33661
rect 30677 33589 30723 33627
rect 30677 33555 30683 33589
rect 30717 33555 30723 33589
rect 30677 33517 30723 33555
rect 30677 33483 30683 33517
rect 30717 33483 30723 33517
rect 30677 33445 30723 33483
rect 30677 33411 30683 33445
rect 30717 33411 30723 33445
rect 30677 33373 30723 33411
rect 30677 33339 30683 33373
rect 30717 33339 30723 33373
rect 30677 33301 30723 33339
rect 30677 33267 30683 33301
rect 30717 33267 30723 33301
rect 30677 33229 30723 33267
rect 30677 33195 30683 33229
rect 30717 33195 30723 33229
rect 30677 33157 30723 33195
rect 30677 33123 30683 33157
rect 30717 33123 30723 33157
rect 30677 33085 30723 33123
rect 30677 33051 30683 33085
rect 30717 33051 30723 33085
rect 30677 33013 30723 33051
rect 30677 32979 30683 33013
rect 30717 32979 30723 33013
rect 30677 32941 30723 32979
rect 30677 32907 30683 32941
rect 30717 32907 30723 32941
rect 30677 32869 30723 32907
rect 30677 32835 30683 32869
rect 30717 32835 30723 32869
rect 30677 32797 30723 32835
rect 30677 32763 30683 32797
rect 30717 32763 30723 32797
rect 30677 32725 30723 32763
rect 30677 32691 30683 32725
rect 30717 32691 30723 32725
rect 30677 32653 30723 32691
rect 30677 32619 30683 32653
rect 30717 32619 30723 32653
rect 30677 32581 30723 32619
rect 30677 32547 30683 32581
rect 30717 32547 30723 32581
rect 30677 32509 30723 32547
rect 30677 32475 30683 32509
rect 30717 32475 30723 32509
rect 30677 32437 30723 32475
rect 30677 32403 30683 32437
rect 30717 32403 30723 32437
rect 30677 32387 30723 32403
rect 31135 33661 31181 33677
rect 31135 33627 31141 33661
rect 31175 33627 31181 33661
rect 31135 33589 31181 33627
rect 31135 33555 31141 33589
rect 31175 33555 31181 33589
rect 31135 33517 31181 33555
rect 31135 33483 31141 33517
rect 31175 33483 31181 33517
rect 31135 33445 31181 33483
rect 31135 33411 31141 33445
rect 31175 33411 31181 33445
rect 31135 33373 31181 33411
rect 31135 33339 31141 33373
rect 31175 33339 31181 33373
rect 31135 33301 31181 33339
rect 31135 33267 31141 33301
rect 31175 33267 31181 33301
rect 31135 33229 31181 33267
rect 31135 33195 31141 33229
rect 31175 33195 31181 33229
rect 31135 33157 31181 33195
rect 31135 33123 31141 33157
rect 31175 33123 31181 33157
rect 31135 33085 31181 33123
rect 31135 33051 31141 33085
rect 31175 33051 31181 33085
rect 31135 33013 31181 33051
rect 31135 32979 31141 33013
rect 31175 32979 31181 33013
rect 31135 32941 31181 32979
rect 31135 32907 31141 32941
rect 31175 32907 31181 32941
rect 31135 32869 31181 32907
rect 31135 32835 31141 32869
rect 31175 32835 31181 32869
rect 31135 32797 31181 32835
rect 31135 32763 31141 32797
rect 31175 32763 31181 32797
rect 31135 32725 31181 32763
rect 31135 32691 31141 32725
rect 31175 32691 31181 32725
rect 31135 32653 31181 32691
rect 31135 32619 31141 32653
rect 31175 32619 31181 32653
rect 31135 32581 31181 32619
rect 31135 32547 31141 32581
rect 31175 32547 31181 32581
rect 31135 32509 31181 32547
rect 31135 32475 31141 32509
rect 31175 32475 31181 32509
rect 31135 32437 31181 32475
rect 31135 32403 31141 32437
rect 31175 32403 31181 32437
rect 31135 32387 31181 32403
rect 31593 33661 31639 33677
rect 31593 33627 31599 33661
rect 31633 33627 31639 33661
rect 31593 33589 31639 33627
rect 31593 33555 31599 33589
rect 31633 33555 31639 33589
rect 31593 33517 31639 33555
rect 31593 33483 31599 33517
rect 31633 33483 31639 33517
rect 31593 33445 31639 33483
rect 31593 33411 31599 33445
rect 31633 33411 31639 33445
rect 31593 33373 31639 33411
rect 31593 33339 31599 33373
rect 31633 33339 31639 33373
rect 31593 33301 31639 33339
rect 31593 33267 31599 33301
rect 31633 33267 31639 33301
rect 31593 33229 31639 33267
rect 31593 33195 31599 33229
rect 31633 33195 31639 33229
rect 31593 33157 31639 33195
rect 31593 33123 31599 33157
rect 31633 33123 31639 33157
rect 31593 33085 31639 33123
rect 31593 33051 31599 33085
rect 31633 33051 31639 33085
rect 31593 33013 31639 33051
rect 31593 32979 31599 33013
rect 31633 32979 31639 33013
rect 31593 32941 31639 32979
rect 31593 32907 31599 32941
rect 31633 32907 31639 32941
rect 31593 32869 31639 32907
rect 31593 32835 31599 32869
rect 31633 32835 31639 32869
rect 31593 32797 31639 32835
rect 31593 32763 31599 32797
rect 31633 32763 31639 32797
rect 31593 32725 31639 32763
rect 31593 32691 31599 32725
rect 31633 32691 31639 32725
rect 31593 32653 31639 32691
rect 31593 32619 31599 32653
rect 31633 32619 31639 32653
rect 31593 32581 31639 32619
rect 31593 32547 31599 32581
rect 31633 32547 31639 32581
rect 31593 32509 31639 32547
rect 31593 32475 31599 32509
rect 31633 32475 31639 32509
rect 31593 32437 31639 32475
rect 31593 32403 31599 32437
rect 31633 32403 31639 32437
rect 31593 32387 31639 32403
rect 32051 33661 32097 33677
rect 32051 33627 32057 33661
rect 32091 33627 32097 33661
rect 32051 33589 32097 33627
rect 32051 33555 32057 33589
rect 32091 33555 32097 33589
rect 32051 33517 32097 33555
rect 32051 33483 32057 33517
rect 32091 33483 32097 33517
rect 32051 33445 32097 33483
rect 32051 33411 32057 33445
rect 32091 33411 32097 33445
rect 32051 33373 32097 33411
rect 32051 33339 32057 33373
rect 32091 33339 32097 33373
rect 32051 33301 32097 33339
rect 32051 33267 32057 33301
rect 32091 33267 32097 33301
rect 32051 33229 32097 33267
rect 32051 33195 32057 33229
rect 32091 33195 32097 33229
rect 32051 33157 32097 33195
rect 32051 33123 32057 33157
rect 32091 33123 32097 33157
rect 32051 33085 32097 33123
rect 32051 33051 32057 33085
rect 32091 33051 32097 33085
rect 32051 33013 32097 33051
rect 32051 32979 32057 33013
rect 32091 32979 32097 33013
rect 32051 32941 32097 32979
rect 32051 32907 32057 32941
rect 32091 32907 32097 32941
rect 32051 32869 32097 32907
rect 32051 32835 32057 32869
rect 32091 32835 32097 32869
rect 32051 32797 32097 32835
rect 32051 32763 32057 32797
rect 32091 32763 32097 32797
rect 32051 32725 32097 32763
rect 32051 32691 32057 32725
rect 32091 32691 32097 32725
rect 32051 32653 32097 32691
rect 32051 32619 32057 32653
rect 32091 32619 32097 32653
rect 32051 32581 32097 32619
rect 32051 32547 32057 32581
rect 32091 32547 32097 32581
rect 32051 32509 32097 32547
rect 32051 32475 32057 32509
rect 32091 32475 32097 32509
rect 32051 32437 32097 32475
rect 32051 32403 32057 32437
rect 32091 32403 32097 32437
rect 32051 32387 32097 32403
rect 32509 33661 32555 33677
rect 32509 33627 32515 33661
rect 32549 33627 32555 33661
rect 32509 33589 32555 33627
rect 32509 33555 32515 33589
rect 32549 33555 32555 33589
rect 32509 33517 32555 33555
rect 32509 33483 32515 33517
rect 32549 33483 32555 33517
rect 32509 33445 32555 33483
rect 32509 33411 32515 33445
rect 32549 33411 32555 33445
rect 32509 33373 32555 33411
rect 32509 33339 32515 33373
rect 32549 33339 32555 33373
rect 32509 33301 32555 33339
rect 32509 33267 32515 33301
rect 32549 33267 32555 33301
rect 32509 33229 32555 33267
rect 32509 33195 32515 33229
rect 32549 33195 32555 33229
rect 32509 33157 32555 33195
rect 32509 33123 32515 33157
rect 32549 33123 32555 33157
rect 32509 33085 32555 33123
rect 32509 33051 32515 33085
rect 32549 33051 32555 33085
rect 32509 33013 32555 33051
rect 32509 32979 32515 33013
rect 32549 32979 32555 33013
rect 32509 32941 32555 32979
rect 32509 32907 32515 32941
rect 32549 32907 32555 32941
rect 32509 32869 32555 32907
rect 32509 32835 32515 32869
rect 32549 32835 32555 32869
rect 32509 32797 32555 32835
rect 32509 32763 32515 32797
rect 32549 32763 32555 32797
rect 32509 32725 32555 32763
rect 32509 32691 32515 32725
rect 32549 32691 32555 32725
rect 32509 32653 32555 32691
rect 32509 32619 32515 32653
rect 32549 32619 32555 32653
rect 32509 32581 32555 32619
rect 32509 32547 32515 32581
rect 32549 32547 32555 32581
rect 32509 32509 32555 32547
rect 32509 32475 32515 32509
rect 32549 32475 32555 32509
rect 32509 32437 32555 32475
rect 32509 32403 32515 32437
rect 32549 32403 32555 32437
rect 32509 32387 32555 32403
rect 32967 33661 33013 33677
rect 32967 33627 32973 33661
rect 33007 33627 33013 33661
rect 32967 33589 33013 33627
rect 32967 33555 32973 33589
rect 33007 33555 33013 33589
rect 32967 33517 33013 33555
rect 32967 33483 32973 33517
rect 33007 33483 33013 33517
rect 32967 33445 33013 33483
rect 32967 33411 32973 33445
rect 33007 33411 33013 33445
rect 32967 33373 33013 33411
rect 32967 33339 32973 33373
rect 33007 33339 33013 33373
rect 32967 33301 33013 33339
rect 32967 33267 32973 33301
rect 33007 33267 33013 33301
rect 32967 33229 33013 33267
rect 32967 33195 32973 33229
rect 33007 33195 33013 33229
rect 32967 33157 33013 33195
rect 32967 33123 32973 33157
rect 33007 33123 33013 33157
rect 32967 33085 33013 33123
rect 32967 33051 32973 33085
rect 33007 33051 33013 33085
rect 32967 33013 33013 33051
rect 32967 32979 32973 33013
rect 33007 32979 33013 33013
rect 32967 32941 33013 32979
rect 32967 32907 32973 32941
rect 33007 32907 33013 32941
rect 32967 32869 33013 32907
rect 32967 32835 32973 32869
rect 33007 32835 33013 32869
rect 32967 32797 33013 32835
rect 32967 32763 32973 32797
rect 33007 32763 33013 32797
rect 32967 32725 33013 32763
rect 32967 32691 32973 32725
rect 33007 32691 33013 32725
rect 32967 32653 33013 32691
rect 32967 32619 32973 32653
rect 33007 32619 33013 32653
rect 32967 32581 33013 32619
rect 32967 32547 32973 32581
rect 33007 32547 33013 32581
rect 32967 32509 33013 32547
rect 32967 32475 32973 32509
rect 33007 32475 33013 32509
rect 32967 32437 33013 32475
rect 32967 32403 32973 32437
rect 33007 32403 33013 32437
rect 32967 32387 33013 32403
rect 33425 33661 33471 33677
rect 33425 33627 33431 33661
rect 33465 33627 33471 33661
rect 33425 33589 33471 33627
rect 33425 33555 33431 33589
rect 33465 33555 33471 33589
rect 33425 33517 33471 33555
rect 33425 33483 33431 33517
rect 33465 33483 33471 33517
rect 33425 33445 33471 33483
rect 33425 33411 33431 33445
rect 33465 33411 33471 33445
rect 33425 33373 33471 33411
rect 33425 33339 33431 33373
rect 33465 33339 33471 33373
rect 33425 33301 33471 33339
rect 33425 33267 33431 33301
rect 33465 33267 33471 33301
rect 33425 33229 33471 33267
rect 33425 33195 33431 33229
rect 33465 33195 33471 33229
rect 33425 33157 33471 33195
rect 33425 33123 33431 33157
rect 33465 33123 33471 33157
rect 33425 33085 33471 33123
rect 33425 33051 33431 33085
rect 33465 33051 33471 33085
rect 33425 33013 33471 33051
rect 33425 32979 33431 33013
rect 33465 32979 33471 33013
rect 33425 32941 33471 32979
rect 33425 32907 33431 32941
rect 33465 32907 33471 32941
rect 33425 32869 33471 32907
rect 33425 32835 33431 32869
rect 33465 32835 33471 32869
rect 33425 32797 33471 32835
rect 33425 32763 33431 32797
rect 33465 32763 33471 32797
rect 33425 32725 33471 32763
rect 33425 32691 33431 32725
rect 33465 32691 33471 32725
rect 33425 32653 33471 32691
rect 33425 32619 33431 32653
rect 33465 32619 33471 32653
rect 33425 32581 33471 32619
rect 33425 32547 33431 32581
rect 33465 32547 33471 32581
rect 33425 32509 33471 32547
rect 33425 32475 33431 32509
rect 33465 32475 33471 32509
rect 33425 32437 33471 32475
rect 33425 32403 33431 32437
rect 33465 32403 33471 32437
rect 33425 32387 33471 32403
rect 33883 33661 33929 33677
rect 33883 33627 33889 33661
rect 33923 33627 33929 33661
rect 33883 33589 33929 33627
rect 33883 33555 33889 33589
rect 33923 33555 33929 33589
rect 33883 33517 33929 33555
rect 33883 33483 33889 33517
rect 33923 33483 33929 33517
rect 33883 33445 33929 33483
rect 33883 33411 33889 33445
rect 33923 33411 33929 33445
rect 33883 33373 33929 33411
rect 33883 33339 33889 33373
rect 33923 33339 33929 33373
rect 33883 33301 33929 33339
rect 33883 33267 33889 33301
rect 33923 33267 33929 33301
rect 33883 33229 33929 33267
rect 33883 33195 33889 33229
rect 33923 33195 33929 33229
rect 33883 33157 33929 33195
rect 33883 33123 33889 33157
rect 33923 33123 33929 33157
rect 33883 33085 33929 33123
rect 33883 33051 33889 33085
rect 33923 33051 33929 33085
rect 33883 33013 33929 33051
rect 33883 32979 33889 33013
rect 33923 32979 33929 33013
rect 33883 32941 33929 32979
rect 33883 32907 33889 32941
rect 33923 32907 33929 32941
rect 33883 32869 33929 32907
rect 33883 32835 33889 32869
rect 33923 32835 33929 32869
rect 33883 32797 33929 32835
rect 33883 32763 33889 32797
rect 33923 32763 33929 32797
rect 33883 32725 33929 32763
rect 33883 32691 33889 32725
rect 33923 32691 33929 32725
rect 33883 32653 33929 32691
rect 33883 32619 33889 32653
rect 33923 32619 33929 32653
rect 33883 32581 33929 32619
rect 33883 32547 33889 32581
rect 33923 32547 33929 32581
rect 33883 32509 33929 32547
rect 33883 32475 33889 32509
rect 33923 32475 33929 32509
rect 33883 32437 33929 32475
rect 33883 32403 33889 32437
rect 33923 32403 33929 32437
rect 33883 32387 33929 32403
rect 34341 33661 34387 33677
rect 34341 33627 34347 33661
rect 34381 33627 34387 33661
rect 34341 33589 34387 33627
rect 34341 33555 34347 33589
rect 34381 33555 34387 33589
rect 34341 33517 34387 33555
rect 34341 33483 34347 33517
rect 34381 33483 34387 33517
rect 34341 33445 34387 33483
rect 34341 33411 34347 33445
rect 34381 33411 34387 33445
rect 34341 33373 34387 33411
rect 34341 33339 34347 33373
rect 34381 33339 34387 33373
rect 34341 33301 34387 33339
rect 34341 33267 34347 33301
rect 34381 33267 34387 33301
rect 34341 33229 34387 33267
rect 34341 33195 34347 33229
rect 34381 33195 34387 33229
rect 34341 33157 34387 33195
rect 34341 33123 34347 33157
rect 34381 33123 34387 33157
rect 34341 33085 34387 33123
rect 34341 33051 34347 33085
rect 34381 33051 34387 33085
rect 34341 33013 34387 33051
rect 34341 32979 34347 33013
rect 34381 32979 34387 33013
rect 34341 32941 34387 32979
rect 34341 32907 34347 32941
rect 34381 32907 34387 32941
rect 34341 32869 34387 32907
rect 34341 32835 34347 32869
rect 34381 32835 34387 32869
rect 34341 32797 34387 32835
rect 34341 32763 34347 32797
rect 34381 32763 34387 32797
rect 34341 32725 34387 32763
rect 34341 32691 34347 32725
rect 34381 32691 34387 32725
rect 34341 32653 34387 32691
rect 34341 32619 34347 32653
rect 34381 32619 34387 32653
rect 34341 32581 34387 32619
rect 34341 32547 34347 32581
rect 34381 32547 34387 32581
rect 34341 32509 34387 32547
rect 34341 32475 34347 32509
rect 34381 32475 34387 32509
rect 34341 32437 34387 32475
rect 34341 32403 34347 32437
rect 34381 32403 34387 32437
rect 34341 32387 34387 32403
rect 34799 33661 34845 33677
rect 34799 33627 34805 33661
rect 34839 33627 34845 33661
rect 34799 33589 34845 33627
rect 34799 33555 34805 33589
rect 34839 33555 34845 33589
rect 34799 33517 34845 33555
rect 34799 33483 34805 33517
rect 34839 33483 34845 33517
rect 34799 33445 34845 33483
rect 34799 33411 34805 33445
rect 34839 33411 34845 33445
rect 34799 33373 34845 33411
rect 34799 33339 34805 33373
rect 34839 33339 34845 33373
rect 34799 33301 34845 33339
rect 34799 33267 34805 33301
rect 34839 33267 34845 33301
rect 34799 33229 34845 33267
rect 34799 33195 34805 33229
rect 34839 33195 34845 33229
rect 34799 33157 34845 33195
rect 34799 33123 34805 33157
rect 34839 33123 34845 33157
rect 34799 33085 34845 33123
rect 34799 33051 34805 33085
rect 34839 33051 34845 33085
rect 34799 33013 34845 33051
rect 34799 32979 34805 33013
rect 34839 32979 34845 33013
rect 34799 32941 34845 32979
rect 34799 32907 34805 32941
rect 34839 32907 34845 32941
rect 34799 32869 34845 32907
rect 34799 32835 34805 32869
rect 34839 32835 34845 32869
rect 34799 32797 34845 32835
rect 34799 32763 34805 32797
rect 34839 32763 34845 32797
rect 34799 32725 34845 32763
rect 34799 32691 34805 32725
rect 34839 32691 34845 32725
rect 34799 32653 34845 32691
rect 34799 32619 34805 32653
rect 34839 32619 34845 32653
rect 34799 32581 34845 32619
rect 34799 32547 34805 32581
rect 34839 32547 34845 32581
rect 34799 32509 34845 32547
rect 34799 32475 34805 32509
rect 34839 32475 34845 32509
rect 34799 32437 34845 32475
rect 34799 32403 34805 32437
rect 34839 32403 34845 32437
rect 34799 32387 34845 32403
rect 35257 33661 35303 33677
rect 35257 33627 35263 33661
rect 35297 33627 35303 33661
rect 35257 33589 35303 33627
rect 35257 33555 35263 33589
rect 35297 33555 35303 33589
rect 35257 33517 35303 33555
rect 35257 33483 35263 33517
rect 35297 33483 35303 33517
rect 35257 33445 35303 33483
rect 35257 33411 35263 33445
rect 35297 33411 35303 33445
rect 35257 33373 35303 33411
rect 35257 33339 35263 33373
rect 35297 33339 35303 33373
rect 35257 33301 35303 33339
rect 35257 33267 35263 33301
rect 35297 33267 35303 33301
rect 35257 33229 35303 33267
rect 35257 33195 35263 33229
rect 35297 33195 35303 33229
rect 35257 33157 35303 33195
rect 35257 33123 35263 33157
rect 35297 33123 35303 33157
rect 35257 33085 35303 33123
rect 35257 33051 35263 33085
rect 35297 33051 35303 33085
rect 35257 33013 35303 33051
rect 35257 32979 35263 33013
rect 35297 32979 35303 33013
rect 35257 32941 35303 32979
rect 35257 32907 35263 32941
rect 35297 32907 35303 32941
rect 35257 32869 35303 32907
rect 35257 32835 35263 32869
rect 35297 32835 35303 32869
rect 35257 32797 35303 32835
rect 35257 32763 35263 32797
rect 35297 32763 35303 32797
rect 35257 32725 35303 32763
rect 35257 32691 35263 32725
rect 35297 32691 35303 32725
rect 35257 32653 35303 32691
rect 35257 32619 35263 32653
rect 35297 32619 35303 32653
rect 35257 32581 35303 32619
rect 35257 32547 35263 32581
rect 35297 32547 35303 32581
rect 35257 32509 35303 32547
rect 35257 32475 35263 32509
rect 35297 32475 35303 32509
rect 35257 32437 35303 32475
rect 35257 32403 35263 32437
rect 35297 32403 35303 32437
rect 35257 32387 35303 32403
rect 35715 33661 35761 33677
rect 35715 33627 35721 33661
rect 35755 33627 35761 33661
rect 35715 33589 35761 33627
rect 35715 33555 35721 33589
rect 35755 33555 35761 33589
rect 35715 33517 35761 33555
rect 35715 33483 35721 33517
rect 35755 33483 35761 33517
rect 35715 33445 35761 33483
rect 35715 33411 35721 33445
rect 35755 33411 35761 33445
rect 35715 33373 35761 33411
rect 35715 33339 35721 33373
rect 35755 33339 35761 33373
rect 35715 33301 35761 33339
rect 35715 33267 35721 33301
rect 35755 33267 35761 33301
rect 35715 33229 35761 33267
rect 35715 33195 35721 33229
rect 35755 33195 35761 33229
rect 35715 33157 35761 33195
rect 35715 33123 35721 33157
rect 35755 33123 35761 33157
rect 35715 33085 35761 33123
rect 35715 33051 35721 33085
rect 35755 33051 35761 33085
rect 35715 33013 35761 33051
rect 35715 32979 35721 33013
rect 35755 32979 35761 33013
rect 35715 32941 35761 32979
rect 35715 32907 35721 32941
rect 35755 32907 35761 32941
rect 35715 32869 35761 32907
rect 35715 32835 35721 32869
rect 35755 32835 35761 32869
rect 35715 32797 35761 32835
rect 35715 32763 35721 32797
rect 35755 32763 35761 32797
rect 35715 32725 35761 32763
rect 35715 32691 35721 32725
rect 35755 32691 35761 32725
rect 35715 32653 35761 32691
rect 35715 32619 35721 32653
rect 35755 32619 35761 32653
rect 35715 32581 35761 32619
rect 35715 32547 35721 32581
rect 35755 32547 35761 32581
rect 35715 32509 35761 32547
rect 35715 32475 35721 32509
rect 35755 32475 35761 32509
rect 35715 32437 35761 32475
rect 35715 32403 35721 32437
rect 35755 32403 35761 32437
rect 35715 32387 35761 32403
rect 36173 33661 36219 33677
rect 36173 33627 36179 33661
rect 36213 33627 36219 33661
rect 36173 33589 36219 33627
rect 36173 33555 36179 33589
rect 36213 33555 36219 33589
rect 36173 33517 36219 33555
rect 36173 33483 36179 33517
rect 36213 33483 36219 33517
rect 36173 33445 36219 33483
rect 36173 33411 36179 33445
rect 36213 33411 36219 33445
rect 36173 33373 36219 33411
rect 36173 33339 36179 33373
rect 36213 33339 36219 33373
rect 36173 33301 36219 33339
rect 36173 33267 36179 33301
rect 36213 33267 36219 33301
rect 36173 33229 36219 33267
rect 36173 33195 36179 33229
rect 36213 33195 36219 33229
rect 36173 33157 36219 33195
rect 36173 33123 36179 33157
rect 36213 33123 36219 33157
rect 36173 33085 36219 33123
rect 36173 33051 36179 33085
rect 36213 33051 36219 33085
rect 36173 33013 36219 33051
rect 36173 32979 36179 33013
rect 36213 32979 36219 33013
rect 36173 32941 36219 32979
rect 36173 32907 36179 32941
rect 36213 32907 36219 32941
rect 36173 32869 36219 32907
rect 36173 32835 36179 32869
rect 36213 32835 36219 32869
rect 36173 32797 36219 32835
rect 36173 32763 36179 32797
rect 36213 32763 36219 32797
rect 36173 32725 36219 32763
rect 36173 32691 36179 32725
rect 36213 32691 36219 32725
rect 36173 32653 36219 32691
rect 36173 32619 36179 32653
rect 36213 32619 36219 32653
rect 36173 32581 36219 32619
rect 36173 32547 36179 32581
rect 36213 32547 36219 32581
rect 36173 32509 36219 32547
rect 36173 32475 36179 32509
rect 36213 32475 36219 32509
rect 36173 32437 36219 32475
rect 36173 32403 36179 32437
rect 36213 32403 36219 32437
rect 36173 32387 36219 32403
rect 36631 33661 36677 33677
rect 36631 33627 36637 33661
rect 36671 33627 36677 33661
rect 36631 33589 36677 33627
rect 36631 33555 36637 33589
rect 36671 33555 36677 33589
rect 36631 33517 36677 33555
rect 36631 33483 36637 33517
rect 36671 33483 36677 33517
rect 36631 33445 36677 33483
rect 36631 33411 36637 33445
rect 36671 33411 36677 33445
rect 36631 33373 36677 33411
rect 36631 33339 36637 33373
rect 36671 33339 36677 33373
rect 36631 33301 36677 33339
rect 36631 33267 36637 33301
rect 36671 33267 36677 33301
rect 36631 33229 36677 33267
rect 36631 33195 36637 33229
rect 36671 33195 36677 33229
rect 36631 33157 36677 33195
rect 36631 33123 36637 33157
rect 36671 33123 36677 33157
rect 36631 33085 36677 33123
rect 36631 33051 36637 33085
rect 36671 33051 36677 33085
rect 36631 33013 36677 33051
rect 36631 32979 36637 33013
rect 36671 32979 36677 33013
rect 36631 32941 36677 32979
rect 36631 32907 36637 32941
rect 36671 32907 36677 32941
rect 36631 32869 36677 32907
rect 36631 32835 36637 32869
rect 36671 32835 36677 32869
rect 36631 32797 36677 32835
rect 36631 32763 36637 32797
rect 36671 32763 36677 32797
rect 36631 32725 36677 32763
rect 36631 32691 36637 32725
rect 36671 32691 36677 32725
rect 36631 32653 36677 32691
rect 36631 32619 36637 32653
rect 36671 32619 36677 32653
rect 36631 32581 36677 32619
rect 36631 32547 36637 32581
rect 36671 32547 36677 32581
rect 36631 32509 36677 32547
rect 36631 32475 36637 32509
rect 36671 32475 36677 32509
rect 36631 32437 36677 32475
rect 36631 32403 36637 32437
rect 36671 32403 36677 32437
rect 36631 32387 36677 32403
rect 37089 33661 37135 33677
rect 37089 33627 37095 33661
rect 37129 33627 37135 33661
rect 37089 33589 37135 33627
rect 37089 33555 37095 33589
rect 37129 33555 37135 33589
rect 37089 33517 37135 33555
rect 37089 33483 37095 33517
rect 37129 33483 37135 33517
rect 37089 33445 37135 33483
rect 37089 33411 37095 33445
rect 37129 33411 37135 33445
rect 37089 33373 37135 33411
rect 37089 33339 37095 33373
rect 37129 33339 37135 33373
rect 37089 33301 37135 33339
rect 37089 33267 37095 33301
rect 37129 33267 37135 33301
rect 37089 33229 37135 33267
rect 37089 33195 37095 33229
rect 37129 33195 37135 33229
rect 37089 33157 37135 33195
rect 37089 33123 37095 33157
rect 37129 33123 37135 33157
rect 37089 33085 37135 33123
rect 37089 33051 37095 33085
rect 37129 33051 37135 33085
rect 37089 33013 37135 33051
rect 37089 32979 37095 33013
rect 37129 32979 37135 33013
rect 37089 32941 37135 32979
rect 37089 32907 37095 32941
rect 37129 32907 37135 32941
rect 37089 32869 37135 32907
rect 37089 32835 37095 32869
rect 37129 32835 37135 32869
rect 37089 32797 37135 32835
rect 37089 32763 37095 32797
rect 37129 32763 37135 32797
rect 37089 32725 37135 32763
rect 37089 32691 37095 32725
rect 37129 32691 37135 32725
rect 37089 32653 37135 32691
rect 37089 32619 37095 32653
rect 37129 32619 37135 32653
rect 37089 32581 37135 32619
rect 37089 32547 37095 32581
rect 37129 32547 37135 32581
rect 37089 32509 37135 32547
rect 37089 32475 37095 32509
rect 37129 32475 37135 32509
rect 37089 32437 37135 32475
rect 37089 32403 37095 32437
rect 37129 32403 37135 32437
rect 37089 32387 37135 32403
rect 37547 33661 37593 33677
rect 37547 33627 37553 33661
rect 37587 33627 37593 33661
rect 37547 33589 37593 33627
rect 37547 33555 37553 33589
rect 37587 33555 37593 33589
rect 37547 33517 37593 33555
rect 37547 33483 37553 33517
rect 37587 33483 37593 33517
rect 37547 33445 37593 33483
rect 37547 33411 37553 33445
rect 37587 33411 37593 33445
rect 37547 33373 37593 33411
rect 37547 33339 37553 33373
rect 37587 33339 37593 33373
rect 37547 33301 37593 33339
rect 37547 33267 37553 33301
rect 37587 33267 37593 33301
rect 37547 33229 37593 33267
rect 37547 33195 37553 33229
rect 37587 33195 37593 33229
rect 37547 33157 37593 33195
rect 37547 33123 37553 33157
rect 37587 33123 37593 33157
rect 37547 33085 37593 33123
rect 37547 33051 37553 33085
rect 37587 33051 37593 33085
rect 37547 33013 37593 33051
rect 37547 32979 37553 33013
rect 37587 32979 37593 33013
rect 37547 32941 37593 32979
rect 37547 32907 37553 32941
rect 37587 32907 37593 32941
rect 37547 32869 37593 32907
rect 37547 32835 37553 32869
rect 37587 32835 37593 32869
rect 37547 32797 37593 32835
rect 37547 32763 37553 32797
rect 37587 32763 37593 32797
rect 37547 32725 37593 32763
rect 37547 32691 37553 32725
rect 37587 32691 37593 32725
rect 37547 32653 37593 32691
rect 37547 32619 37553 32653
rect 37587 32619 37593 32653
rect 37547 32581 37593 32619
rect 37547 32547 37553 32581
rect 37587 32547 37593 32581
rect 37547 32509 37593 32547
rect 37547 32475 37553 32509
rect 37587 32475 37593 32509
rect 37547 32437 37593 32475
rect 37547 32403 37553 32437
rect 37587 32403 37593 32437
rect 37547 32387 37593 32403
rect 38005 33661 38051 33677
rect 38005 33627 38011 33661
rect 38045 33627 38051 33661
rect 38005 33589 38051 33627
rect 38005 33555 38011 33589
rect 38045 33555 38051 33589
rect 38005 33517 38051 33555
rect 38005 33483 38011 33517
rect 38045 33483 38051 33517
rect 38005 33445 38051 33483
rect 38005 33411 38011 33445
rect 38045 33411 38051 33445
rect 38005 33373 38051 33411
rect 38005 33339 38011 33373
rect 38045 33339 38051 33373
rect 38005 33301 38051 33339
rect 38005 33267 38011 33301
rect 38045 33267 38051 33301
rect 38005 33229 38051 33267
rect 38005 33195 38011 33229
rect 38045 33195 38051 33229
rect 38005 33157 38051 33195
rect 38005 33123 38011 33157
rect 38045 33123 38051 33157
rect 38005 33085 38051 33123
rect 38005 33051 38011 33085
rect 38045 33051 38051 33085
rect 38005 33013 38051 33051
rect 38005 32979 38011 33013
rect 38045 32979 38051 33013
rect 38005 32941 38051 32979
rect 38005 32907 38011 32941
rect 38045 32907 38051 32941
rect 38005 32869 38051 32907
rect 38005 32835 38011 32869
rect 38045 32835 38051 32869
rect 38005 32797 38051 32835
rect 38005 32763 38011 32797
rect 38045 32763 38051 32797
rect 38005 32725 38051 32763
rect 38005 32691 38011 32725
rect 38045 32691 38051 32725
rect 38005 32653 38051 32691
rect 38005 32619 38011 32653
rect 38045 32619 38051 32653
rect 38005 32581 38051 32619
rect 38005 32547 38011 32581
rect 38045 32547 38051 32581
rect 38005 32509 38051 32547
rect 38005 32475 38011 32509
rect 38045 32475 38051 32509
rect 38005 32437 38051 32475
rect 38005 32403 38011 32437
rect 38045 32403 38051 32437
rect 38005 32387 38051 32403
rect 38463 33661 38509 33677
rect 38463 33627 38469 33661
rect 38503 33627 38509 33661
rect 38463 33589 38509 33627
rect 38463 33555 38469 33589
rect 38503 33555 38509 33589
rect 38463 33517 38509 33555
rect 38463 33483 38469 33517
rect 38503 33483 38509 33517
rect 38463 33445 38509 33483
rect 38463 33411 38469 33445
rect 38503 33411 38509 33445
rect 38463 33373 38509 33411
rect 38463 33339 38469 33373
rect 38503 33339 38509 33373
rect 38463 33301 38509 33339
rect 38463 33267 38469 33301
rect 38503 33267 38509 33301
rect 38463 33229 38509 33267
rect 38463 33195 38469 33229
rect 38503 33195 38509 33229
rect 38463 33157 38509 33195
rect 38463 33123 38469 33157
rect 38503 33123 38509 33157
rect 38463 33085 38509 33123
rect 38463 33051 38469 33085
rect 38503 33051 38509 33085
rect 38463 33013 38509 33051
rect 38463 32979 38469 33013
rect 38503 32979 38509 33013
rect 38463 32941 38509 32979
rect 38463 32907 38469 32941
rect 38503 32907 38509 32941
rect 38463 32869 38509 32907
rect 38463 32835 38469 32869
rect 38503 32835 38509 32869
rect 38463 32797 38509 32835
rect 38463 32763 38469 32797
rect 38503 32763 38509 32797
rect 38463 32725 38509 32763
rect 38463 32691 38469 32725
rect 38503 32691 38509 32725
rect 38463 32653 38509 32691
rect 38463 32619 38469 32653
rect 38503 32619 38509 32653
rect 38463 32581 38509 32619
rect 38463 32547 38469 32581
rect 38503 32547 38509 32581
rect 38463 32509 38509 32547
rect 38463 32475 38469 32509
rect 38503 32475 38509 32509
rect 38463 32437 38509 32475
rect 38463 32403 38469 32437
rect 38503 32403 38509 32437
rect 38463 32387 38509 32403
rect 38921 33661 38967 33677
rect 38921 33627 38927 33661
rect 38961 33627 38967 33661
rect 38921 33589 38967 33627
rect 38921 33555 38927 33589
rect 38961 33555 38967 33589
rect 38921 33517 38967 33555
rect 38921 33483 38927 33517
rect 38961 33483 38967 33517
rect 38921 33445 38967 33483
rect 38921 33411 38927 33445
rect 38961 33411 38967 33445
rect 38921 33373 38967 33411
rect 38921 33339 38927 33373
rect 38961 33339 38967 33373
rect 38921 33301 38967 33339
rect 38921 33267 38927 33301
rect 38961 33267 38967 33301
rect 38921 33229 38967 33267
rect 38921 33195 38927 33229
rect 38961 33195 38967 33229
rect 38921 33157 38967 33195
rect 38921 33123 38927 33157
rect 38961 33123 38967 33157
rect 38921 33085 38967 33123
rect 38921 33051 38927 33085
rect 38961 33051 38967 33085
rect 38921 33013 38967 33051
rect 38921 32979 38927 33013
rect 38961 32979 38967 33013
rect 38921 32941 38967 32979
rect 38921 32907 38927 32941
rect 38961 32907 38967 32941
rect 38921 32869 38967 32907
rect 38921 32835 38927 32869
rect 38961 32835 38967 32869
rect 38921 32797 38967 32835
rect 38921 32763 38927 32797
rect 38961 32763 38967 32797
rect 38921 32725 38967 32763
rect 38921 32691 38927 32725
rect 38961 32691 38967 32725
rect 38921 32653 38967 32691
rect 38921 32619 38927 32653
rect 38961 32619 38967 32653
rect 38921 32581 38967 32619
rect 38921 32547 38927 32581
rect 38961 32547 38967 32581
rect 38921 32509 38967 32547
rect 38921 32475 38927 32509
rect 38961 32475 38967 32509
rect 38921 32437 38967 32475
rect 38921 32403 38927 32437
rect 38961 32403 38967 32437
rect 38921 32387 38967 32403
rect 39379 33661 39425 33677
rect 39379 33627 39385 33661
rect 39419 33627 39425 33661
rect 39379 33589 39425 33627
rect 39379 33555 39385 33589
rect 39419 33555 39425 33589
rect 39379 33517 39425 33555
rect 39379 33483 39385 33517
rect 39419 33483 39425 33517
rect 39379 33445 39425 33483
rect 39379 33411 39385 33445
rect 39419 33411 39425 33445
rect 39379 33373 39425 33411
rect 39379 33339 39385 33373
rect 39419 33339 39425 33373
rect 39379 33301 39425 33339
rect 39379 33267 39385 33301
rect 39419 33267 39425 33301
rect 39379 33229 39425 33267
rect 39379 33195 39385 33229
rect 39419 33195 39425 33229
rect 39379 33157 39425 33195
rect 39379 33123 39385 33157
rect 39419 33123 39425 33157
rect 39379 33085 39425 33123
rect 39379 33051 39385 33085
rect 39419 33051 39425 33085
rect 39379 33013 39425 33051
rect 39379 32979 39385 33013
rect 39419 32979 39425 33013
rect 39379 32941 39425 32979
rect 39379 32907 39385 32941
rect 39419 32907 39425 32941
rect 39379 32869 39425 32907
rect 39379 32835 39385 32869
rect 39419 32835 39425 32869
rect 39379 32797 39425 32835
rect 39379 32763 39385 32797
rect 39419 32763 39425 32797
rect 39379 32725 39425 32763
rect 39379 32691 39385 32725
rect 39419 32691 39425 32725
rect 39379 32653 39425 32691
rect 39379 32619 39385 32653
rect 39419 32619 39425 32653
rect 39379 32581 39425 32619
rect 39379 32547 39385 32581
rect 39419 32547 39425 32581
rect 39379 32509 39425 32547
rect 39379 32475 39385 32509
rect 39419 32475 39425 32509
rect 39379 32437 39425 32475
rect 39379 32403 39385 32437
rect 39419 32403 39425 32437
rect 39379 32387 39425 32403
rect 39837 33661 39883 33677
rect 39837 33627 39843 33661
rect 39877 33627 39883 33661
rect 39837 33589 39883 33627
rect 39837 33555 39843 33589
rect 39877 33555 39883 33589
rect 39837 33517 39883 33555
rect 39837 33483 39843 33517
rect 39877 33483 39883 33517
rect 39837 33445 39883 33483
rect 39837 33411 39843 33445
rect 39877 33411 39883 33445
rect 39837 33373 39883 33411
rect 39837 33339 39843 33373
rect 39877 33339 39883 33373
rect 39837 33301 39883 33339
rect 39837 33267 39843 33301
rect 39877 33267 39883 33301
rect 39837 33229 39883 33267
rect 39837 33195 39843 33229
rect 39877 33195 39883 33229
rect 39837 33157 39883 33195
rect 39837 33123 39843 33157
rect 39877 33123 39883 33157
rect 39837 33085 39883 33123
rect 39837 33051 39843 33085
rect 39877 33051 39883 33085
rect 39837 33013 39883 33051
rect 39837 32979 39843 33013
rect 39877 32979 39883 33013
rect 39837 32941 39883 32979
rect 39837 32907 39843 32941
rect 39877 32907 39883 32941
rect 39837 32869 39883 32907
rect 39837 32835 39843 32869
rect 39877 32835 39883 32869
rect 39837 32797 39883 32835
rect 39837 32763 39843 32797
rect 39877 32763 39883 32797
rect 39837 32725 39883 32763
rect 39837 32691 39843 32725
rect 39877 32691 39883 32725
rect 39837 32653 39883 32691
rect 39837 32619 39843 32653
rect 39877 32619 39883 32653
rect 39837 32581 39883 32619
rect 39837 32547 39843 32581
rect 39877 32547 39883 32581
rect 39837 32509 39883 32547
rect 39837 32475 39843 32509
rect 39877 32475 39883 32509
rect 39837 32437 39883 32475
rect 39837 32403 39843 32437
rect 39877 32416 39883 32437
rect 40295 33661 40341 33677
rect 40295 33627 40301 33661
rect 40335 33627 40341 33661
rect 40295 33589 40341 33627
rect 40295 33555 40301 33589
rect 40335 33555 40341 33589
rect 40295 33517 40341 33555
rect 40295 33483 40301 33517
rect 40335 33483 40341 33517
rect 40295 33445 40341 33483
rect 40295 33411 40301 33445
rect 40335 33411 40341 33445
rect 40295 33373 40341 33411
rect 40295 33339 40301 33373
rect 40335 33339 40341 33373
rect 40295 33301 40341 33339
rect 40295 33267 40301 33301
rect 40335 33267 40341 33301
rect 40295 33229 40341 33267
rect 40295 33195 40301 33229
rect 40335 33195 40341 33229
rect 40295 33157 40341 33195
rect 40295 33123 40301 33157
rect 40335 33123 40341 33157
rect 40295 33085 40341 33123
rect 40295 33051 40301 33085
rect 40335 33051 40341 33085
rect 40295 33013 40341 33051
rect 40295 32979 40301 33013
rect 40335 32979 40341 33013
rect 40295 32941 40341 32979
rect 40295 32907 40301 32941
rect 40335 32907 40341 32941
rect 40295 32869 40341 32907
rect 40295 32835 40301 32869
rect 40335 32835 40341 32869
rect 40295 32797 40341 32835
rect 40295 32763 40301 32797
rect 40335 32763 40341 32797
rect 40295 32725 40341 32763
rect 40295 32691 40301 32725
rect 40335 32691 40341 32725
rect 40295 32653 40341 32691
rect 40295 32619 40301 32653
rect 40335 32619 40341 32653
rect 40295 32581 40341 32619
rect 40295 32547 40301 32581
rect 40335 32547 40341 32581
rect 40295 32509 40341 32547
rect 40295 32475 40301 32509
rect 40335 32475 40341 32509
rect 40295 32437 40341 32475
rect 40034 32416 40040 32428
rect 39877 32403 40040 32416
rect 39837 32388 40040 32403
rect 39837 32387 39883 32388
rect 40034 32376 40040 32388
rect 40092 32376 40098 32428
rect 40295 32403 40301 32437
rect 40335 32403 40341 32437
rect 40295 32387 40341 32403
rect 40753 33661 40799 33677
rect 40753 33627 40759 33661
rect 40793 33627 40799 33661
rect 40753 33589 40799 33627
rect 40753 33555 40759 33589
rect 40793 33555 40799 33589
rect 40753 33517 40799 33555
rect 40753 33483 40759 33517
rect 40793 33483 40799 33517
rect 40753 33445 40799 33483
rect 40753 33411 40759 33445
rect 40793 33411 40799 33445
rect 40753 33373 40799 33411
rect 40753 33339 40759 33373
rect 40793 33339 40799 33373
rect 40753 33301 40799 33339
rect 40753 33267 40759 33301
rect 40793 33267 40799 33301
rect 40753 33229 40799 33267
rect 40753 33195 40759 33229
rect 40793 33195 40799 33229
rect 40753 33157 40799 33195
rect 40753 33123 40759 33157
rect 40793 33123 40799 33157
rect 40753 33085 40799 33123
rect 40753 33051 40759 33085
rect 40793 33051 40799 33085
rect 40753 33013 40799 33051
rect 40753 32979 40759 33013
rect 40793 32979 40799 33013
rect 40753 32941 40799 32979
rect 40753 32907 40759 32941
rect 40793 32907 40799 32941
rect 40753 32869 40799 32907
rect 40753 32835 40759 32869
rect 40793 32835 40799 32869
rect 40753 32797 40799 32835
rect 40753 32763 40759 32797
rect 40793 32763 40799 32797
rect 40753 32725 40799 32763
rect 40753 32691 40759 32725
rect 40793 32691 40799 32725
rect 40753 32653 40799 32691
rect 40753 32619 40759 32653
rect 40793 32619 40799 32653
rect 40753 32581 40799 32619
rect 40753 32547 40759 32581
rect 40793 32547 40799 32581
rect 40753 32509 40799 32547
rect 40753 32475 40759 32509
rect 40793 32475 40799 32509
rect 40753 32437 40799 32475
rect 40753 32403 40759 32437
rect 40793 32403 40799 32437
rect 40753 32387 40799 32403
rect 41211 33661 41257 33677
rect 41211 33627 41217 33661
rect 41251 33627 41257 33661
rect 41211 33589 41257 33627
rect 41211 33555 41217 33589
rect 41251 33555 41257 33589
rect 41211 33517 41257 33555
rect 41211 33483 41217 33517
rect 41251 33483 41257 33517
rect 41211 33445 41257 33483
rect 41211 33411 41217 33445
rect 41251 33411 41257 33445
rect 41211 33373 41257 33411
rect 41211 33339 41217 33373
rect 41251 33339 41257 33373
rect 41211 33301 41257 33339
rect 41211 33267 41217 33301
rect 41251 33267 41257 33301
rect 41211 33229 41257 33267
rect 41211 33195 41217 33229
rect 41251 33195 41257 33229
rect 41211 33157 41257 33195
rect 41211 33123 41217 33157
rect 41251 33123 41257 33157
rect 41211 33085 41257 33123
rect 41211 33051 41217 33085
rect 41251 33051 41257 33085
rect 41211 33013 41257 33051
rect 41211 32979 41217 33013
rect 41251 32979 41257 33013
rect 41211 32941 41257 32979
rect 41211 32907 41217 32941
rect 41251 32907 41257 32941
rect 41211 32869 41257 32907
rect 41211 32835 41217 32869
rect 41251 32835 41257 32869
rect 41211 32797 41257 32835
rect 41211 32763 41217 32797
rect 41251 32763 41257 32797
rect 41211 32725 41257 32763
rect 41211 32691 41217 32725
rect 41251 32691 41257 32725
rect 41211 32653 41257 32691
rect 41211 32619 41217 32653
rect 41251 32619 41257 32653
rect 41211 32581 41257 32619
rect 41211 32547 41217 32581
rect 41251 32547 41257 32581
rect 41211 32509 41257 32547
rect 41211 32475 41217 32509
rect 41251 32475 41257 32509
rect 41211 32437 41257 32475
rect 41211 32403 41217 32437
rect 41251 32403 41257 32437
rect 41211 32387 41257 32403
rect 41669 33661 41715 33677
rect 41669 33627 41675 33661
rect 41709 33627 41715 33661
rect 41669 33589 41715 33627
rect 41669 33555 41675 33589
rect 41709 33555 41715 33589
rect 41669 33517 41715 33555
rect 41669 33483 41675 33517
rect 41709 33483 41715 33517
rect 41669 33445 41715 33483
rect 41669 33411 41675 33445
rect 41709 33411 41715 33445
rect 41669 33373 41715 33411
rect 41669 33339 41675 33373
rect 41709 33339 41715 33373
rect 41669 33301 41715 33339
rect 41669 33267 41675 33301
rect 41709 33267 41715 33301
rect 41669 33229 41715 33267
rect 41669 33195 41675 33229
rect 41709 33195 41715 33229
rect 41669 33157 41715 33195
rect 41669 33123 41675 33157
rect 41709 33123 41715 33157
rect 41669 33085 41715 33123
rect 41669 33051 41675 33085
rect 41709 33051 41715 33085
rect 41669 33013 41715 33051
rect 41669 32979 41675 33013
rect 41709 32979 41715 33013
rect 41669 32941 41715 32979
rect 41669 32907 41675 32941
rect 41709 32907 41715 32941
rect 41669 32869 41715 32907
rect 41669 32835 41675 32869
rect 41709 32835 41715 32869
rect 41669 32797 41715 32835
rect 41669 32763 41675 32797
rect 41709 32763 41715 32797
rect 41669 32725 41715 32763
rect 41669 32691 41675 32725
rect 41709 32691 41715 32725
rect 41669 32653 41715 32691
rect 41669 32619 41675 32653
rect 41709 32619 41715 32653
rect 41669 32581 41715 32619
rect 41669 32547 41675 32581
rect 41709 32547 41715 32581
rect 41669 32509 41715 32547
rect 41669 32475 41675 32509
rect 41709 32475 41715 32509
rect 41669 32437 41715 32475
rect 41669 32403 41675 32437
rect 41709 32403 41715 32437
rect 41669 32387 41715 32403
rect 26878 32280 26884 32292
rect 26823 32252 26884 32280
rect 26878 32240 26884 32252
rect 26936 32240 26942 32292
rect 14182 32172 14188 32224
rect 14240 32172 14246 32224
rect 14185 32147 14197 32172
rect 14231 32147 14243 32172
rect 14185 32141 14243 32147
rect 900 32090 47736 32092
rect 900 31974 922 32090
rect 2510 32049 46126 32090
rect 2510 32015 6787 32049
rect 6821 32015 7187 32049
rect 7221 32015 7587 32049
rect 7621 32015 7987 32049
rect 8021 32015 8387 32049
rect 8421 32015 8787 32049
rect 8821 32015 9187 32049
rect 9221 32015 9587 32049
rect 9621 32015 9987 32049
rect 10021 32015 10387 32049
rect 10421 32015 10787 32049
rect 10821 32015 11187 32049
rect 11221 32015 11587 32049
rect 11621 32015 11987 32049
rect 12021 32015 12387 32049
rect 12421 32015 12787 32049
rect 12821 32015 13187 32049
rect 13221 32015 13587 32049
rect 13621 32015 14331 32049
rect 14365 32015 14731 32049
rect 14765 32015 15131 32049
rect 15165 32015 15531 32049
rect 15565 32015 15931 32049
rect 15965 32015 16331 32049
rect 16365 32015 16731 32049
rect 16765 32015 17131 32049
rect 17165 32015 17531 32049
rect 17565 32015 17931 32049
rect 17965 32015 18331 32049
rect 18365 32015 18731 32049
rect 18765 32015 19131 32049
rect 19165 32015 19531 32049
rect 19565 32015 19931 32049
rect 19965 32015 20331 32049
rect 20365 32015 20731 32049
rect 20765 32015 21131 32049
rect 21165 32015 21531 32049
rect 21565 32015 21931 32049
rect 21965 32015 22331 32049
rect 22365 32015 22731 32049
rect 22765 32015 23131 32049
rect 23165 32015 23531 32049
rect 23565 32015 23931 32049
rect 23965 32015 24331 32049
rect 24365 32015 24731 32049
rect 24765 32015 25131 32049
rect 25165 32015 25531 32049
rect 25565 32015 25931 32049
rect 25965 32015 26331 32049
rect 26365 32015 26731 32049
rect 26765 32015 27131 32049
rect 27165 32015 27531 32049
rect 27565 32015 27931 32049
rect 27965 32015 28331 32049
rect 28365 32015 28731 32049
rect 28765 32015 29131 32049
rect 29165 32015 29531 32049
rect 29565 32015 29931 32049
rect 29965 32015 30331 32049
rect 30365 32015 30731 32049
rect 30765 32015 31131 32049
rect 31165 32015 31531 32049
rect 31565 32015 31931 32049
rect 31965 32015 32331 32049
rect 32365 32015 32731 32049
rect 32765 32015 33131 32049
rect 33165 32015 33531 32049
rect 33565 32015 33931 32049
rect 33965 32015 34331 32049
rect 34365 32015 34731 32049
rect 34765 32015 35131 32049
rect 35165 32015 35531 32049
rect 35565 32015 35931 32049
rect 35965 32015 36331 32049
rect 36365 32015 36731 32049
rect 36765 32015 37131 32049
rect 37165 32015 37531 32049
rect 37565 32015 37931 32049
rect 37965 32015 38331 32049
rect 38365 32015 38731 32049
rect 38765 32015 39131 32049
rect 39165 32015 39531 32049
rect 39565 32015 39931 32049
rect 39965 32015 40331 32049
rect 40365 32015 40731 32049
rect 40765 32015 41131 32049
rect 41165 32015 41531 32049
rect 41565 32015 46126 32049
rect 2510 31974 46126 32015
rect 47714 31974 47736 32090
rect 900 31972 47736 31974
rect 3348 30210 45288 30212
rect 3348 30094 3370 30210
rect 4958 30169 43678 30210
rect 4958 30135 6197 30169
rect 6231 30135 6597 30169
rect 6631 30135 6997 30169
rect 7031 30135 7397 30169
rect 7431 30135 7797 30169
rect 7831 30135 8197 30169
rect 8231 30135 8597 30169
rect 8631 30135 8997 30169
rect 9031 30135 9397 30169
rect 9431 30135 9797 30169
rect 9831 30135 10197 30169
rect 10231 30135 10597 30169
rect 10631 30135 10997 30169
rect 11031 30135 11397 30169
rect 11431 30135 11797 30169
rect 11831 30135 12197 30169
rect 12231 30135 12597 30169
rect 12631 30135 12997 30169
rect 13031 30135 13397 30169
rect 13431 30135 13797 30169
rect 13831 30135 14197 30169
rect 14231 30135 14597 30169
rect 14631 30135 14997 30169
rect 15031 30135 15397 30169
rect 15431 30135 15797 30169
rect 15831 30135 16197 30169
rect 16231 30135 16597 30169
rect 16631 30135 16997 30169
rect 17031 30135 17397 30169
rect 17431 30135 17797 30169
rect 17831 30135 18197 30169
rect 18231 30135 18597 30169
rect 18631 30135 18997 30169
rect 19031 30135 19397 30169
rect 19431 30135 19797 30169
rect 19831 30135 20197 30169
rect 20231 30135 20597 30169
rect 20631 30135 20997 30169
rect 21031 30135 21397 30169
rect 21431 30135 21797 30169
rect 21831 30135 22197 30169
rect 22231 30135 22597 30169
rect 22631 30135 22997 30169
rect 23031 30135 23397 30169
rect 23431 30135 23797 30169
rect 23831 30135 24197 30169
rect 24231 30135 24597 30169
rect 24631 30135 24997 30169
rect 25031 30135 25397 30169
rect 25431 30135 25797 30169
rect 25831 30135 26197 30169
rect 26231 30135 26597 30169
rect 26631 30135 26997 30169
rect 27031 30135 27397 30169
rect 27431 30135 27797 30169
rect 27831 30135 28197 30169
rect 28231 30135 28597 30169
rect 28631 30135 28997 30169
rect 29031 30135 29397 30169
rect 29431 30135 29797 30169
rect 29831 30135 30197 30169
rect 30231 30135 30597 30169
rect 30631 30135 30997 30169
rect 31031 30135 31397 30169
rect 31431 30135 31797 30169
rect 31831 30135 32197 30169
rect 32231 30135 32597 30169
rect 32631 30135 32997 30169
rect 33031 30135 33397 30169
rect 33431 30135 34225 30169
rect 34259 30135 34625 30169
rect 34659 30135 35025 30169
rect 35059 30135 35425 30169
rect 35459 30135 35825 30169
rect 35859 30135 36225 30169
rect 36259 30135 36625 30169
rect 36659 30135 37577 30169
rect 37611 30135 37777 30169
rect 37811 30135 37977 30169
rect 38011 30135 38177 30169
rect 38211 30135 38377 30169
rect 38411 30135 38577 30169
rect 38611 30135 38777 30169
rect 38811 30135 38977 30169
rect 39011 30135 39177 30169
rect 39211 30135 39377 30169
rect 39411 30135 39577 30169
rect 39611 30135 40321 30169
rect 40355 30135 40521 30169
rect 40555 30135 40721 30169
rect 40755 30135 40921 30169
rect 40955 30135 41121 30169
rect 41155 30135 41321 30169
rect 41355 30135 41521 30169
rect 41555 30135 41721 30169
rect 41755 30135 41921 30169
rect 41955 30135 42121 30169
rect 42155 30135 42321 30169
rect 42355 30135 43678 30169
rect 4958 30094 43678 30135
rect 45266 30094 45288 30210
rect 3348 30092 45288 30094
rect 17512 29917 17540 30092
rect 6055 29901 6101 29917
rect 6055 29867 6061 29901
rect 6095 29867 6101 29901
rect 6055 29829 6101 29867
rect 6055 29795 6061 29829
rect 6095 29795 6101 29829
rect 6055 29757 6101 29795
rect 6055 29723 6061 29757
rect 6095 29723 6101 29757
rect 6055 29685 6101 29723
rect 6055 29651 6061 29685
rect 6095 29651 6101 29685
rect 6055 29613 6101 29651
rect 6055 29579 6061 29613
rect 6095 29579 6101 29613
rect 6055 29541 6101 29579
rect 6055 29507 6061 29541
rect 6095 29507 6101 29541
rect 6055 29469 6101 29507
rect 6055 29435 6061 29469
rect 6095 29435 6101 29469
rect 6055 29397 6101 29435
rect 6055 29363 6061 29397
rect 6095 29363 6101 29397
rect 6055 29325 6101 29363
rect 6055 29291 6061 29325
rect 6095 29291 6101 29325
rect 6055 29253 6101 29291
rect 6055 29219 6061 29253
rect 6095 29219 6101 29253
rect 6055 29181 6101 29219
rect 6055 29147 6061 29181
rect 6095 29147 6101 29181
rect 6055 29109 6101 29147
rect 6055 29075 6061 29109
rect 6095 29075 6101 29109
rect 6055 29037 6101 29075
rect 6055 29003 6061 29037
rect 6095 29003 6101 29037
rect 6055 28965 6101 29003
rect 6055 28931 6061 28965
rect 6095 28931 6101 28965
rect 6055 28893 6101 28931
rect 6055 28859 6061 28893
rect 6095 28859 6101 28893
rect 6055 28821 6101 28859
rect 6055 28787 6061 28821
rect 6095 28787 6101 28821
rect 6055 28749 6101 28787
rect 6055 28715 6061 28749
rect 6095 28715 6101 28749
rect 6055 28677 6101 28715
rect 6055 28643 6061 28677
rect 6095 28643 6101 28677
rect 6055 28627 6101 28643
rect 6513 29901 6559 29917
rect 6513 29867 6519 29901
rect 6553 29867 6559 29901
rect 6513 29829 6559 29867
rect 6513 29795 6519 29829
rect 6553 29795 6559 29829
rect 6513 29757 6559 29795
rect 6513 29723 6519 29757
rect 6553 29723 6559 29757
rect 6513 29685 6559 29723
rect 6513 29651 6519 29685
rect 6553 29651 6559 29685
rect 6513 29613 6559 29651
rect 6513 29579 6519 29613
rect 6553 29579 6559 29613
rect 6513 29541 6559 29579
rect 6513 29507 6519 29541
rect 6553 29507 6559 29541
rect 6513 29469 6559 29507
rect 6513 29435 6519 29469
rect 6553 29435 6559 29469
rect 6513 29397 6559 29435
rect 6513 29363 6519 29397
rect 6553 29363 6559 29397
rect 6513 29325 6559 29363
rect 6513 29291 6519 29325
rect 6553 29291 6559 29325
rect 6513 29253 6559 29291
rect 6513 29219 6519 29253
rect 6553 29219 6559 29253
rect 6513 29181 6559 29219
rect 6513 29147 6519 29181
rect 6553 29147 6559 29181
rect 6513 29109 6559 29147
rect 6513 29075 6519 29109
rect 6553 29075 6559 29109
rect 6513 29037 6559 29075
rect 6513 29003 6519 29037
rect 6553 29003 6559 29037
rect 6513 28965 6559 29003
rect 6513 28931 6519 28965
rect 6553 28931 6559 28965
rect 6513 28893 6559 28931
rect 6513 28859 6519 28893
rect 6553 28859 6559 28893
rect 6513 28821 6559 28859
rect 6513 28787 6519 28821
rect 6553 28787 6559 28821
rect 6513 28749 6559 28787
rect 6513 28715 6519 28749
rect 6553 28715 6559 28749
rect 6513 28677 6559 28715
rect 6513 28643 6519 28677
rect 6553 28643 6559 28677
rect 6513 28627 6559 28643
rect 6971 29901 7017 29917
rect 6971 29867 6977 29901
rect 7011 29867 7017 29901
rect 6971 29829 7017 29867
rect 6971 29795 6977 29829
rect 7011 29795 7017 29829
rect 6971 29757 7017 29795
rect 6971 29723 6977 29757
rect 7011 29723 7017 29757
rect 6971 29685 7017 29723
rect 6971 29651 6977 29685
rect 7011 29651 7017 29685
rect 6971 29613 7017 29651
rect 6971 29579 6977 29613
rect 7011 29579 7017 29613
rect 6971 29541 7017 29579
rect 6971 29507 6977 29541
rect 7011 29507 7017 29541
rect 6971 29469 7017 29507
rect 6971 29435 6977 29469
rect 7011 29435 7017 29469
rect 6971 29397 7017 29435
rect 6971 29363 6977 29397
rect 7011 29363 7017 29397
rect 6971 29325 7017 29363
rect 6971 29291 6977 29325
rect 7011 29291 7017 29325
rect 6971 29253 7017 29291
rect 6971 29219 6977 29253
rect 7011 29219 7017 29253
rect 6971 29181 7017 29219
rect 6971 29147 6977 29181
rect 7011 29147 7017 29181
rect 6971 29109 7017 29147
rect 6971 29075 6977 29109
rect 7011 29075 7017 29109
rect 6971 29037 7017 29075
rect 6971 29003 6977 29037
rect 7011 29003 7017 29037
rect 6971 28965 7017 29003
rect 6971 28931 6977 28965
rect 7011 28931 7017 28965
rect 6971 28893 7017 28931
rect 6971 28859 6977 28893
rect 7011 28859 7017 28893
rect 6971 28821 7017 28859
rect 6971 28787 6977 28821
rect 7011 28787 7017 28821
rect 6971 28749 7017 28787
rect 6971 28715 6977 28749
rect 7011 28715 7017 28749
rect 6971 28677 7017 28715
rect 6971 28643 6977 28677
rect 7011 28643 7017 28677
rect 6971 28627 7017 28643
rect 7429 29901 7475 29917
rect 7429 29867 7435 29901
rect 7469 29867 7475 29901
rect 7429 29829 7475 29867
rect 7429 29795 7435 29829
rect 7469 29795 7475 29829
rect 7429 29757 7475 29795
rect 7429 29723 7435 29757
rect 7469 29723 7475 29757
rect 7429 29685 7475 29723
rect 7429 29651 7435 29685
rect 7469 29651 7475 29685
rect 7429 29613 7475 29651
rect 7429 29579 7435 29613
rect 7469 29579 7475 29613
rect 7429 29541 7475 29579
rect 7429 29507 7435 29541
rect 7469 29507 7475 29541
rect 7429 29469 7475 29507
rect 7429 29435 7435 29469
rect 7469 29435 7475 29469
rect 7429 29397 7475 29435
rect 7429 29363 7435 29397
rect 7469 29363 7475 29397
rect 7429 29325 7475 29363
rect 7429 29291 7435 29325
rect 7469 29291 7475 29325
rect 7429 29253 7475 29291
rect 7429 29219 7435 29253
rect 7469 29219 7475 29253
rect 7429 29181 7475 29219
rect 7429 29147 7435 29181
rect 7469 29147 7475 29181
rect 7429 29109 7475 29147
rect 7429 29075 7435 29109
rect 7469 29075 7475 29109
rect 7429 29037 7475 29075
rect 7429 29003 7435 29037
rect 7469 29003 7475 29037
rect 7429 28965 7475 29003
rect 7429 28931 7435 28965
rect 7469 28931 7475 28965
rect 7429 28893 7475 28931
rect 7429 28859 7435 28893
rect 7469 28859 7475 28893
rect 7429 28821 7475 28859
rect 7429 28787 7435 28821
rect 7469 28787 7475 28821
rect 7429 28749 7475 28787
rect 7429 28715 7435 28749
rect 7469 28715 7475 28749
rect 7429 28677 7475 28715
rect 7429 28643 7435 28677
rect 7469 28643 7475 28677
rect 7429 28627 7475 28643
rect 7887 29901 7933 29917
rect 7887 29867 7893 29901
rect 7927 29867 7933 29901
rect 7887 29829 7933 29867
rect 7887 29795 7893 29829
rect 7927 29795 7933 29829
rect 7887 29757 7933 29795
rect 7887 29723 7893 29757
rect 7927 29723 7933 29757
rect 7887 29685 7933 29723
rect 7887 29651 7893 29685
rect 7927 29651 7933 29685
rect 7887 29613 7933 29651
rect 7887 29579 7893 29613
rect 7927 29579 7933 29613
rect 7887 29541 7933 29579
rect 7887 29507 7893 29541
rect 7927 29507 7933 29541
rect 7887 29469 7933 29507
rect 7887 29435 7893 29469
rect 7927 29435 7933 29469
rect 7887 29397 7933 29435
rect 7887 29363 7893 29397
rect 7927 29363 7933 29397
rect 7887 29325 7933 29363
rect 7887 29291 7893 29325
rect 7927 29291 7933 29325
rect 7887 29253 7933 29291
rect 7887 29219 7893 29253
rect 7927 29219 7933 29253
rect 7887 29181 7933 29219
rect 7887 29147 7893 29181
rect 7927 29147 7933 29181
rect 7887 29109 7933 29147
rect 7887 29075 7893 29109
rect 7927 29075 7933 29109
rect 7887 29037 7933 29075
rect 7887 29003 7893 29037
rect 7927 29003 7933 29037
rect 7887 28965 7933 29003
rect 7887 28931 7893 28965
rect 7927 28931 7933 28965
rect 7887 28893 7933 28931
rect 7887 28859 7893 28893
rect 7927 28859 7933 28893
rect 7887 28821 7933 28859
rect 7887 28787 7893 28821
rect 7927 28787 7933 28821
rect 7887 28749 7933 28787
rect 7887 28715 7893 28749
rect 7927 28715 7933 28749
rect 7887 28677 7933 28715
rect 7887 28643 7893 28677
rect 7927 28643 7933 28677
rect 7887 28627 7933 28643
rect 8345 29901 8391 29917
rect 8345 29867 8351 29901
rect 8385 29867 8391 29901
rect 8345 29829 8391 29867
rect 8345 29795 8351 29829
rect 8385 29795 8391 29829
rect 8345 29757 8391 29795
rect 8345 29723 8351 29757
rect 8385 29723 8391 29757
rect 8345 29685 8391 29723
rect 8345 29651 8351 29685
rect 8385 29651 8391 29685
rect 8345 29613 8391 29651
rect 8345 29579 8351 29613
rect 8385 29579 8391 29613
rect 8345 29541 8391 29579
rect 8345 29507 8351 29541
rect 8385 29507 8391 29541
rect 8345 29469 8391 29507
rect 8345 29435 8351 29469
rect 8385 29435 8391 29469
rect 8345 29397 8391 29435
rect 8345 29363 8351 29397
rect 8385 29363 8391 29397
rect 8345 29325 8391 29363
rect 8345 29291 8351 29325
rect 8385 29291 8391 29325
rect 8345 29253 8391 29291
rect 8345 29219 8351 29253
rect 8385 29219 8391 29253
rect 8345 29181 8391 29219
rect 8345 29147 8351 29181
rect 8385 29147 8391 29181
rect 8345 29109 8391 29147
rect 8345 29075 8351 29109
rect 8385 29075 8391 29109
rect 8345 29037 8391 29075
rect 8345 29003 8351 29037
rect 8385 29003 8391 29037
rect 8345 28965 8391 29003
rect 8345 28931 8351 28965
rect 8385 28931 8391 28965
rect 8345 28893 8391 28931
rect 8345 28859 8351 28893
rect 8385 28859 8391 28893
rect 8345 28821 8391 28859
rect 8345 28787 8351 28821
rect 8385 28787 8391 28821
rect 8345 28749 8391 28787
rect 8345 28715 8351 28749
rect 8385 28715 8391 28749
rect 8345 28677 8391 28715
rect 8345 28643 8351 28677
rect 8385 28643 8391 28677
rect 8345 28627 8391 28643
rect 8803 29901 8849 29917
rect 8803 29867 8809 29901
rect 8843 29867 8849 29901
rect 8803 29829 8849 29867
rect 8803 29795 8809 29829
rect 8843 29795 8849 29829
rect 8803 29757 8849 29795
rect 8803 29723 8809 29757
rect 8843 29723 8849 29757
rect 8803 29685 8849 29723
rect 8803 29651 8809 29685
rect 8843 29651 8849 29685
rect 8803 29613 8849 29651
rect 8803 29579 8809 29613
rect 8843 29579 8849 29613
rect 8803 29541 8849 29579
rect 8803 29507 8809 29541
rect 8843 29507 8849 29541
rect 8803 29469 8849 29507
rect 8803 29435 8809 29469
rect 8843 29435 8849 29469
rect 8803 29397 8849 29435
rect 8803 29363 8809 29397
rect 8843 29363 8849 29397
rect 8803 29325 8849 29363
rect 8803 29291 8809 29325
rect 8843 29291 8849 29325
rect 8803 29253 8849 29291
rect 8803 29219 8809 29253
rect 8843 29219 8849 29253
rect 8803 29181 8849 29219
rect 8803 29147 8809 29181
rect 8843 29147 8849 29181
rect 8803 29109 8849 29147
rect 8803 29075 8809 29109
rect 8843 29075 8849 29109
rect 8803 29037 8849 29075
rect 8803 29003 8809 29037
rect 8843 29003 8849 29037
rect 8803 28965 8849 29003
rect 8803 28931 8809 28965
rect 8843 28931 8849 28965
rect 8803 28893 8849 28931
rect 8803 28859 8809 28893
rect 8843 28859 8849 28893
rect 8803 28821 8849 28859
rect 8803 28787 8809 28821
rect 8843 28787 8849 28821
rect 8803 28749 8849 28787
rect 8803 28715 8809 28749
rect 8843 28715 8849 28749
rect 8803 28677 8849 28715
rect 8803 28643 8809 28677
rect 8843 28643 8849 28677
rect 8803 28627 8849 28643
rect 9261 29901 9307 29917
rect 9261 29867 9267 29901
rect 9301 29867 9307 29901
rect 9261 29829 9307 29867
rect 9261 29795 9267 29829
rect 9301 29795 9307 29829
rect 9261 29757 9307 29795
rect 9261 29723 9267 29757
rect 9301 29723 9307 29757
rect 9261 29685 9307 29723
rect 9261 29651 9267 29685
rect 9301 29651 9307 29685
rect 9261 29613 9307 29651
rect 9261 29579 9267 29613
rect 9301 29579 9307 29613
rect 9261 29541 9307 29579
rect 9261 29507 9267 29541
rect 9301 29507 9307 29541
rect 9261 29469 9307 29507
rect 9261 29435 9267 29469
rect 9301 29435 9307 29469
rect 9261 29397 9307 29435
rect 9261 29363 9267 29397
rect 9301 29363 9307 29397
rect 9261 29325 9307 29363
rect 9261 29291 9267 29325
rect 9301 29291 9307 29325
rect 9261 29253 9307 29291
rect 9261 29219 9267 29253
rect 9301 29219 9307 29253
rect 9261 29181 9307 29219
rect 9261 29147 9267 29181
rect 9301 29147 9307 29181
rect 9261 29109 9307 29147
rect 9261 29075 9267 29109
rect 9301 29075 9307 29109
rect 9261 29037 9307 29075
rect 9261 29003 9267 29037
rect 9301 29003 9307 29037
rect 9261 28965 9307 29003
rect 9261 28931 9267 28965
rect 9301 28931 9307 28965
rect 9261 28893 9307 28931
rect 9261 28859 9267 28893
rect 9301 28859 9307 28893
rect 9261 28821 9307 28859
rect 9261 28787 9267 28821
rect 9301 28787 9307 28821
rect 9261 28749 9307 28787
rect 9261 28715 9267 28749
rect 9301 28715 9307 28749
rect 9261 28677 9307 28715
rect 9261 28643 9267 28677
rect 9301 28643 9307 28677
rect 9261 28627 9307 28643
rect 9719 29901 9765 29917
rect 9719 29867 9725 29901
rect 9759 29867 9765 29901
rect 9719 29829 9765 29867
rect 9719 29795 9725 29829
rect 9759 29795 9765 29829
rect 9719 29757 9765 29795
rect 9719 29723 9725 29757
rect 9759 29723 9765 29757
rect 9719 29685 9765 29723
rect 9719 29651 9725 29685
rect 9759 29651 9765 29685
rect 9719 29613 9765 29651
rect 9719 29579 9725 29613
rect 9759 29579 9765 29613
rect 9719 29541 9765 29579
rect 9719 29507 9725 29541
rect 9759 29507 9765 29541
rect 9719 29469 9765 29507
rect 9719 29435 9725 29469
rect 9759 29435 9765 29469
rect 9719 29397 9765 29435
rect 9719 29363 9725 29397
rect 9759 29363 9765 29397
rect 9719 29325 9765 29363
rect 9719 29291 9725 29325
rect 9759 29291 9765 29325
rect 9719 29253 9765 29291
rect 9719 29219 9725 29253
rect 9759 29219 9765 29253
rect 9719 29181 9765 29219
rect 9719 29147 9725 29181
rect 9759 29147 9765 29181
rect 9719 29109 9765 29147
rect 9719 29075 9725 29109
rect 9759 29075 9765 29109
rect 9719 29037 9765 29075
rect 9719 29003 9725 29037
rect 9759 29003 9765 29037
rect 9719 28965 9765 29003
rect 9719 28931 9725 28965
rect 9759 28931 9765 28965
rect 9719 28893 9765 28931
rect 9719 28859 9725 28893
rect 9759 28859 9765 28893
rect 9719 28821 9765 28859
rect 9719 28787 9725 28821
rect 9759 28787 9765 28821
rect 9719 28749 9765 28787
rect 9719 28715 9725 28749
rect 9759 28715 9765 28749
rect 9719 28677 9765 28715
rect 9719 28643 9725 28677
rect 9759 28643 9765 28677
rect 9719 28627 9765 28643
rect 10177 29901 10223 29917
rect 10177 29867 10183 29901
rect 10217 29867 10223 29901
rect 10177 29829 10223 29867
rect 10177 29795 10183 29829
rect 10217 29795 10223 29829
rect 10177 29757 10223 29795
rect 10177 29723 10183 29757
rect 10217 29723 10223 29757
rect 10177 29685 10223 29723
rect 10177 29651 10183 29685
rect 10217 29651 10223 29685
rect 10177 29613 10223 29651
rect 10177 29579 10183 29613
rect 10217 29579 10223 29613
rect 10177 29541 10223 29579
rect 10177 29507 10183 29541
rect 10217 29507 10223 29541
rect 10177 29469 10223 29507
rect 10177 29435 10183 29469
rect 10217 29435 10223 29469
rect 10177 29397 10223 29435
rect 10177 29363 10183 29397
rect 10217 29363 10223 29397
rect 10177 29325 10223 29363
rect 10177 29291 10183 29325
rect 10217 29291 10223 29325
rect 10177 29253 10223 29291
rect 10177 29219 10183 29253
rect 10217 29219 10223 29253
rect 10177 29181 10223 29219
rect 10177 29147 10183 29181
rect 10217 29147 10223 29181
rect 10177 29109 10223 29147
rect 10177 29075 10183 29109
rect 10217 29075 10223 29109
rect 10177 29037 10223 29075
rect 10177 29003 10183 29037
rect 10217 29003 10223 29037
rect 10177 28965 10223 29003
rect 10177 28931 10183 28965
rect 10217 28931 10223 28965
rect 10177 28893 10223 28931
rect 10177 28859 10183 28893
rect 10217 28859 10223 28893
rect 10177 28821 10223 28859
rect 10177 28787 10183 28821
rect 10217 28787 10223 28821
rect 10177 28749 10223 28787
rect 10177 28715 10183 28749
rect 10217 28715 10223 28749
rect 10177 28677 10223 28715
rect 10177 28643 10183 28677
rect 10217 28643 10223 28677
rect 10177 28627 10223 28643
rect 10635 29901 10681 29917
rect 10635 29867 10641 29901
rect 10675 29867 10681 29901
rect 10635 29829 10681 29867
rect 10635 29795 10641 29829
rect 10675 29795 10681 29829
rect 10635 29757 10681 29795
rect 10635 29723 10641 29757
rect 10675 29723 10681 29757
rect 10635 29685 10681 29723
rect 10635 29651 10641 29685
rect 10675 29651 10681 29685
rect 10635 29613 10681 29651
rect 10635 29579 10641 29613
rect 10675 29579 10681 29613
rect 10635 29541 10681 29579
rect 10635 29507 10641 29541
rect 10675 29507 10681 29541
rect 10635 29469 10681 29507
rect 10635 29435 10641 29469
rect 10675 29435 10681 29469
rect 10635 29397 10681 29435
rect 10635 29363 10641 29397
rect 10675 29363 10681 29397
rect 10635 29325 10681 29363
rect 10635 29291 10641 29325
rect 10675 29291 10681 29325
rect 10635 29253 10681 29291
rect 10635 29219 10641 29253
rect 10675 29219 10681 29253
rect 10635 29181 10681 29219
rect 10635 29147 10641 29181
rect 10675 29147 10681 29181
rect 10635 29109 10681 29147
rect 10635 29075 10641 29109
rect 10675 29075 10681 29109
rect 10635 29037 10681 29075
rect 10635 29003 10641 29037
rect 10675 29003 10681 29037
rect 10635 28965 10681 29003
rect 10635 28931 10641 28965
rect 10675 28931 10681 28965
rect 10635 28893 10681 28931
rect 10635 28859 10641 28893
rect 10675 28859 10681 28893
rect 10635 28821 10681 28859
rect 10635 28787 10641 28821
rect 10675 28787 10681 28821
rect 10635 28749 10681 28787
rect 10635 28715 10641 28749
rect 10675 28715 10681 28749
rect 10635 28677 10681 28715
rect 10635 28643 10641 28677
rect 10675 28643 10681 28677
rect 10635 28627 10681 28643
rect 11093 29901 11139 29917
rect 11093 29867 11099 29901
rect 11133 29867 11139 29901
rect 11093 29829 11139 29867
rect 11093 29795 11099 29829
rect 11133 29795 11139 29829
rect 11093 29757 11139 29795
rect 11093 29723 11099 29757
rect 11133 29723 11139 29757
rect 11093 29685 11139 29723
rect 11093 29651 11099 29685
rect 11133 29651 11139 29685
rect 11093 29613 11139 29651
rect 11093 29579 11099 29613
rect 11133 29579 11139 29613
rect 11093 29541 11139 29579
rect 11093 29507 11099 29541
rect 11133 29507 11139 29541
rect 11093 29469 11139 29507
rect 11093 29435 11099 29469
rect 11133 29435 11139 29469
rect 11093 29397 11139 29435
rect 11093 29363 11099 29397
rect 11133 29363 11139 29397
rect 11093 29325 11139 29363
rect 11093 29291 11099 29325
rect 11133 29291 11139 29325
rect 11093 29253 11139 29291
rect 11093 29219 11099 29253
rect 11133 29219 11139 29253
rect 11093 29181 11139 29219
rect 11093 29147 11099 29181
rect 11133 29147 11139 29181
rect 11093 29109 11139 29147
rect 11093 29075 11099 29109
rect 11133 29075 11139 29109
rect 11093 29037 11139 29075
rect 11093 29003 11099 29037
rect 11133 29003 11139 29037
rect 11093 28965 11139 29003
rect 11093 28931 11099 28965
rect 11133 28931 11139 28965
rect 11093 28893 11139 28931
rect 11093 28859 11099 28893
rect 11133 28859 11139 28893
rect 11093 28821 11139 28859
rect 11093 28787 11099 28821
rect 11133 28787 11139 28821
rect 11093 28749 11139 28787
rect 11093 28715 11099 28749
rect 11133 28715 11139 28749
rect 11093 28677 11139 28715
rect 11093 28643 11099 28677
rect 11133 28643 11139 28677
rect 11093 28627 11139 28643
rect 11551 29901 11597 29917
rect 11551 29867 11557 29901
rect 11591 29867 11597 29901
rect 11551 29829 11597 29867
rect 11551 29795 11557 29829
rect 11591 29795 11597 29829
rect 11551 29757 11597 29795
rect 11551 29723 11557 29757
rect 11591 29723 11597 29757
rect 11551 29685 11597 29723
rect 11551 29651 11557 29685
rect 11591 29651 11597 29685
rect 11551 29613 11597 29651
rect 11551 29579 11557 29613
rect 11591 29579 11597 29613
rect 11551 29541 11597 29579
rect 11551 29507 11557 29541
rect 11591 29507 11597 29541
rect 11551 29469 11597 29507
rect 11551 29435 11557 29469
rect 11591 29435 11597 29469
rect 11551 29397 11597 29435
rect 11551 29363 11557 29397
rect 11591 29363 11597 29397
rect 11551 29325 11597 29363
rect 11551 29291 11557 29325
rect 11591 29291 11597 29325
rect 11551 29253 11597 29291
rect 11551 29219 11557 29253
rect 11591 29219 11597 29253
rect 11551 29181 11597 29219
rect 11551 29147 11557 29181
rect 11591 29147 11597 29181
rect 11551 29109 11597 29147
rect 11551 29075 11557 29109
rect 11591 29075 11597 29109
rect 11551 29037 11597 29075
rect 11551 29003 11557 29037
rect 11591 29003 11597 29037
rect 11551 28965 11597 29003
rect 11551 28931 11557 28965
rect 11591 28931 11597 28965
rect 11551 28893 11597 28931
rect 11551 28859 11557 28893
rect 11591 28859 11597 28893
rect 11551 28821 11597 28859
rect 11551 28787 11557 28821
rect 11591 28787 11597 28821
rect 11551 28749 11597 28787
rect 11551 28715 11557 28749
rect 11591 28715 11597 28749
rect 11551 28677 11597 28715
rect 11551 28643 11557 28677
rect 11591 28643 11597 28677
rect 11551 28627 11597 28643
rect 12009 29901 12055 29917
rect 12009 29867 12015 29901
rect 12049 29867 12055 29901
rect 12009 29829 12055 29867
rect 12009 29795 12015 29829
rect 12049 29795 12055 29829
rect 12009 29757 12055 29795
rect 12009 29723 12015 29757
rect 12049 29723 12055 29757
rect 12009 29685 12055 29723
rect 12009 29651 12015 29685
rect 12049 29651 12055 29685
rect 12009 29613 12055 29651
rect 12009 29579 12015 29613
rect 12049 29579 12055 29613
rect 12009 29541 12055 29579
rect 12009 29507 12015 29541
rect 12049 29507 12055 29541
rect 12009 29469 12055 29507
rect 12009 29435 12015 29469
rect 12049 29435 12055 29469
rect 12009 29397 12055 29435
rect 12009 29363 12015 29397
rect 12049 29363 12055 29397
rect 12009 29325 12055 29363
rect 12009 29291 12015 29325
rect 12049 29291 12055 29325
rect 12009 29253 12055 29291
rect 12009 29219 12015 29253
rect 12049 29219 12055 29253
rect 12009 29181 12055 29219
rect 12009 29147 12015 29181
rect 12049 29147 12055 29181
rect 12009 29109 12055 29147
rect 12009 29075 12015 29109
rect 12049 29075 12055 29109
rect 12009 29037 12055 29075
rect 12009 29003 12015 29037
rect 12049 29003 12055 29037
rect 12009 28965 12055 29003
rect 12009 28931 12015 28965
rect 12049 28931 12055 28965
rect 12009 28893 12055 28931
rect 12009 28859 12015 28893
rect 12049 28859 12055 28893
rect 12009 28821 12055 28859
rect 12009 28787 12015 28821
rect 12049 28787 12055 28821
rect 12009 28749 12055 28787
rect 12009 28715 12015 28749
rect 12049 28715 12055 28749
rect 12009 28677 12055 28715
rect 12009 28643 12015 28677
rect 12049 28643 12055 28677
rect 12009 28627 12055 28643
rect 12467 29901 12513 29917
rect 12467 29867 12473 29901
rect 12507 29867 12513 29901
rect 12467 29829 12513 29867
rect 12467 29795 12473 29829
rect 12507 29795 12513 29829
rect 12467 29757 12513 29795
rect 12467 29723 12473 29757
rect 12507 29723 12513 29757
rect 12467 29685 12513 29723
rect 12467 29651 12473 29685
rect 12507 29651 12513 29685
rect 12467 29613 12513 29651
rect 12467 29579 12473 29613
rect 12507 29579 12513 29613
rect 12467 29541 12513 29579
rect 12467 29507 12473 29541
rect 12507 29507 12513 29541
rect 12467 29469 12513 29507
rect 12467 29435 12473 29469
rect 12507 29435 12513 29469
rect 12467 29397 12513 29435
rect 12467 29363 12473 29397
rect 12507 29363 12513 29397
rect 12467 29325 12513 29363
rect 12467 29291 12473 29325
rect 12507 29291 12513 29325
rect 12467 29253 12513 29291
rect 12467 29219 12473 29253
rect 12507 29219 12513 29253
rect 12467 29181 12513 29219
rect 12467 29147 12473 29181
rect 12507 29147 12513 29181
rect 12467 29109 12513 29147
rect 12467 29075 12473 29109
rect 12507 29075 12513 29109
rect 12467 29037 12513 29075
rect 12467 29003 12473 29037
rect 12507 29003 12513 29037
rect 12467 28965 12513 29003
rect 12467 28931 12473 28965
rect 12507 28931 12513 28965
rect 12467 28893 12513 28931
rect 12467 28859 12473 28893
rect 12507 28859 12513 28893
rect 12467 28821 12513 28859
rect 12467 28787 12473 28821
rect 12507 28787 12513 28821
rect 12467 28749 12513 28787
rect 12467 28715 12473 28749
rect 12507 28715 12513 28749
rect 12467 28677 12513 28715
rect 12467 28643 12473 28677
rect 12507 28643 12513 28677
rect 12467 28627 12513 28643
rect 12925 29901 12971 29917
rect 12925 29867 12931 29901
rect 12965 29867 12971 29901
rect 12925 29829 12971 29867
rect 12925 29795 12931 29829
rect 12965 29795 12971 29829
rect 12925 29757 12971 29795
rect 12925 29723 12931 29757
rect 12965 29723 12971 29757
rect 12925 29685 12971 29723
rect 12925 29651 12931 29685
rect 12965 29651 12971 29685
rect 12925 29613 12971 29651
rect 12925 29579 12931 29613
rect 12965 29579 12971 29613
rect 12925 29541 12971 29579
rect 12925 29507 12931 29541
rect 12965 29507 12971 29541
rect 12925 29469 12971 29507
rect 12925 29435 12931 29469
rect 12965 29435 12971 29469
rect 12925 29397 12971 29435
rect 12925 29363 12931 29397
rect 12965 29363 12971 29397
rect 12925 29325 12971 29363
rect 12925 29291 12931 29325
rect 12965 29291 12971 29325
rect 12925 29253 12971 29291
rect 12925 29219 12931 29253
rect 12965 29219 12971 29253
rect 12925 29181 12971 29219
rect 12925 29147 12931 29181
rect 12965 29147 12971 29181
rect 12925 29109 12971 29147
rect 12925 29075 12931 29109
rect 12965 29075 12971 29109
rect 12925 29037 12971 29075
rect 12925 29003 12931 29037
rect 12965 29003 12971 29037
rect 12925 28965 12971 29003
rect 12925 28931 12931 28965
rect 12965 28931 12971 28965
rect 12925 28893 12971 28931
rect 12925 28859 12931 28893
rect 12965 28859 12971 28893
rect 12925 28821 12971 28859
rect 12925 28787 12931 28821
rect 12965 28787 12971 28821
rect 12925 28749 12971 28787
rect 12925 28715 12931 28749
rect 12965 28715 12971 28749
rect 12925 28677 12971 28715
rect 12925 28643 12931 28677
rect 12965 28643 12971 28677
rect 12925 28627 12971 28643
rect 13383 29901 13429 29917
rect 13383 29867 13389 29901
rect 13423 29867 13429 29901
rect 13383 29829 13429 29867
rect 13383 29795 13389 29829
rect 13423 29795 13429 29829
rect 13383 29757 13429 29795
rect 13383 29723 13389 29757
rect 13423 29723 13429 29757
rect 13383 29685 13429 29723
rect 13383 29651 13389 29685
rect 13423 29651 13429 29685
rect 13383 29613 13429 29651
rect 13383 29579 13389 29613
rect 13423 29579 13429 29613
rect 13383 29541 13429 29579
rect 13383 29507 13389 29541
rect 13423 29507 13429 29541
rect 13383 29469 13429 29507
rect 13383 29435 13389 29469
rect 13423 29435 13429 29469
rect 13383 29397 13429 29435
rect 13383 29363 13389 29397
rect 13423 29363 13429 29397
rect 13383 29325 13429 29363
rect 13383 29291 13389 29325
rect 13423 29291 13429 29325
rect 13383 29253 13429 29291
rect 13383 29219 13389 29253
rect 13423 29219 13429 29253
rect 13383 29181 13429 29219
rect 13383 29147 13389 29181
rect 13423 29147 13429 29181
rect 13383 29109 13429 29147
rect 13383 29075 13389 29109
rect 13423 29075 13429 29109
rect 13383 29037 13429 29075
rect 13383 29003 13389 29037
rect 13423 29003 13429 29037
rect 13383 28965 13429 29003
rect 13383 28931 13389 28965
rect 13423 28931 13429 28965
rect 13383 28893 13429 28931
rect 13383 28859 13389 28893
rect 13423 28859 13429 28893
rect 13383 28821 13429 28859
rect 13383 28787 13389 28821
rect 13423 28787 13429 28821
rect 13383 28749 13429 28787
rect 13383 28715 13389 28749
rect 13423 28715 13429 28749
rect 13383 28677 13429 28715
rect 13383 28643 13389 28677
rect 13423 28643 13429 28677
rect 13383 28627 13429 28643
rect 13841 29901 13887 29917
rect 13841 29867 13847 29901
rect 13881 29867 13887 29901
rect 13841 29829 13887 29867
rect 13841 29795 13847 29829
rect 13881 29795 13887 29829
rect 13841 29757 13887 29795
rect 13841 29723 13847 29757
rect 13881 29723 13887 29757
rect 13841 29685 13887 29723
rect 13841 29651 13847 29685
rect 13881 29651 13887 29685
rect 13841 29613 13887 29651
rect 13841 29579 13847 29613
rect 13881 29579 13887 29613
rect 13841 29541 13887 29579
rect 13841 29507 13847 29541
rect 13881 29507 13887 29541
rect 13841 29469 13887 29507
rect 13841 29435 13847 29469
rect 13881 29435 13887 29469
rect 13841 29397 13887 29435
rect 13841 29363 13847 29397
rect 13881 29363 13887 29397
rect 13841 29325 13887 29363
rect 13841 29291 13847 29325
rect 13881 29291 13887 29325
rect 13841 29253 13887 29291
rect 13841 29219 13847 29253
rect 13881 29219 13887 29253
rect 13841 29181 13887 29219
rect 13841 29147 13847 29181
rect 13881 29147 13887 29181
rect 13841 29109 13887 29147
rect 13841 29075 13847 29109
rect 13881 29075 13887 29109
rect 13841 29037 13887 29075
rect 13841 29003 13847 29037
rect 13881 29003 13887 29037
rect 13841 28965 13887 29003
rect 13841 28931 13847 28965
rect 13881 28931 13887 28965
rect 13841 28893 13887 28931
rect 13841 28859 13847 28893
rect 13881 28859 13887 28893
rect 13841 28821 13887 28859
rect 13841 28787 13847 28821
rect 13881 28787 13887 28821
rect 13841 28749 13887 28787
rect 13841 28715 13847 28749
rect 13881 28715 13887 28749
rect 13841 28677 13887 28715
rect 13841 28643 13847 28677
rect 13881 28643 13887 28677
rect 13841 28627 13887 28643
rect 14299 29901 14345 29917
rect 14299 29867 14305 29901
rect 14339 29867 14345 29901
rect 14299 29829 14345 29867
rect 14299 29795 14305 29829
rect 14339 29795 14345 29829
rect 14299 29757 14345 29795
rect 14299 29723 14305 29757
rect 14339 29723 14345 29757
rect 14299 29685 14345 29723
rect 14299 29651 14305 29685
rect 14339 29651 14345 29685
rect 14299 29613 14345 29651
rect 14299 29579 14305 29613
rect 14339 29579 14345 29613
rect 14299 29541 14345 29579
rect 14299 29507 14305 29541
rect 14339 29507 14345 29541
rect 14299 29469 14345 29507
rect 14299 29435 14305 29469
rect 14339 29435 14345 29469
rect 14299 29397 14345 29435
rect 14299 29363 14305 29397
rect 14339 29363 14345 29397
rect 14299 29325 14345 29363
rect 14299 29291 14305 29325
rect 14339 29291 14345 29325
rect 14299 29253 14345 29291
rect 14299 29219 14305 29253
rect 14339 29219 14345 29253
rect 14299 29181 14345 29219
rect 14299 29147 14305 29181
rect 14339 29147 14345 29181
rect 14299 29109 14345 29147
rect 14299 29075 14305 29109
rect 14339 29075 14345 29109
rect 14299 29037 14345 29075
rect 14299 29003 14305 29037
rect 14339 29003 14345 29037
rect 14299 28965 14345 29003
rect 14299 28931 14305 28965
rect 14339 28931 14345 28965
rect 14299 28893 14345 28931
rect 14299 28859 14305 28893
rect 14339 28859 14345 28893
rect 14299 28821 14345 28859
rect 14299 28787 14305 28821
rect 14339 28787 14345 28821
rect 14299 28749 14345 28787
rect 14299 28715 14305 28749
rect 14339 28715 14345 28749
rect 14299 28677 14345 28715
rect 14299 28643 14305 28677
rect 14339 28643 14345 28677
rect 14299 28627 14345 28643
rect 14757 29901 14803 29917
rect 14757 29867 14763 29901
rect 14797 29867 14803 29901
rect 14757 29829 14803 29867
rect 14757 29795 14763 29829
rect 14797 29795 14803 29829
rect 14757 29757 14803 29795
rect 14757 29723 14763 29757
rect 14797 29723 14803 29757
rect 14757 29685 14803 29723
rect 14757 29651 14763 29685
rect 14797 29651 14803 29685
rect 14757 29613 14803 29651
rect 14757 29579 14763 29613
rect 14797 29579 14803 29613
rect 14757 29541 14803 29579
rect 14757 29507 14763 29541
rect 14797 29507 14803 29541
rect 14757 29469 14803 29507
rect 14757 29435 14763 29469
rect 14797 29435 14803 29469
rect 14757 29397 14803 29435
rect 14757 29363 14763 29397
rect 14797 29363 14803 29397
rect 14757 29325 14803 29363
rect 14757 29291 14763 29325
rect 14797 29291 14803 29325
rect 14757 29253 14803 29291
rect 14757 29219 14763 29253
rect 14797 29219 14803 29253
rect 14757 29181 14803 29219
rect 14757 29147 14763 29181
rect 14797 29147 14803 29181
rect 14757 29109 14803 29147
rect 14757 29075 14763 29109
rect 14797 29075 14803 29109
rect 14757 29037 14803 29075
rect 14757 29003 14763 29037
rect 14797 29003 14803 29037
rect 14757 28965 14803 29003
rect 14757 28931 14763 28965
rect 14797 28931 14803 28965
rect 14757 28893 14803 28931
rect 14757 28859 14763 28893
rect 14797 28859 14803 28893
rect 14757 28821 14803 28859
rect 14757 28787 14763 28821
rect 14797 28787 14803 28821
rect 14757 28749 14803 28787
rect 14757 28715 14763 28749
rect 14797 28715 14803 28749
rect 14757 28677 14803 28715
rect 14757 28643 14763 28677
rect 14797 28643 14803 28677
rect 14757 28627 14803 28643
rect 15215 29901 15261 29917
rect 15215 29867 15221 29901
rect 15255 29867 15261 29901
rect 15215 29829 15261 29867
rect 15215 29795 15221 29829
rect 15255 29795 15261 29829
rect 15215 29757 15261 29795
rect 15215 29723 15221 29757
rect 15255 29723 15261 29757
rect 15215 29685 15261 29723
rect 15215 29651 15221 29685
rect 15255 29651 15261 29685
rect 15215 29613 15261 29651
rect 15215 29579 15221 29613
rect 15255 29579 15261 29613
rect 15215 29541 15261 29579
rect 15215 29507 15221 29541
rect 15255 29507 15261 29541
rect 15215 29469 15261 29507
rect 15215 29435 15221 29469
rect 15255 29435 15261 29469
rect 15215 29397 15261 29435
rect 15215 29363 15221 29397
rect 15255 29363 15261 29397
rect 15215 29325 15261 29363
rect 15215 29291 15221 29325
rect 15255 29291 15261 29325
rect 15215 29253 15261 29291
rect 15215 29219 15221 29253
rect 15255 29219 15261 29253
rect 15215 29181 15261 29219
rect 15215 29147 15221 29181
rect 15255 29147 15261 29181
rect 15215 29109 15261 29147
rect 15215 29075 15221 29109
rect 15255 29075 15261 29109
rect 15215 29037 15261 29075
rect 15215 29003 15221 29037
rect 15255 29003 15261 29037
rect 15215 28965 15261 29003
rect 15215 28931 15221 28965
rect 15255 28931 15261 28965
rect 15215 28893 15261 28931
rect 15215 28859 15221 28893
rect 15255 28859 15261 28893
rect 15215 28821 15261 28859
rect 15215 28787 15221 28821
rect 15255 28787 15261 28821
rect 15215 28749 15261 28787
rect 15215 28715 15221 28749
rect 15255 28715 15261 28749
rect 15215 28677 15261 28715
rect 15215 28643 15221 28677
rect 15255 28643 15261 28677
rect 15215 28627 15261 28643
rect 15673 29901 15719 29917
rect 15673 29867 15679 29901
rect 15713 29867 15719 29901
rect 15673 29829 15719 29867
rect 15673 29795 15679 29829
rect 15713 29795 15719 29829
rect 15673 29757 15719 29795
rect 15673 29723 15679 29757
rect 15713 29723 15719 29757
rect 15673 29685 15719 29723
rect 15673 29651 15679 29685
rect 15713 29651 15719 29685
rect 15673 29613 15719 29651
rect 15673 29579 15679 29613
rect 15713 29579 15719 29613
rect 15673 29541 15719 29579
rect 15673 29507 15679 29541
rect 15713 29507 15719 29541
rect 15673 29469 15719 29507
rect 15673 29435 15679 29469
rect 15713 29435 15719 29469
rect 15673 29397 15719 29435
rect 15673 29363 15679 29397
rect 15713 29363 15719 29397
rect 15673 29325 15719 29363
rect 15673 29291 15679 29325
rect 15713 29291 15719 29325
rect 15673 29253 15719 29291
rect 15673 29219 15679 29253
rect 15713 29219 15719 29253
rect 15673 29181 15719 29219
rect 15673 29147 15679 29181
rect 15713 29147 15719 29181
rect 15673 29109 15719 29147
rect 15673 29075 15679 29109
rect 15713 29075 15719 29109
rect 15673 29037 15719 29075
rect 15673 29003 15679 29037
rect 15713 29003 15719 29037
rect 15673 28965 15719 29003
rect 15673 28931 15679 28965
rect 15713 28931 15719 28965
rect 15673 28893 15719 28931
rect 15673 28859 15679 28893
rect 15713 28859 15719 28893
rect 15673 28821 15719 28859
rect 15673 28787 15679 28821
rect 15713 28787 15719 28821
rect 15673 28749 15719 28787
rect 15673 28715 15679 28749
rect 15713 28715 15719 28749
rect 15673 28677 15719 28715
rect 15673 28643 15679 28677
rect 15713 28643 15719 28677
rect 15673 28627 15719 28643
rect 16131 29901 16177 29917
rect 16131 29867 16137 29901
rect 16171 29867 16177 29901
rect 16131 29829 16177 29867
rect 16131 29795 16137 29829
rect 16171 29795 16177 29829
rect 16131 29757 16177 29795
rect 16131 29723 16137 29757
rect 16171 29723 16177 29757
rect 16131 29685 16177 29723
rect 16131 29651 16137 29685
rect 16171 29651 16177 29685
rect 16131 29613 16177 29651
rect 16131 29579 16137 29613
rect 16171 29579 16177 29613
rect 16131 29541 16177 29579
rect 16131 29507 16137 29541
rect 16171 29507 16177 29541
rect 16131 29469 16177 29507
rect 16131 29435 16137 29469
rect 16171 29435 16177 29469
rect 16131 29397 16177 29435
rect 16131 29363 16137 29397
rect 16171 29363 16177 29397
rect 16131 29325 16177 29363
rect 16131 29291 16137 29325
rect 16171 29291 16177 29325
rect 16131 29253 16177 29291
rect 16131 29219 16137 29253
rect 16171 29219 16177 29253
rect 16131 29181 16177 29219
rect 16131 29147 16137 29181
rect 16171 29147 16177 29181
rect 16131 29109 16177 29147
rect 16131 29075 16137 29109
rect 16171 29075 16177 29109
rect 16131 29037 16177 29075
rect 16131 29003 16137 29037
rect 16171 29003 16177 29037
rect 16131 28965 16177 29003
rect 16131 28931 16137 28965
rect 16171 28931 16177 28965
rect 16131 28893 16177 28931
rect 16131 28859 16137 28893
rect 16171 28859 16177 28893
rect 16131 28821 16177 28859
rect 16131 28787 16137 28821
rect 16171 28787 16177 28821
rect 16131 28749 16177 28787
rect 16131 28715 16137 28749
rect 16171 28715 16177 28749
rect 16131 28677 16177 28715
rect 16131 28643 16137 28677
rect 16171 28643 16177 28677
rect 16131 28627 16177 28643
rect 16589 29901 16635 29917
rect 16589 29867 16595 29901
rect 16629 29867 16635 29901
rect 16589 29829 16635 29867
rect 16589 29795 16595 29829
rect 16629 29795 16635 29829
rect 16589 29757 16635 29795
rect 16589 29723 16595 29757
rect 16629 29723 16635 29757
rect 16589 29685 16635 29723
rect 16589 29651 16595 29685
rect 16629 29651 16635 29685
rect 16589 29613 16635 29651
rect 16589 29579 16595 29613
rect 16629 29579 16635 29613
rect 16589 29541 16635 29579
rect 16589 29507 16595 29541
rect 16629 29507 16635 29541
rect 16589 29469 16635 29507
rect 16589 29435 16595 29469
rect 16629 29435 16635 29469
rect 16589 29397 16635 29435
rect 16589 29363 16595 29397
rect 16629 29363 16635 29397
rect 16589 29325 16635 29363
rect 16589 29291 16595 29325
rect 16629 29291 16635 29325
rect 16589 29253 16635 29291
rect 16589 29219 16595 29253
rect 16629 29219 16635 29253
rect 16589 29181 16635 29219
rect 16589 29147 16595 29181
rect 16629 29147 16635 29181
rect 16589 29109 16635 29147
rect 16589 29075 16595 29109
rect 16629 29075 16635 29109
rect 16589 29037 16635 29075
rect 16589 29003 16595 29037
rect 16629 29003 16635 29037
rect 16589 28965 16635 29003
rect 16589 28931 16595 28965
rect 16629 28931 16635 28965
rect 16589 28893 16635 28931
rect 16589 28859 16595 28893
rect 16629 28859 16635 28893
rect 16589 28821 16635 28859
rect 16589 28787 16595 28821
rect 16629 28787 16635 28821
rect 16589 28749 16635 28787
rect 16589 28715 16595 28749
rect 16629 28715 16635 28749
rect 16589 28677 16635 28715
rect 16589 28643 16595 28677
rect 16629 28643 16635 28677
rect 16589 28627 16635 28643
rect 17047 29901 17093 29917
rect 17047 29867 17053 29901
rect 17087 29867 17093 29901
rect 17047 29829 17093 29867
rect 17047 29795 17053 29829
rect 17087 29795 17093 29829
rect 17047 29757 17093 29795
rect 17047 29723 17053 29757
rect 17087 29723 17093 29757
rect 17047 29685 17093 29723
rect 17047 29651 17053 29685
rect 17087 29651 17093 29685
rect 17047 29613 17093 29651
rect 17047 29579 17053 29613
rect 17087 29579 17093 29613
rect 17047 29541 17093 29579
rect 17047 29507 17053 29541
rect 17087 29507 17093 29541
rect 17047 29469 17093 29507
rect 17047 29435 17053 29469
rect 17087 29435 17093 29469
rect 17047 29397 17093 29435
rect 17047 29363 17053 29397
rect 17087 29363 17093 29397
rect 17047 29325 17093 29363
rect 17047 29291 17053 29325
rect 17087 29291 17093 29325
rect 17047 29253 17093 29291
rect 17047 29219 17053 29253
rect 17087 29219 17093 29253
rect 17047 29181 17093 29219
rect 17047 29147 17053 29181
rect 17087 29147 17093 29181
rect 17047 29109 17093 29147
rect 17047 29075 17053 29109
rect 17087 29075 17093 29109
rect 17047 29037 17093 29075
rect 17047 29003 17053 29037
rect 17087 29003 17093 29037
rect 17047 28965 17093 29003
rect 17047 28931 17053 28965
rect 17087 28931 17093 28965
rect 17047 28893 17093 28931
rect 17047 28859 17053 28893
rect 17087 28859 17093 28893
rect 17047 28821 17093 28859
rect 17047 28787 17053 28821
rect 17087 28787 17093 28821
rect 17047 28749 17093 28787
rect 17047 28715 17053 28749
rect 17087 28715 17093 28749
rect 17047 28677 17093 28715
rect 17047 28643 17053 28677
rect 17087 28643 17093 28677
rect 17047 28627 17093 28643
rect 17505 29901 17551 29917
rect 17505 29867 17511 29901
rect 17545 29867 17551 29901
rect 17505 29829 17551 29867
rect 17505 29795 17511 29829
rect 17545 29795 17551 29829
rect 17505 29757 17551 29795
rect 17505 29723 17511 29757
rect 17545 29723 17551 29757
rect 17505 29685 17551 29723
rect 17505 29651 17511 29685
rect 17545 29651 17551 29685
rect 17505 29613 17551 29651
rect 17505 29579 17511 29613
rect 17545 29579 17551 29613
rect 17505 29541 17551 29579
rect 17505 29507 17511 29541
rect 17545 29507 17551 29541
rect 17505 29469 17551 29507
rect 17505 29435 17511 29469
rect 17545 29435 17551 29469
rect 17505 29397 17551 29435
rect 17505 29363 17511 29397
rect 17545 29363 17551 29397
rect 17505 29325 17551 29363
rect 17505 29291 17511 29325
rect 17545 29291 17551 29325
rect 17505 29253 17551 29291
rect 17505 29219 17511 29253
rect 17545 29219 17551 29253
rect 17505 29181 17551 29219
rect 17505 29147 17511 29181
rect 17545 29147 17551 29181
rect 17505 29109 17551 29147
rect 17505 29075 17511 29109
rect 17545 29075 17551 29109
rect 17505 29037 17551 29075
rect 17505 29003 17511 29037
rect 17545 29003 17551 29037
rect 17505 28965 17551 29003
rect 17505 28931 17511 28965
rect 17545 28931 17551 28965
rect 17505 28893 17551 28931
rect 17505 28859 17511 28893
rect 17545 28859 17551 28893
rect 17505 28821 17551 28859
rect 17505 28787 17511 28821
rect 17545 28787 17551 28821
rect 17505 28749 17551 28787
rect 17505 28715 17511 28749
rect 17545 28715 17551 28749
rect 17505 28677 17551 28715
rect 17505 28643 17511 28677
rect 17545 28643 17551 28677
rect 17505 28627 17551 28643
rect 17963 29901 18009 29917
rect 17963 29867 17969 29901
rect 18003 29867 18009 29901
rect 17963 29829 18009 29867
rect 17963 29795 17969 29829
rect 18003 29795 18009 29829
rect 17963 29757 18009 29795
rect 17963 29723 17969 29757
rect 18003 29723 18009 29757
rect 17963 29685 18009 29723
rect 17963 29651 17969 29685
rect 18003 29651 18009 29685
rect 17963 29613 18009 29651
rect 17963 29579 17969 29613
rect 18003 29579 18009 29613
rect 17963 29541 18009 29579
rect 17963 29507 17969 29541
rect 18003 29507 18009 29541
rect 17963 29469 18009 29507
rect 17963 29435 17969 29469
rect 18003 29435 18009 29469
rect 17963 29397 18009 29435
rect 17963 29363 17969 29397
rect 18003 29363 18009 29397
rect 17963 29325 18009 29363
rect 17963 29291 17969 29325
rect 18003 29291 18009 29325
rect 17963 29253 18009 29291
rect 17963 29219 17969 29253
rect 18003 29219 18009 29253
rect 17963 29181 18009 29219
rect 17963 29147 17969 29181
rect 18003 29147 18009 29181
rect 17963 29109 18009 29147
rect 17963 29075 17969 29109
rect 18003 29075 18009 29109
rect 17963 29037 18009 29075
rect 17963 29003 17969 29037
rect 18003 29003 18009 29037
rect 17963 28965 18009 29003
rect 17963 28931 17969 28965
rect 18003 28931 18009 28965
rect 17963 28893 18009 28931
rect 17963 28859 17969 28893
rect 18003 28859 18009 28893
rect 17963 28821 18009 28859
rect 17963 28787 17969 28821
rect 18003 28787 18009 28821
rect 17963 28749 18009 28787
rect 17963 28715 17969 28749
rect 18003 28715 18009 28749
rect 17963 28677 18009 28715
rect 17963 28643 17969 28677
rect 18003 28643 18009 28677
rect 17963 28627 18009 28643
rect 18421 29901 18467 29917
rect 18421 29867 18427 29901
rect 18461 29867 18467 29901
rect 18421 29829 18467 29867
rect 18421 29795 18427 29829
rect 18461 29795 18467 29829
rect 18421 29757 18467 29795
rect 18421 29723 18427 29757
rect 18461 29723 18467 29757
rect 18421 29685 18467 29723
rect 18421 29651 18427 29685
rect 18461 29651 18467 29685
rect 18421 29613 18467 29651
rect 18421 29579 18427 29613
rect 18461 29579 18467 29613
rect 18421 29541 18467 29579
rect 18421 29507 18427 29541
rect 18461 29507 18467 29541
rect 18421 29469 18467 29507
rect 18421 29435 18427 29469
rect 18461 29435 18467 29469
rect 18421 29397 18467 29435
rect 18421 29363 18427 29397
rect 18461 29363 18467 29397
rect 18421 29325 18467 29363
rect 18421 29291 18427 29325
rect 18461 29291 18467 29325
rect 18421 29253 18467 29291
rect 18421 29219 18427 29253
rect 18461 29219 18467 29253
rect 18421 29181 18467 29219
rect 18421 29147 18427 29181
rect 18461 29147 18467 29181
rect 18421 29109 18467 29147
rect 18421 29075 18427 29109
rect 18461 29075 18467 29109
rect 18421 29037 18467 29075
rect 18421 29003 18427 29037
rect 18461 29003 18467 29037
rect 18421 28965 18467 29003
rect 18421 28931 18427 28965
rect 18461 28931 18467 28965
rect 18421 28893 18467 28931
rect 18421 28859 18427 28893
rect 18461 28859 18467 28893
rect 18421 28821 18467 28859
rect 18421 28787 18427 28821
rect 18461 28787 18467 28821
rect 18421 28749 18467 28787
rect 18421 28715 18427 28749
rect 18461 28715 18467 28749
rect 18421 28677 18467 28715
rect 18879 29901 18925 29917
rect 18879 29867 18885 29901
rect 18919 29867 18925 29901
rect 18879 29829 18925 29867
rect 18879 29795 18885 29829
rect 18919 29795 18925 29829
rect 18879 29757 18925 29795
rect 18879 29723 18885 29757
rect 18919 29723 18925 29757
rect 18879 29685 18925 29723
rect 18879 29651 18885 29685
rect 18919 29651 18925 29685
rect 18879 29613 18925 29651
rect 18879 29579 18885 29613
rect 18919 29579 18925 29613
rect 18879 29541 18925 29579
rect 18879 29507 18885 29541
rect 18919 29507 18925 29541
rect 18879 29469 18925 29507
rect 18879 29435 18885 29469
rect 18919 29435 18925 29469
rect 18879 29397 18925 29435
rect 18879 29363 18885 29397
rect 18919 29363 18925 29397
rect 18879 29325 18925 29363
rect 18879 29291 18885 29325
rect 18919 29291 18925 29325
rect 18879 29253 18925 29291
rect 18879 29219 18885 29253
rect 18919 29219 18925 29253
rect 18879 29181 18925 29219
rect 18879 29147 18885 29181
rect 18919 29147 18925 29181
rect 18879 29109 18925 29147
rect 18879 29075 18885 29109
rect 18919 29075 18925 29109
rect 18879 29037 18925 29075
rect 18879 29003 18885 29037
rect 18919 29003 18925 29037
rect 18879 28965 18925 29003
rect 18879 28931 18885 28965
rect 18919 28931 18925 28965
rect 18879 28893 18925 28931
rect 18879 28859 18885 28893
rect 18919 28859 18925 28893
rect 18879 28821 18925 28859
rect 18879 28787 18885 28821
rect 18919 28787 18925 28821
rect 18879 28749 18925 28787
rect 18879 28715 18885 28749
rect 18919 28715 18925 28749
rect 18879 28688 18925 28715
rect 19337 29901 19383 29917
rect 19337 29867 19343 29901
rect 19377 29867 19383 29901
rect 19337 29829 19383 29867
rect 19337 29795 19343 29829
rect 19377 29795 19383 29829
rect 19337 29757 19383 29795
rect 19337 29723 19343 29757
rect 19377 29723 19383 29757
rect 19337 29685 19383 29723
rect 19337 29651 19343 29685
rect 19377 29651 19383 29685
rect 19337 29613 19383 29651
rect 19337 29579 19343 29613
rect 19377 29579 19383 29613
rect 19337 29541 19383 29579
rect 19337 29507 19343 29541
rect 19377 29507 19383 29541
rect 19337 29469 19383 29507
rect 19337 29435 19343 29469
rect 19377 29435 19383 29469
rect 19337 29397 19383 29435
rect 19337 29363 19343 29397
rect 19377 29363 19383 29397
rect 19337 29325 19383 29363
rect 19337 29291 19343 29325
rect 19377 29291 19383 29325
rect 19337 29253 19383 29291
rect 19337 29219 19343 29253
rect 19377 29219 19383 29253
rect 19337 29181 19383 29219
rect 19337 29147 19343 29181
rect 19377 29147 19383 29181
rect 19337 29109 19383 29147
rect 19337 29075 19343 29109
rect 19377 29075 19383 29109
rect 19337 29037 19383 29075
rect 19337 29003 19343 29037
rect 19377 29003 19383 29037
rect 19337 28965 19383 29003
rect 19337 28931 19343 28965
rect 19377 28931 19383 28965
rect 19337 28893 19383 28931
rect 19337 28859 19343 28893
rect 19377 28859 19383 28893
rect 19337 28821 19383 28859
rect 19337 28787 19343 28821
rect 19377 28787 19383 28821
rect 19337 28749 19383 28787
rect 19337 28715 19343 28749
rect 19377 28715 19383 28749
rect 18421 28643 18427 28677
rect 18461 28643 18467 28677
rect 18421 28627 18467 28643
rect 18874 28636 18880 28688
rect 18932 28636 18938 28688
rect 19337 28677 19383 28715
rect 19337 28643 19343 28677
rect 19377 28643 19383 28677
rect 18879 28627 18925 28636
rect 19337 28627 19383 28643
rect 19795 29901 19841 29917
rect 19795 29867 19801 29901
rect 19835 29867 19841 29901
rect 19795 29829 19841 29867
rect 19795 29795 19801 29829
rect 19835 29795 19841 29829
rect 19795 29757 19841 29795
rect 19795 29723 19801 29757
rect 19835 29723 19841 29757
rect 19795 29685 19841 29723
rect 19795 29651 19801 29685
rect 19835 29651 19841 29685
rect 19795 29613 19841 29651
rect 19795 29579 19801 29613
rect 19835 29579 19841 29613
rect 19795 29541 19841 29579
rect 19795 29507 19801 29541
rect 19835 29507 19841 29541
rect 19795 29469 19841 29507
rect 19795 29435 19801 29469
rect 19835 29435 19841 29469
rect 19795 29397 19841 29435
rect 19795 29363 19801 29397
rect 19835 29363 19841 29397
rect 19795 29325 19841 29363
rect 19795 29291 19801 29325
rect 19835 29291 19841 29325
rect 19795 29253 19841 29291
rect 19795 29219 19801 29253
rect 19835 29219 19841 29253
rect 19795 29181 19841 29219
rect 19795 29147 19801 29181
rect 19835 29147 19841 29181
rect 19795 29109 19841 29147
rect 19795 29075 19801 29109
rect 19835 29075 19841 29109
rect 19795 29037 19841 29075
rect 19795 29003 19801 29037
rect 19835 29003 19841 29037
rect 19795 28965 19841 29003
rect 19795 28931 19801 28965
rect 19835 28931 19841 28965
rect 19795 28893 19841 28931
rect 19795 28859 19801 28893
rect 19835 28859 19841 28893
rect 19795 28821 19841 28859
rect 19795 28787 19801 28821
rect 19835 28787 19841 28821
rect 19795 28749 19841 28787
rect 19795 28715 19801 28749
rect 19835 28715 19841 28749
rect 19795 28677 19841 28715
rect 19795 28643 19801 28677
rect 19835 28643 19841 28677
rect 19795 28627 19841 28643
rect 20253 29901 20299 29917
rect 20253 29867 20259 29901
rect 20293 29867 20299 29901
rect 20253 29829 20299 29867
rect 20253 29795 20259 29829
rect 20293 29795 20299 29829
rect 20253 29757 20299 29795
rect 20253 29723 20259 29757
rect 20293 29723 20299 29757
rect 20253 29685 20299 29723
rect 20253 29651 20259 29685
rect 20293 29651 20299 29685
rect 20253 29613 20299 29651
rect 20253 29579 20259 29613
rect 20293 29579 20299 29613
rect 20253 29541 20299 29579
rect 20253 29507 20259 29541
rect 20293 29507 20299 29541
rect 20253 29469 20299 29507
rect 20253 29435 20259 29469
rect 20293 29435 20299 29469
rect 20253 29397 20299 29435
rect 20253 29363 20259 29397
rect 20293 29363 20299 29397
rect 20253 29325 20299 29363
rect 20253 29291 20259 29325
rect 20293 29291 20299 29325
rect 20253 29253 20299 29291
rect 20253 29219 20259 29253
rect 20293 29219 20299 29253
rect 20253 29181 20299 29219
rect 20253 29147 20259 29181
rect 20293 29147 20299 29181
rect 20253 29109 20299 29147
rect 20253 29075 20259 29109
rect 20293 29075 20299 29109
rect 20253 29037 20299 29075
rect 20253 29003 20259 29037
rect 20293 29003 20299 29037
rect 20253 28965 20299 29003
rect 20253 28931 20259 28965
rect 20293 28931 20299 28965
rect 20253 28893 20299 28931
rect 20253 28859 20259 28893
rect 20293 28859 20299 28893
rect 20253 28821 20299 28859
rect 20253 28787 20259 28821
rect 20293 28787 20299 28821
rect 20253 28749 20299 28787
rect 20253 28715 20259 28749
rect 20293 28715 20299 28749
rect 20253 28677 20299 28715
rect 20253 28643 20259 28677
rect 20293 28643 20299 28677
rect 20253 28627 20299 28643
rect 20711 29901 20757 29917
rect 20711 29867 20717 29901
rect 20751 29867 20757 29901
rect 20711 29829 20757 29867
rect 20711 29795 20717 29829
rect 20751 29795 20757 29829
rect 20711 29757 20757 29795
rect 20711 29723 20717 29757
rect 20751 29723 20757 29757
rect 20711 29685 20757 29723
rect 20711 29651 20717 29685
rect 20751 29651 20757 29685
rect 20711 29613 20757 29651
rect 20711 29579 20717 29613
rect 20751 29579 20757 29613
rect 20711 29541 20757 29579
rect 20711 29507 20717 29541
rect 20751 29507 20757 29541
rect 20711 29469 20757 29507
rect 20711 29435 20717 29469
rect 20751 29435 20757 29469
rect 20711 29397 20757 29435
rect 20711 29363 20717 29397
rect 20751 29363 20757 29397
rect 20711 29325 20757 29363
rect 20711 29291 20717 29325
rect 20751 29291 20757 29325
rect 20711 29253 20757 29291
rect 20711 29219 20717 29253
rect 20751 29219 20757 29253
rect 20711 29181 20757 29219
rect 20711 29147 20717 29181
rect 20751 29147 20757 29181
rect 20711 29109 20757 29147
rect 20711 29075 20717 29109
rect 20751 29075 20757 29109
rect 20711 29037 20757 29075
rect 20711 29003 20717 29037
rect 20751 29003 20757 29037
rect 20711 28965 20757 29003
rect 20711 28931 20717 28965
rect 20751 28931 20757 28965
rect 20711 28893 20757 28931
rect 20711 28859 20717 28893
rect 20751 28859 20757 28893
rect 20711 28821 20757 28859
rect 20711 28787 20717 28821
rect 20751 28787 20757 28821
rect 20711 28749 20757 28787
rect 20711 28715 20717 28749
rect 20751 28715 20757 28749
rect 20711 28677 20757 28715
rect 20711 28643 20717 28677
rect 20751 28643 20757 28677
rect 20711 28627 20757 28643
rect 21169 29901 21215 29917
rect 21169 29867 21175 29901
rect 21209 29867 21215 29901
rect 21169 29829 21215 29867
rect 21169 29795 21175 29829
rect 21209 29795 21215 29829
rect 21169 29757 21215 29795
rect 21169 29723 21175 29757
rect 21209 29723 21215 29757
rect 21169 29685 21215 29723
rect 21169 29651 21175 29685
rect 21209 29651 21215 29685
rect 21169 29613 21215 29651
rect 21169 29579 21175 29613
rect 21209 29579 21215 29613
rect 21169 29541 21215 29579
rect 21169 29507 21175 29541
rect 21209 29507 21215 29541
rect 21169 29469 21215 29507
rect 21169 29435 21175 29469
rect 21209 29435 21215 29469
rect 21169 29397 21215 29435
rect 21169 29363 21175 29397
rect 21209 29363 21215 29397
rect 21169 29325 21215 29363
rect 21169 29291 21175 29325
rect 21209 29291 21215 29325
rect 21169 29253 21215 29291
rect 21169 29219 21175 29253
rect 21209 29219 21215 29253
rect 21169 29181 21215 29219
rect 21169 29147 21175 29181
rect 21209 29147 21215 29181
rect 21169 29109 21215 29147
rect 21169 29075 21175 29109
rect 21209 29075 21215 29109
rect 21169 29037 21215 29075
rect 21169 29003 21175 29037
rect 21209 29003 21215 29037
rect 21169 28965 21215 29003
rect 21169 28931 21175 28965
rect 21209 28931 21215 28965
rect 21169 28893 21215 28931
rect 21169 28859 21175 28893
rect 21209 28859 21215 28893
rect 21169 28821 21215 28859
rect 21169 28787 21175 28821
rect 21209 28787 21215 28821
rect 21169 28749 21215 28787
rect 21169 28715 21175 28749
rect 21209 28715 21215 28749
rect 21169 28677 21215 28715
rect 21169 28643 21175 28677
rect 21209 28643 21215 28677
rect 21169 28627 21215 28643
rect 21627 29901 21673 29917
rect 21627 29867 21633 29901
rect 21667 29867 21673 29901
rect 21627 29829 21673 29867
rect 21627 29795 21633 29829
rect 21667 29795 21673 29829
rect 21627 29757 21673 29795
rect 21627 29723 21633 29757
rect 21667 29723 21673 29757
rect 21627 29685 21673 29723
rect 21627 29651 21633 29685
rect 21667 29651 21673 29685
rect 21627 29613 21673 29651
rect 21627 29579 21633 29613
rect 21667 29579 21673 29613
rect 21627 29541 21673 29579
rect 21627 29507 21633 29541
rect 21667 29507 21673 29541
rect 21627 29469 21673 29507
rect 21627 29435 21633 29469
rect 21667 29435 21673 29469
rect 21627 29397 21673 29435
rect 21627 29363 21633 29397
rect 21667 29363 21673 29397
rect 21627 29325 21673 29363
rect 21627 29291 21633 29325
rect 21667 29291 21673 29325
rect 21627 29253 21673 29291
rect 21627 29219 21633 29253
rect 21667 29219 21673 29253
rect 21627 29181 21673 29219
rect 21627 29147 21633 29181
rect 21667 29147 21673 29181
rect 21627 29109 21673 29147
rect 21627 29075 21633 29109
rect 21667 29075 21673 29109
rect 21627 29037 21673 29075
rect 21627 29003 21633 29037
rect 21667 29003 21673 29037
rect 21627 28965 21673 29003
rect 21627 28931 21633 28965
rect 21667 28931 21673 28965
rect 21627 28893 21673 28931
rect 21627 28859 21633 28893
rect 21667 28859 21673 28893
rect 21627 28821 21673 28859
rect 21627 28787 21633 28821
rect 21667 28787 21673 28821
rect 21627 28749 21673 28787
rect 21627 28715 21633 28749
rect 21667 28715 21673 28749
rect 21627 28677 21673 28715
rect 21627 28643 21633 28677
rect 21667 28643 21673 28677
rect 21627 28627 21673 28643
rect 22085 29901 22131 29917
rect 22085 29867 22091 29901
rect 22125 29867 22131 29901
rect 22085 29829 22131 29867
rect 22085 29795 22091 29829
rect 22125 29795 22131 29829
rect 22085 29757 22131 29795
rect 22085 29723 22091 29757
rect 22125 29723 22131 29757
rect 22085 29685 22131 29723
rect 22085 29651 22091 29685
rect 22125 29651 22131 29685
rect 22085 29613 22131 29651
rect 22085 29579 22091 29613
rect 22125 29579 22131 29613
rect 22085 29541 22131 29579
rect 22085 29507 22091 29541
rect 22125 29507 22131 29541
rect 22085 29469 22131 29507
rect 22085 29435 22091 29469
rect 22125 29435 22131 29469
rect 22085 29397 22131 29435
rect 22085 29363 22091 29397
rect 22125 29363 22131 29397
rect 22085 29325 22131 29363
rect 22085 29291 22091 29325
rect 22125 29291 22131 29325
rect 22085 29253 22131 29291
rect 22085 29219 22091 29253
rect 22125 29219 22131 29253
rect 22085 29181 22131 29219
rect 22085 29147 22091 29181
rect 22125 29147 22131 29181
rect 22085 29109 22131 29147
rect 22085 29075 22091 29109
rect 22125 29075 22131 29109
rect 22085 29037 22131 29075
rect 22085 29003 22091 29037
rect 22125 29003 22131 29037
rect 22085 28965 22131 29003
rect 22085 28931 22091 28965
rect 22125 28931 22131 28965
rect 22085 28893 22131 28931
rect 22085 28859 22091 28893
rect 22125 28859 22131 28893
rect 22085 28821 22131 28859
rect 22085 28787 22091 28821
rect 22125 28787 22131 28821
rect 22085 28749 22131 28787
rect 22085 28715 22091 28749
rect 22125 28715 22131 28749
rect 22085 28677 22131 28715
rect 22085 28643 22091 28677
rect 22125 28643 22131 28677
rect 22085 28627 22131 28643
rect 22543 29901 22589 29917
rect 22543 29867 22549 29901
rect 22583 29867 22589 29901
rect 22543 29829 22589 29867
rect 22543 29795 22549 29829
rect 22583 29795 22589 29829
rect 22543 29757 22589 29795
rect 22543 29723 22549 29757
rect 22583 29723 22589 29757
rect 22543 29685 22589 29723
rect 22543 29651 22549 29685
rect 22583 29651 22589 29685
rect 22543 29613 22589 29651
rect 22543 29579 22549 29613
rect 22583 29579 22589 29613
rect 22543 29541 22589 29579
rect 22543 29507 22549 29541
rect 22583 29507 22589 29541
rect 22543 29469 22589 29507
rect 22543 29435 22549 29469
rect 22583 29435 22589 29469
rect 22543 29397 22589 29435
rect 22543 29363 22549 29397
rect 22583 29363 22589 29397
rect 22543 29325 22589 29363
rect 22543 29291 22549 29325
rect 22583 29291 22589 29325
rect 22543 29253 22589 29291
rect 22543 29219 22549 29253
rect 22583 29219 22589 29253
rect 22543 29181 22589 29219
rect 22543 29147 22549 29181
rect 22583 29147 22589 29181
rect 22543 29109 22589 29147
rect 22543 29075 22549 29109
rect 22583 29075 22589 29109
rect 22543 29037 22589 29075
rect 22543 29003 22549 29037
rect 22583 29003 22589 29037
rect 22543 28965 22589 29003
rect 22543 28931 22549 28965
rect 22583 28931 22589 28965
rect 22543 28893 22589 28931
rect 22543 28859 22549 28893
rect 22583 28859 22589 28893
rect 22543 28821 22589 28859
rect 22543 28787 22549 28821
rect 22583 28787 22589 28821
rect 22543 28749 22589 28787
rect 22543 28715 22549 28749
rect 22583 28715 22589 28749
rect 22543 28677 22589 28715
rect 22543 28643 22549 28677
rect 22583 28643 22589 28677
rect 22543 28627 22589 28643
rect 23001 29901 23047 29917
rect 23001 29867 23007 29901
rect 23041 29867 23047 29901
rect 23001 29829 23047 29867
rect 23001 29795 23007 29829
rect 23041 29795 23047 29829
rect 23001 29757 23047 29795
rect 23001 29723 23007 29757
rect 23041 29723 23047 29757
rect 23001 29685 23047 29723
rect 23001 29651 23007 29685
rect 23041 29651 23047 29685
rect 23001 29613 23047 29651
rect 23001 29579 23007 29613
rect 23041 29579 23047 29613
rect 23001 29541 23047 29579
rect 23001 29507 23007 29541
rect 23041 29507 23047 29541
rect 23001 29469 23047 29507
rect 23001 29435 23007 29469
rect 23041 29435 23047 29469
rect 23001 29397 23047 29435
rect 23001 29363 23007 29397
rect 23041 29363 23047 29397
rect 23001 29325 23047 29363
rect 23001 29291 23007 29325
rect 23041 29291 23047 29325
rect 23001 29253 23047 29291
rect 23001 29219 23007 29253
rect 23041 29219 23047 29253
rect 23001 29181 23047 29219
rect 23001 29147 23007 29181
rect 23041 29147 23047 29181
rect 23001 29109 23047 29147
rect 23001 29075 23007 29109
rect 23041 29075 23047 29109
rect 23001 29037 23047 29075
rect 23001 29003 23007 29037
rect 23041 29003 23047 29037
rect 23001 28965 23047 29003
rect 23001 28931 23007 28965
rect 23041 28931 23047 28965
rect 23001 28893 23047 28931
rect 23001 28859 23007 28893
rect 23041 28859 23047 28893
rect 23001 28821 23047 28859
rect 23001 28787 23007 28821
rect 23041 28787 23047 28821
rect 23001 28749 23047 28787
rect 23001 28715 23007 28749
rect 23041 28715 23047 28749
rect 23001 28677 23047 28715
rect 23001 28643 23007 28677
rect 23041 28643 23047 28677
rect 23001 28627 23047 28643
rect 23459 29901 23505 29917
rect 23459 29867 23465 29901
rect 23499 29867 23505 29901
rect 23459 29829 23505 29867
rect 23459 29795 23465 29829
rect 23499 29795 23505 29829
rect 23459 29757 23505 29795
rect 23459 29723 23465 29757
rect 23499 29723 23505 29757
rect 23459 29685 23505 29723
rect 23459 29651 23465 29685
rect 23499 29651 23505 29685
rect 23459 29613 23505 29651
rect 23459 29579 23465 29613
rect 23499 29579 23505 29613
rect 23459 29541 23505 29579
rect 23459 29507 23465 29541
rect 23499 29507 23505 29541
rect 23459 29469 23505 29507
rect 23459 29435 23465 29469
rect 23499 29435 23505 29469
rect 23459 29397 23505 29435
rect 23459 29363 23465 29397
rect 23499 29363 23505 29397
rect 23459 29325 23505 29363
rect 23459 29291 23465 29325
rect 23499 29291 23505 29325
rect 23459 29253 23505 29291
rect 23459 29219 23465 29253
rect 23499 29219 23505 29253
rect 23459 29181 23505 29219
rect 23459 29147 23465 29181
rect 23499 29147 23505 29181
rect 23459 29109 23505 29147
rect 23459 29075 23465 29109
rect 23499 29075 23505 29109
rect 23459 29037 23505 29075
rect 23459 29003 23465 29037
rect 23499 29003 23505 29037
rect 23459 28965 23505 29003
rect 23459 28931 23465 28965
rect 23499 28931 23505 28965
rect 23459 28893 23505 28931
rect 23459 28859 23465 28893
rect 23499 28859 23505 28893
rect 23459 28821 23505 28859
rect 23459 28787 23465 28821
rect 23499 28787 23505 28821
rect 23459 28749 23505 28787
rect 23459 28715 23465 28749
rect 23499 28715 23505 28749
rect 23459 28677 23505 28715
rect 23459 28643 23465 28677
rect 23499 28643 23505 28677
rect 23459 28627 23505 28643
rect 23917 29901 23963 29917
rect 23917 29867 23923 29901
rect 23957 29867 23963 29901
rect 23917 29829 23963 29867
rect 23917 29795 23923 29829
rect 23957 29795 23963 29829
rect 23917 29757 23963 29795
rect 23917 29723 23923 29757
rect 23957 29723 23963 29757
rect 23917 29685 23963 29723
rect 23917 29651 23923 29685
rect 23957 29651 23963 29685
rect 23917 29613 23963 29651
rect 23917 29579 23923 29613
rect 23957 29579 23963 29613
rect 23917 29541 23963 29579
rect 23917 29507 23923 29541
rect 23957 29507 23963 29541
rect 23917 29469 23963 29507
rect 23917 29435 23923 29469
rect 23957 29435 23963 29469
rect 23917 29397 23963 29435
rect 23917 29363 23923 29397
rect 23957 29363 23963 29397
rect 23917 29325 23963 29363
rect 23917 29291 23923 29325
rect 23957 29291 23963 29325
rect 23917 29253 23963 29291
rect 23917 29219 23923 29253
rect 23957 29219 23963 29253
rect 23917 29181 23963 29219
rect 23917 29147 23923 29181
rect 23957 29147 23963 29181
rect 23917 29109 23963 29147
rect 23917 29075 23923 29109
rect 23957 29075 23963 29109
rect 23917 29037 23963 29075
rect 23917 29003 23923 29037
rect 23957 29003 23963 29037
rect 23917 28965 23963 29003
rect 23917 28931 23923 28965
rect 23957 28931 23963 28965
rect 23917 28893 23963 28931
rect 23917 28859 23923 28893
rect 23957 28859 23963 28893
rect 23917 28821 23963 28859
rect 23917 28787 23923 28821
rect 23957 28787 23963 28821
rect 23917 28749 23963 28787
rect 23917 28715 23923 28749
rect 23957 28715 23963 28749
rect 23917 28677 23963 28715
rect 23917 28643 23923 28677
rect 23957 28643 23963 28677
rect 23917 28627 23963 28643
rect 24375 29901 24421 29917
rect 24375 29867 24381 29901
rect 24415 29867 24421 29901
rect 24375 29829 24421 29867
rect 24375 29795 24381 29829
rect 24415 29795 24421 29829
rect 24375 29757 24421 29795
rect 24375 29723 24381 29757
rect 24415 29723 24421 29757
rect 24375 29685 24421 29723
rect 24375 29651 24381 29685
rect 24415 29651 24421 29685
rect 24375 29613 24421 29651
rect 24375 29579 24381 29613
rect 24415 29579 24421 29613
rect 24375 29541 24421 29579
rect 24375 29507 24381 29541
rect 24415 29507 24421 29541
rect 24375 29469 24421 29507
rect 24375 29435 24381 29469
rect 24415 29435 24421 29469
rect 24375 29397 24421 29435
rect 24375 29363 24381 29397
rect 24415 29363 24421 29397
rect 24375 29325 24421 29363
rect 24375 29291 24381 29325
rect 24415 29291 24421 29325
rect 24375 29253 24421 29291
rect 24375 29219 24381 29253
rect 24415 29219 24421 29253
rect 24375 29181 24421 29219
rect 24375 29147 24381 29181
rect 24415 29147 24421 29181
rect 24375 29109 24421 29147
rect 24375 29075 24381 29109
rect 24415 29075 24421 29109
rect 24375 29037 24421 29075
rect 24375 29003 24381 29037
rect 24415 29003 24421 29037
rect 24375 28965 24421 29003
rect 24375 28931 24381 28965
rect 24415 28931 24421 28965
rect 24375 28893 24421 28931
rect 24375 28859 24381 28893
rect 24415 28859 24421 28893
rect 24375 28821 24421 28859
rect 24375 28787 24381 28821
rect 24415 28787 24421 28821
rect 24375 28749 24421 28787
rect 24375 28715 24381 28749
rect 24415 28715 24421 28749
rect 24375 28677 24421 28715
rect 24375 28643 24381 28677
rect 24415 28643 24421 28677
rect 24375 28627 24421 28643
rect 24833 29901 24879 29917
rect 24833 29867 24839 29901
rect 24873 29867 24879 29901
rect 24833 29829 24879 29867
rect 24833 29795 24839 29829
rect 24873 29795 24879 29829
rect 24833 29757 24879 29795
rect 24833 29723 24839 29757
rect 24873 29723 24879 29757
rect 24833 29685 24879 29723
rect 24833 29651 24839 29685
rect 24873 29651 24879 29685
rect 24833 29613 24879 29651
rect 24833 29579 24839 29613
rect 24873 29579 24879 29613
rect 24833 29541 24879 29579
rect 24833 29507 24839 29541
rect 24873 29507 24879 29541
rect 24833 29469 24879 29507
rect 24833 29435 24839 29469
rect 24873 29435 24879 29469
rect 24833 29397 24879 29435
rect 24833 29363 24839 29397
rect 24873 29363 24879 29397
rect 24833 29325 24879 29363
rect 24833 29291 24839 29325
rect 24873 29291 24879 29325
rect 24833 29253 24879 29291
rect 24833 29219 24839 29253
rect 24873 29219 24879 29253
rect 24833 29181 24879 29219
rect 24833 29147 24839 29181
rect 24873 29147 24879 29181
rect 24833 29109 24879 29147
rect 24833 29075 24839 29109
rect 24873 29075 24879 29109
rect 24833 29037 24879 29075
rect 24833 29003 24839 29037
rect 24873 29003 24879 29037
rect 24833 28965 24879 29003
rect 24833 28931 24839 28965
rect 24873 28931 24879 28965
rect 24833 28893 24879 28931
rect 24833 28859 24839 28893
rect 24873 28859 24879 28893
rect 24833 28821 24879 28859
rect 24833 28787 24839 28821
rect 24873 28787 24879 28821
rect 24833 28749 24879 28787
rect 24833 28715 24839 28749
rect 24873 28715 24879 28749
rect 24833 28677 24879 28715
rect 24833 28643 24839 28677
rect 24873 28643 24879 28677
rect 24833 28627 24879 28643
rect 25291 29901 25337 29917
rect 25291 29867 25297 29901
rect 25331 29867 25337 29901
rect 25291 29829 25337 29867
rect 25291 29795 25297 29829
rect 25331 29795 25337 29829
rect 25291 29757 25337 29795
rect 25291 29723 25297 29757
rect 25331 29723 25337 29757
rect 25291 29685 25337 29723
rect 25291 29651 25297 29685
rect 25331 29651 25337 29685
rect 25291 29613 25337 29651
rect 25291 29579 25297 29613
rect 25331 29579 25337 29613
rect 25291 29541 25337 29579
rect 25291 29507 25297 29541
rect 25331 29507 25337 29541
rect 25291 29469 25337 29507
rect 25291 29435 25297 29469
rect 25331 29435 25337 29469
rect 25291 29397 25337 29435
rect 25291 29363 25297 29397
rect 25331 29363 25337 29397
rect 25291 29325 25337 29363
rect 25291 29291 25297 29325
rect 25331 29291 25337 29325
rect 25291 29253 25337 29291
rect 25291 29219 25297 29253
rect 25331 29219 25337 29253
rect 25291 29181 25337 29219
rect 25291 29147 25297 29181
rect 25331 29147 25337 29181
rect 25291 29109 25337 29147
rect 25291 29075 25297 29109
rect 25331 29075 25337 29109
rect 25291 29037 25337 29075
rect 25291 29003 25297 29037
rect 25331 29003 25337 29037
rect 25291 28965 25337 29003
rect 25291 28931 25297 28965
rect 25331 28931 25337 28965
rect 25291 28893 25337 28931
rect 25291 28859 25297 28893
rect 25331 28859 25337 28893
rect 25291 28821 25337 28859
rect 25291 28787 25297 28821
rect 25331 28787 25337 28821
rect 25291 28749 25337 28787
rect 25291 28715 25297 28749
rect 25331 28715 25337 28749
rect 25291 28677 25337 28715
rect 25291 28643 25297 28677
rect 25331 28643 25337 28677
rect 25291 28627 25337 28643
rect 25749 29901 25795 29917
rect 25749 29867 25755 29901
rect 25789 29867 25795 29901
rect 25749 29829 25795 29867
rect 25749 29795 25755 29829
rect 25789 29795 25795 29829
rect 25749 29757 25795 29795
rect 25749 29723 25755 29757
rect 25789 29723 25795 29757
rect 25749 29685 25795 29723
rect 25749 29651 25755 29685
rect 25789 29651 25795 29685
rect 25749 29613 25795 29651
rect 25749 29579 25755 29613
rect 25789 29579 25795 29613
rect 25749 29541 25795 29579
rect 25749 29507 25755 29541
rect 25789 29507 25795 29541
rect 25749 29469 25795 29507
rect 25749 29435 25755 29469
rect 25789 29435 25795 29469
rect 25749 29397 25795 29435
rect 25749 29363 25755 29397
rect 25789 29363 25795 29397
rect 25749 29325 25795 29363
rect 25749 29291 25755 29325
rect 25789 29291 25795 29325
rect 25749 29253 25795 29291
rect 25749 29219 25755 29253
rect 25789 29219 25795 29253
rect 25749 29181 25795 29219
rect 25749 29147 25755 29181
rect 25789 29147 25795 29181
rect 25749 29109 25795 29147
rect 25749 29075 25755 29109
rect 25789 29075 25795 29109
rect 25749 29037 25795 29075
rect 25749 29003 25755 29037
rect 25789 29003 25795 29037
rect 25749 28965 25795 29003
rect 25749 28931 25755 28965
rect 25789 28931 25795 28965
rect 25749 28893 25795 28931
rect 25749 28859 25755 28893
rect 25789 28859 25795 28893
rect 25749 28821 25795 28859
rect 25749 28787 25755 28821
rect 25789 28787 25795 28821
rect 25749 28749 25795 28787
rect 25749 28715 25755 28749
rect 25789 28715 25795 28749
rect 25749 28677 25795 28715
rect 25749 28643 25755 28677
rect 25789 28643 25795 28677
rect 25749 28627 25795 28643
rect 26207 29901 26253 29917
rect 26207 29867 26213 29901
rect 26247 29867 26253 29901
rect 26207 29829 26253 29867
rect 26207 29795 26213 29829
rect 26247 29795 26253 29829
rect 26207 29757 26253 29795
rect 26207 29723 26213 29757
rect 26247 29723 26253 29757
rect 26207 29685 26253 29723
rect 26207 29651 26213 29685
rect 26247 29651 26253 29685
rect 26207 29613 26253 29651
rect 26207 29579 26213 29613
rect 26247 29579 26253 29613
rect 26207 29541 26253 29579
rect 26207 29507 26213 29541
rect 26247 29507 26253 29541
rect 26207 29469 26253 29507
rect 26207 29435 26213 29469
rect 26247 29435 26253 29469
rect 26207 29397 26253 29435
rect 26207 29363 26213 29397
rect 26247 29363 26253 29397
rect 26207 29325 26253 29363
rect 26207 29291 26213 29325
rect 26247 29291 26253 29325
rect 26207 29253 26253 29291
rect 26207 29219 26213 29253
rect 26247 29219 26253 29253
rect 26207 29181 26253 29219
rect 26207 29147 26213 29181
rect 26247 29147 26253 29181
rect 26207 29109 26253 29147
rect 26207 29075 26213 29109
rect 26247 29075 26253 29109
rect 26207 29037 26253 29075
rect 26207 29003 26213 29037
rect 26247 29003 26253 29037
rect 26207 28965 26253 29003
rect 26207 28931 26213 28965
rect 26247 28931 26253 28965
rect 26207 28893 26253 28931
rect 26207 28859 26213 28893
rect 26247 28859 26253 28893
rect 26207 28821 26253 28859
rect 26207 28787 26213 28821
rect 26247 28787 26253 28821
rect 26207 28749 26253 28787
rect 26207 28715 26213 28749
rect 26247 28715 26253 28749
rect 26207 28677 26253 28715
rect 26207 28643 26213 28677
rect 26247 28643 26253 28677
rect 26207 28627 26253 28643
rect 26665 29901 26711 29917
rect 26665 29867 26671 29901
rect 26705 29867 26711 29901
rect 26665 29829 26711 29867
rect 26665 29795 26671 29829
rect 26705 29795 26711 29829
rect 26665 29757 26711 29795
rect 26665 29723 26671 29757
rect 26705 29723 26711 29757
rect 26665 29685 26711 29723
rect 26665 29651 26671 29685
rect 26705 29651 26711 29685
rect 26665 29613 26711 29651
rect 26665 29579 26671 29613
rect 26705 29579 26711 29613
rect 26665 29541 26711 29579
rect 26665 29507 26671 29541
rect 26705 29507 26711 29541
rect 26665 29469 26711 29507
rect 26665 29435 26671 29469
rect 26705 29435 26711 29469
rect 26665 29397 26711 29435
rect 26665 29363 26671 29397
rect 26705 29363 26711 29397
rect 26665 29325 26711 29363
rect 26665 29291 26671 29325
rect 26705 29291 26711 29325
rect 26665 29253 26711 29291
rect 26665 29219 26671 29253
rect 26705 29219 26711 29253
rect 26665 29181 26711 29219
rect 26665 29147 26671 29181
rect 26705 29147 26711 29181
rect 26665 29109 26711 29147
rect 26665 29075 26671 29109
rect 26705 29075 26711 29109
rect 26665 29037 26711 29075
rect 26665 29003 26671 29037
rect 26705 29003 26711 29037
rect 26665 28965 26711 29003
rect 26665 28931 26671 28965
rect 26705 28931 26711 28965
rect 26665 28893 26711 28931
rect 26665 28859 26671 28893
rect 26705 28859 26711 28893
rect 26665 28821 26711 28859
rect 26665 28787 26671 28821
rect 26705 28787 26711 28821
rect 26665 28749 26711 28787
rect 26665 28715 26671 28749
rect 26705 28715 26711 28749
rect 26665 28677 26711 28715
rect 26665 28643 26671 28677
rect 26705 28643 26711 28677
rect 26665 28627 26711 28643
rect 27123 29901 27169 29917
rect 27123 29867 27129 29901
rect 27163 29867 27169 29901
rect 27123 29829 27169 29867
rect 27123 29795 27129 29829
rect 27163 29795 27169 29829
rect 27123 29757 27169 29795
rect 27123 29723 27129 29757
rect 27163 29723 27169 29757
rect 27123 29685 27169 29723
rect 27123 29651 27129 29685
rect 27163 29651 27169 29685
rect 27123 29613 27169 29651
rect 27123 29579 27129 29613
rect 27163 29579 27169 29613
rect 27123 29541 27169 29579
rect 27123 29507 27129 29541
rect 27163 29507 27169 29541
rect 27123 29469 27169 29507
rect 27123 29435 27129 29469
rect 27163 29435 27169 29469
rect 27123 29397 27169 29435
rect 27123 29363 27129 29397
rect 27163 29363 27169 29397
rect 27123 29325 27169 29363
rect 27123 29291 27129 29325
rect 27163 29291 27169 29325
rect 27123 29253 27169 29291
rect 27123 29219 27129 29253
rect 27163 29219 27169 29253
rect 27123 29181 27169 29219
rect 27123 29147 27129 29181
rect 27163 29147 27169 29181
rect 27123 29109 27169 29147
rect 27123 29075 27129 29109
rect 27163 29075 27169 29109
rect 27123 29037 27169 29075
rect 27123 29003 27129 29037
rect 27163 29003 27169 29037
rect 27123 28965 27169 29003
rect 27123 28931 27129 28965
rect 27163 28931 27169 28965
rect 27123 28893 27169 28931
rect 27123 28859 27129 28893
rect 27163 28859 27169 28893
rect 27123 28821 27169 28859
rect 27123 28787 27129 28821
rect 27163 28787 27169 28821
rect 27123 28749 27169 28787
rect 27123 28715 27129 28749
rect 27163 28715 27169 28749
rect 27123 28677 27169 28715
rect 27123 28643 27129 28677
rect 27163 28643 27169 28677
rect 27123 28627 27169 28643
rect 27581 29901 27627 29917
rect 27581 29867 27587 29901
rect 27621 29867 27627 29901
rect 27581 29829 27627 29867
rect 27581 29795 27587 29829
rect 27621 29795 27627 29829
rect 27581 29757 27627 29795
rect 27581 29723 27587 29757
rect 27621 29723 27627 29757
rect 27581 29685 27627 29723
rect 27581 29651 27587 29685
rect 27621 29651 27627 29685
rect 27581 29613 27627 29651
rect 27581 29579 27587 29613
rect 27621 29579 27627 29613
rect 27581 29541 27627 29579
rect 27581 29507 27587 29541
rect 27621 29507 27627 29541
rect 27581 29469 27627 29507
rect 27581 29435 27587 29469
rect 27621 29435 27627 29469
rect 27581 29397 27627 29435
rect 27581 29363 27587 29397
rect 27621 29363 27627 29397
rect 27581 29325 27627 29363
rect 27581 29291 27587 29325
rect 27621 29291 27627 29325
rect 27581 29253 27627 29291
rect 27581 29219 27587 29253
rect 27621 29219 27627 29253
rect 27581 29181 27627 29219
rect 27581 29147 27587 29181
rect 27621 29147 27627 29181
rect 27581 29109 27627 29147
rect 27581 29075 27587 29109
rect 27621 29075 27627 29109
rect 27581 29037 27627 29075
rect 27581 29003 27587 29037
rect 27621 29003 27627 29037
rect 27581 28965 27627 29003
rect 27581 28931 27587 28965
rect 27621 28931 27627 28965
rect 27581 28893 27627 28931
rect 27581 28859 27587 28893
rect 27621 28859 27627 28893
rect 27581 28821 27627 28859
rect 27581 28787 27587 28821
rect 27621 28787 27627 28821
rect 27581 28749 27627 28787
rect 27581 28715 27587 28749
rect 27621 28715 27627 28749
rect 27581 28677 27627 28715
rect 27581 28643 27587 28677
rect 27621 28643 27627 28677
rect 27581 28627 27627 28643
rect 28039 29901 28085 29917
rect 28039 29867 28045 29901
rect 28079 29867 28085 29901
rect 28039 29829 28085 29867
rect 28039 29795 28045 29829
rect 28079 29795 28085 29829
rect 28039 29757 28085 29795
rect 28039 29723 28045 29757
rect 28079 29723 28085 29757
rect 28039 29685 28085 29723
rect 28039 29651 28045 29685
rect 28079 29651 28085 29685
rect 28039 29613 28085 29651
rect 28039 29579 28045 29613
rect 28079 29579 28085 29613
rect 28039 29541 28085 29579
rect 28039 29507 28045 29541
rect 28079 29507 28085 29541
rect 28039 29469 28085 29507
rect 28039 29435 28045 29469
rect 28079 29435 28085 29469
rect 28039 29397 28085 29435
rect 28039 29363 28045 29397
rect 28079 29363 28085 29397
rect 28039 29325 28085 29363
rect 28039 29291 28045 29325
rect 28079 29291 28085 29325
rect 28039 29253 28085 29291
rect 28039 29219 28045 29253
rect 28079 29219 28085 29253
rect 28039 29181 28085 29219
rect 28039 29147 28045 29181
rect 28079 29147 28085 29181
rect 28039 29109 28085 29147
rect 28039 29075 28045 29109
rect 28079 29075 28085 29109
rect 28039 29037 28085 29075
rect 28039 29003 28045 29037
rect 28079 29003 28085 29037
rect 28039 28965 28085 29003
rect 28039 28931 28045 28965
rect 28079 28931 28085 28965
rect 28039 28893 28085 28931
rect 28039 28859 28045 28893
rect 28079 28859 28085 28893
rect 28039 28821 28085 28859
rect 28039 28787 28045 28821
rect 28079 28787 28085 28821
rect 28039 28749 28085 28787
rect 28039 28715 28045 28749
rect 28079 28715 28085 28749
rect 28039 28677 28085 28715
rect 28039 28643 28045 28677
rect 28079 28643 28085 28677
rect 28039 28627 28085 28643
rect 28497 29901 28543 29917
rect 28497 29867 28503 29901
rect 28537 29867 28543 29901
rect 28497 29829 28543 29867
rect 28497 29795 28503 29829
rect 28537 29795 28543 29829
rect 28497 29757 28543 29795
rect 28497 29723 28503 29757
rect 28537 29723 28543 29757
rect 28497 29685 28543 29723
rect 28497 29651 28503 29685
rect 28537 29651 28543 29685
rect 28497 29613 28543 29651
rect 28497 29579 28503 29613
rect 28537 29579 28543 29613
rect 28497 29541 28543 29579
rect 28497 29507 28503 29541
rect 28537 29507 28543 29541
rect 28497 29469 28543 29507
rect 28497 29435 28503 29469
rect 28537 29435 28543 29469
rect 28497 29397 28543 29435
rect 28497 29363 28503 29397
rect 28537 29363 28543 29397
rect 28497 29325 28543 29363
rect 28497 29291 28503 29325
rect 28537 29291 28543 29325
rect 28497 29253 28543 29291
rect 28497 29219 28503 29253
rect 28537 29219 28543 29253
rect 28497 29181 28543 29219
rect 28497 29147 28503 29181
rect 28537 29147 28543 29181
rect 28497 29109 28543 29147
rect 28497 29075 28503 29109
rect 28537 29075 28543 29109
rect 28497 29037 28543 29075
rect 28497 29003 28503 29037
rect 28537 29003 28543 29037
rect 28497 28965 28543 29003
rect 28497 28931 28503 28965
rect 28537 28931 28543 28965
rect 28497 28893 28543 28931
rect 28497 28859 28503 28893
rect 28537 28859 28543 28893
rect 28497 28821 28543 28859
rect 28497 28787 28503 28821
rect 28537 28787 28543 28821
rect 28497 28749 28543 28787
rect 28497 28715 28503 28749
rect 28537 28715 28543 28749
rect 28497 28677 28543 28715
rect 28497 28643 28503 28677
rect 28537 28643 28543 28677
rect 28497 28627 28543 28643
rect 28955 29901 29001 29917
rect 28955 29867 28961 29901
rect 28995 29867 29001 29901
rect 28955 29829 29001 29867
rect 28955 29795 28961 29829
rect 28995 29795 29001 29829
rect 28955 29757 29001 29795
rect 28955 29723 28961 29757
rect 28995 29723 29001 29757
rect 28955 29685 29001 29723
rect 28955 29651 28961 29685
rect 28995 29651 29001 29685
rect 28955 29613 29001 29651
rect 28955 29579 28961 29613
rect 28995 29579 29001 29613
rect 28955 29541 29001 29579
rect 28955 29507 28961 29541
rect 28995 29507 29001 29541
rect 28955 29469 29001 29507
rect 28955 29435 28961 29469
rect 28995 29435 29001 29469
rect 28955 29397 29001 29435
rect 28955 29363 28961 29397
rect 28995 29363 29001 29397
rect 28955 29325 29001 29363
rect 28955 29291 28961 29325
rect 28995 29291 29001 29325
rect 28955 29253 29001 29291
rect 28955 29219 28961 29253
rect 28995 29219 29001 29253
rect 28955 29181 29001 29219
rect 28955 29147 28961 29181
rect 28995 29147 29001 29181
rect 28955 29109 29001 29147
rect 28955 29075 28961 29109
rect 28995 29075 29001 29109
rect 28955 29037 29001 29075
rect 28955 29003 28961 29037
rect 28995 29003 29001 29037
rect 28955 28965 29001 29003
rect 28955 28931 28961 28965
rect 28995 28931 29001 28965
rect 28955 28893 29001 28931
rect 28955 28859 28961 28893
rect 28995 28859 29001 28893
rect 28955 28821 29001 28859
rect 28955 28787 28961 28821
rect 28995 28787 29001 28821
rect 28955 28749 29001 28787
rect 28955 28715 28961 28749
rect 28995 28715 29001 28749
rect 28955 28677 29001 28715
rect 28955 28643 28961 28677
rect 28995 28643 29001 28677
rect 28955 28627 29001 28643
rect 29413 29901 29459 29917
rect 29413 29867 29419 29901
rect 29453 29867 29459 29901
rect 29413 29829 29459 29867
rect 29413 29795 29419 29829
rect 29453 29795 29459 29829
rect 29413 29757 29459 29795
rect 29413 29723 29419 29757
rect 29453 29723 29459 29757
rect 29413 29685 29459 29723
rect 29413 29651 29419 29685
rect 29453 29651 29459 29685
rect 29413 29613 29459 29651
rect 29413 29579 29419 29613
rect 29453 29579 29459 29613
rect 29413 29541 29459 29579
rect 29413 29507 29419 29541
rect 29453 29507 29459 29541
rect 29413 29469 29459 29507
rect 29413 29435 29419 29469
rect 29453 29435 29459 29469
rect 29413 29397 29459 29435
rect 29413 29363 29419 29397
rect 29453 29363 29459 29397
rect 29413 29325 29459 29363
rect 29413 29291 29419 29325
rect 29453 29291 29459 29325
rect 29413 29253 29459 29291
rect 29413 29219 29419 29253
rect 29453 29219 29459 29253
rect 29413 29181 29459 29219
rect 29413 29147 29419 29181
rect 29453 29147 29459 29181
rect 29413 29109 29459 29147
rect 29413 29075 29419 29109
rect 29453 29075 29459 29109
rect 29413 29037 29459 29075
rect 29413 29003 29419 29037
rect 29453 29003 29459 29037
rect 29413 28965 29459 29003
rect 29413 28931 29419 28965
rect 29453 28931 29459 28965
rect 29413 28893 29459 28931
rect 29413 28859 29419 28893
rect 29453 28859 29459 28893
rect 29413 28821 29459 28859
rect 29413 28787 29419 28821
rect 29453 28787 29459 28821
rect 29413 28749 29459 28787
rect 29413 28715 29419 28749
rect 29453 28715 29459 28749
rect 29413 28677 29459 28715
rect 29413 28643 29419 28677
rect 29453 28643 29459 28677
rect 29413 28627 29459 28643
rect 29871 29901 29917 29917
rect 29871 29867 29877 29901
rect 29911 29867 29917 29901
rect 29871 29829 29917 29867
rect 29871 29795 29877 29829
rect 29911 29795 29917 29829
rect 29871 29757 29917 29795
rect 29871 29723 29877 29757
rect 29911 29723 29917 29757
rect 29871 29685 29917 29723
rect 29871 29651 29877 29685
rect 29911 29651 29917 29685
rect 29871 29613 29917 29651
rect 29871 29579 29877 29613
rect 29911 29579 29917 29613
rect 29871 29541 29917 29579
rect 29871 29507 29877 29541
rect 29911 29507 29917 29541
rect 29871 29469 29917 29507
rect 29871 29435 29877 29469
rect 29911 29435 29917 29469
rect 29871 29397 29917 29435
rect 29871 29363 29877 29397
rect 29911 29363 29917 29397
rect 29871 29325 29917 29363
rect 29871 29291 29877 29325
rect 29911 29291 29917 29325
rect 29871 29253 29917 29291
rect 29871 29219 29877 29253
rect 29911 29219 29917 29253
rect 29871 29181 29917 29219
rect 29871 29147 29877 29181
rect 29911 29147 29917 29181
rect 29871 29109 29917 29147
rect 29871 29075 29877 29109
rect 29911 29075 29917 29109
rect 29871 29037 29917 29075
rect 29871 29003 29877 29037
rect 29911 29003 29917 29037
rect 29871 28965 29917 29003
rect 29871 28931 29877 28965
rect 29911 28931 29917 28965
rect 29871 28893 29917 28931
rect 29871 28859 29877 28893
rect 29911 28859 29917 28893
rect 29871 28821 29917 28859
rect 29871 28787 29877 28821
rect 29911 28787 29917 28821
rect 29871 28749 29917 28787
rect 29871 28715 29877 28749
rect 29911 28715 29917 28749
rect 29871 28677 29917 28715
rect 29871 28643 29877 28677
rect 29911 28643 29917 28677
rect 29871 28627 29917 28643
rect 30329 29901 30375 29917
rect 30329 29867 30335 29901
rect 30369 29867 30375 29901
rect 30329 29829 30375 29867
rect 30329 29795 30335 29829
rect 30369 29795 30375 29829
rect 30329 29757 30375 29795
rect 30329 29723 30335 29757
rect 30369 29723 30375 29757
rect 30329 29685 30375 29723
rect 30329 29651 30335 29685
rect 30369 29651 30375 29685
rect 30329 29613 30375 29651
rect 30329 29579 30335 29613
rect 30369 29579 30375 29613
rect 30329 29541 30375 29579
rect 30329 29507 30335 29541
rect 30369 29507 30375 29541
rect 30329 29469 30375 29507
rect 30329 29435 30335 29469
rect 30369 29435 30375 29469
rect 30329 29397 30375 29435
rect 30329 29363 30335 29397
rect 30369 29363 30375 29397
rect 30329 29325 30375 29363
rect 30329 29291 30335 29325
rect 30369 29291 30375 29325
rect 30329 29253 30375 29291
rect 30329 29219 30335 29253
rect 30369 29219 30375 29253
rect 30329 29181 30375 29219
rect 30329 29147 30335 29181
rect 30369 29147 30375 29181
rect 30329 29109 30375 29147
rect 30329 29075 30335 29109
rect 30369 29075 30375 29109
rect 30329 29037 30375 29075
rect 30329 29003 30335 29037
rect 30369 29003 30375 29037
rect 30329 28965 30375 29003
rect 30329 28931 30335 28965
rect 30369 28931 30375 28965
rect 30329 28893 30375 28931
rect 30329 28859 30335 28893
rect 30369 28859 30375 28893
rect 30329 28821 30375 28859
rect 30329 28787 30335 28821
rect 30369 28787 30375 28821
rect 30329 28749 30375 28787
rect 30329 28715 30335 28749
rect 30369 28715 30375 28749
rect 30329 28677 30375 28715
rect 30329 28643 30335 28677
rect 30369 28643 30375 28677
rect 30329 28627 30375 28643
rect 30787 29901 30833 29917
rect 30787 29867 30793 29901
rect 30827 29867 30833 29901
rect 30787 29829 30833 29867
rect 30787 29795 30793 29829
rect 30827 29795 30833 29829
rect 30787 29757 30833 29795
rect 30787 29723 30793 29757
rect 30827 29723 30833 29757
rect 30787 29685 30833 29723
rect 30787 29651 30793 29685
rect 30827 29651 30833 29685
rect 30787 29613 30833 29651
rect 30787 29579 30793 29613
rect 30827 29579 30833 29613
rect 30787 29541 30833 29579
rect 30787 29507 30793 29541
rect 30827 29507 30833 29541
rect 30787 29469 30833 29507
rect 30787 29435 30793 29469
rect 30827 29435 30833 29469
rect 30787 29397 30833 29435
rect 30787 29363 30793 29397
rect 30827 29363 30833 29397
rect 30787 29325 30833 29363
rect 30787 29291 30793 29325
rect 30827 29291 30833 29325
rect 30787 29253 30833 29291
rect 30787 29219 30793 29253
rect 30827 29219 30833 29253
rect 30787 29181 30833 29219
rect 30787 29147 30793 29181
rect 30827 29147 30833 29181
rect 30787 29109 30833 29147
rect 30787 29075 30793 29109
rect 30827 29075 30833 29109
rect 30787 29037 30833 29075
rect 30787 29003 30793 29037
rect 30827 29003 30833 29037
rect 30787 28965 30833 29003
rect 30787 28931 30793 28965
rect 30827 28931 30833 28965
rect 30787 28893 30833 28931
rect 30787 28859 30793 28893
rect 30827 28859 30833 28893
rect 30787 28821 30833 28859
rect 30787 28787 30793 28821
rect 30827 28787 30833 28821
rect 30787 28749 30833 28787
rect 30787 28715 30793 28749
rect 30827 28715 30833 28749
rect 30787 28677 30833 28715
rect 30787 28643 30793 28677
rect 30827 28643 30833 28677
rect 30787 28627 30833 28643
rect 31245 29901 31291 29917
rect 31245 29867 31251 29901
rect 31285 29867 31291 29901
rect 31245 29829 31291 29867
rect 31245 29795 31251 29829
rect 31285 29795 31291 29829
rect 31245 29757 31291 29795
rect 31245 29723 31251 29757
rect 31285 29723 31291 29757
rect 31245 29685 31291 29723
rect 31245 29651 31251 29685
rect 31285 29651 31291 29685
rect 31245 29613 31291 29651
rect 31245 29579 31251 29613
rect 31285 29579 31291 29613
rect 31245 29541 31291 29579
rect 31245 29507 31251 29541
rect 31285 29507 31291 29541
rect 31245 29469 31291 29507
rect 31245 29435 31251 29469
rect 31285 29435 31291 29469
rect 31245 29397 31291 29435
rect 31245 29363 31251 29397
rect 31285 29363 31291 29397
rect 31245 29325 31291 29363
rect 31245 29291 31251 29325
rect 31285 29291 31291 29325
rect 31245 29253 31291 29291
rect 31245 29219 31251 29253
rect 31285 29219 31291 29253
rect 31245 29181 31291 29219
rect 31245 29147 31251 29181
rect 31285 29147 31291 29181
rect 31245 29109 31291 29147
rect 31245 29075 31251 29109
rect 31285 29075 31291 29109
rect 31245 29037 31291 29075
rect 31245 29003 31251 29037
rect 31285 29003 31291 29037
rect 31245 28965 31291 29003
rect 31245 28931 31251 28965
rect 31285 28931 31291 28965
rect 31245 28893 31291 28931
rect 31245 28859 31251 28893
rect 31285 28859 31291 28893
rect 31245 28821 31291 28859
rect 31245 28787 31251 28821
rect 31285 28787 31291 28821
rect 31245 28749 31291 28787
rect 31245 28715 31251 28749
rect 31285 28715 31291 28749
rect 31245 28677 31291 28715
rect 31245 28643 31251 28677
rect 31285 28643 31291 28677
rect 31245 28627 31291 28643
rect 31703 29901 31749 29917
rect 31703 29867 31709 29901
rect 31743 29867 31749 29901
rect 31703 29829 31749 29867
rect 31703 29795 31709 29829
rect 31743 29795 31749 29829
rect 31703 29757 31749 29795
rect 31703 29723 31709 29757
rect 31743 29723 31749 29757
rect 31703 29685 31749 29723
rect 31703 29651 31709 29685
rect 31743 29651 31749 29685
rect 31703 29613 31749 29651
rect 31703 29579 31709 29613
rect 31743 29579 31749 29613
rect 31703 29541 31749 29579
rect 31703 29507 31709 29541
rect 31743 29507 31749 29541
rect 31703 29469 31749 29507
rect 31703 29435 31709 29469
rect 31743 29435 31749 29469
rect 31703 29397 31749 29435
rect 31703 29363 31709 29397
rect 31743 29363 31749 29397
rect 31703 29325 31749 29363
rect 31703 29291 31709 29325
rect 31743 29291 31749 29325
rect 31703 29253 31749 29291
rect 31703 29219 31709 29253
rect 31743 29219 31749 29253
rect 31703 29181 31749 29219
rect 31703 29147 31709 29181
rect 31743 29147 31749 29181
rect 31703 29109 31749 29147
rect 31703 29075 31709 29109
rect 31743 29075 31749 29109
rect 31703 29037 31749 29075
rect 31703 29003 31709 29037
rect 31743 29003 31749 29037
rect 31703 28965 31749 29003
rect 31703 28931 31709 28965
rect 31743 28931 31749 28965
rect 31703 28893 31749 28931
rect 31703 28859 31709 28893
rect 31743 28859 31749 28893
rect 31703 28821 31749 28859
rect 31703 28787 31709 28821
rect 31743 28787 31749 28821
rect 31703 28749 31749 28787
rect 31703 28715 31709 28749
rect 31743 28715 31749 28749
rect 31703 28677 31749 28715
rect 31703 28643 31709 28677
rect 31743 28643 31749 28677
rect 31703 28627 31749 28643
rect 32161 29901 32207 29917
rect 32161 29867 32167 29901
rect 32201 29867 32207 29901
rect 32161 29829 32207 29867
rect 32161 29795 32167 29829
rect 32201 29795 32207 29829
rect 32161 29757 32207 29795
rect 32161 29723 32167 29757
rect 32201 29723 32207 29757
rect 32161 29685 32207 29723
rect 32161 29651 32167 29685
rect 32201 29651 32207 29685
rect 32161 29613 32207 29651
rect 32161 29579 32167 29613
rect 32201 29579 32207 29613
rect 32161 29541 32207 29579
rect 32161 29507 32167 29541
rect 32201 29507 32207 29541
rect 32161 29469 32207 29507
rect 32161 29435 32167 29469
rect 32201 29435 32207 29469
rect 32161 29397 32207 29435
rect 32161 29363 32167 29397
rect 32201 29363 32207 29397
rect 32161 29325 32207 29363
rect 32161 29291 32167 29325
rect 32201 29291 32207 29325
rect 32161 29253 32207 29291
rect 32161 29219 32167 29253
rect 32201 29219 32207 29253
rect 32161 29181 32207 29219
rect 32161 29147 32167 29181
rect 32201 29147 32207 29181
rect 32161 29109 32207 29147
rect 32161 29075 32167 29109
rect 32201 29075 32207 29109
rect 32161 29037 32207 29075
rect 32161 29003 32167 29037
rect 32201 29003 32207 29037
rect 32161 28965 32207 29003
rect 32161 28931 32167 28965
rect 32201 28931 32207 28965
rect 32161 28893 32207 28931
rect 32161 28859 32167 28893
rect 32201 28859 32207 28893
rect 32161 28821 32207 28859
rect 32161 28787 32167 28821
rect 32201 28787 32207 28821
rect 32161 28749 32207 28787
rect 32161 28715 32167 28749
rect 32201 28715 32207 28749
rect 32161 28677 32207 28715
rect 32161 28643 32167 28677
rect 32201 28643 32207 28677
rect 32161 28627 32207 28643
rect 32619 29901 32665 29917
rect 32619 29867 32625 29901
rect 32659 29867 32665 29901
rect 32619 29829 32665 29867
rect 32619 29795 32625 29829
rect 32659 29795 32665 29829
rect 32619 29757 32665 29795
rect 32619 29723 32625 29757
rect 32659 29723 32665 29757
rect 32619 29685 32665 29723
rect 32619 29651 32625 29685
rect 32659 29651 32665 29685
rect 32619 29613 32665 29651
rect 32619 29579 32625 29613
rect 32659 29579 32665 29613
rect 32619 29541 32665 29579
rect 32619 29507 32625 29541
rect 32659 29507 32665 29541
rect 32619 29469 32665 29507
rect 32619 29435 32625 29469
rect 32659 29435 32665 29469
rect 32619 29397 32665 29435
rect 32619 29363 32625 29397
rect 32659 29363 32665 29397
rect 32619 29325 32665 29363
rect 32619 29291 32625 29325
rect 32659 29291 32665 29325
rect 32619 29253 32665 29291
rect 32619 29219 32625 29253
rect 32659 29219 32665 29253
rect 32619 29181 32665 29219
rect 32619 29147 32625 29181
rect 32659 29147 32665 29181
rect 32619 29109 32665 29147
rect 32619 29075 32625 29109
rect 32659 29075 32665 29109
rect 32619 29037 32665 29075
rect 32619 29003 32625 29037
rect 32659 29003 32665 29037
rect 32619 28965 32665 29003
rect 32619 28931 32625 28965
rect 32659 28931 32665 28965
rect 32619 28893 32665 28931
rect 32619 28859 32625 28893
rect 32659 28859 32665 28893
rect 32619 28821 32665 28859
rect 32619 28787 32625 28821
rect 32659 28787 32665 28821
rect 32619 28749 32665 28787
rect 32619 28715 32625 28749
rect 32659 28715 32665 28749
rect 32619 28677 32665 28715
rect 32619 28643 32625 28677
rect 32659 28643 32665 28677
rect 32619 28627 32665 28643
rect 33077 29901 33123 29917
rect 33077 29867 33083 29901
rect 33117 29867 33123 29901
rect 33077 29829 33123 29867
rect 33077 29795 33083 29829
rect 33117 29795 33123 29829
rect 33077 29757 33123 29795
rect 33077 29723 33083 29757
rect 33117 29723 33123 29757
rect 33077 29685 33123 29723
rect 33077 29651 33083 29685
rect 33117 29651 33123 29685
rect 33077 29613 33123 29651
rect 33077 29579 33083 29613
rect 33117 29579 33123 29613
rect 33077 29541 33123 29579
rect 33077 29507 33083 29541
rect 33117 29507 33123 29541
rect 33077 29469 33123 29507
rect 33077 29435 33083 29469
rect 33117 29435 33123 29469
rect 33077 29397 33123 29435
rect 33077 29363 33083 29397
rect 33117 29363 33123 29397
rect 33077 29325 33123 29363
rect 33077 29291 33083 29325
rect 33117 29291 33123 29325
rect 33077 29253 33123 29291
rect 33077 29219 33083 29253
rect 33117 29219 33123 29253
rect 33077 29181 33123 29219
rect 33077 29147 33083 29181
rect 33117 29147 33123 29181
rect 33077 29109 33123 29147
rect 33077 29075 33083 29109
rect 33117 29075 33123 29109
rect 33077 29037 33123 29075
rect 33077 29003 33083 29037
rect 33117 29003 33123 29037
rect 33077 28965 33123 29003
rect 33077 28931 33083 28965
rect 33117 28931 33123 28965
rect 33077 28893 33123 28931
rect 33077 28859 33083 28893
rect 33117 28859 33123 28893
rect 33077 28821 33123 28859
rect 33077 28787 33083 28821
rect 33117 28787 33123 28821
rect 33077 28749 33123 28787
rect 33077 28715 33083 28749
rect 33117 28715 33123 28749
rect 33077 28677 33123 28715
rect 33077 28643 33083 28677
rect 33117 28643 33123 28677
rect 33077 28627 33123 28643
rect 33535 29901 33581 29917
rect 33535 29867 33541 29901
rect 33575 29867 33581 29901
rect 33535 29829 33581 29867
rect 33535 29795 33541 29829
rect 33575 29795 33581 29829
rect 33535 29757 33581 29795
rect 33535 29723 33541 29757
rect 33575 29723 33581 29757
rect 33535 29685 33581 29723
rect 33535 29651 33541 29685
rect 33575 29651 33581 29685
rect 33535 29613 33581 29651
rect 33535 29579 33541 29613
rect 33575 29579 33581 29613
rect 33535 29541 33581 29579
rect 33535 29507 33541 29541
rect 33575 29507 33581 29541
rect 33535 29469 33581 29507
rect 33535 29435 33541 29469
rect 33575 29435 33581 29469
rect 33535 29397 33581 29435
rect 33535 29363 33541 29397
rect 33575 29363 33581 29397
rect 33535 29325 33581 29363
rect 33535 29291 33541 29325
rect 33575 29291 33581 29325
rect 33535 29253 33581 29291
rect 33535 29219 33541 29253
rect 33575 29219 33581 29253
rect 33535 29181 33581 29219
rect 33535 29147 33541 29181
rect 33575 29147 33581 29181
rect 33535 29109 33581 29147
rect 33535 29075 33541 29109
rect 33575 29075 33581 29109
rect 33535 29037 33581 29075
rect 33535 29003 33541 29037
rect 33575 29003 33581 29037
rect 33535 28965 33581 29003
rect 33535 28931 33541 28965
rect 33575 28931 33581 28965
rect 33535 28893 33581 28931
rect 33535 28859 33541 28893
rect 33575 28859 33581 28893
rect 33535 28821 33581 28859
rect 33535 28787 33541 28821
rect 33575 28787 33581 28821
rect 33535 28749 33581 28787
rect 33535 28715 33541 28749
rect 33575 28715 33581 28749
rect 33535 28677 33581 28715
rect 33535 28643 33541 28677
rect 33575 28643 33581 28677
rect 34083 29901 34129 29917
rect 34083 29867 34089 29901
rect 34123 29867 34129 29901
rect 34083 29829 34129 29867
rect 34083 29795 34089 29829
rect 34123 29795 34129 29829
rect 34083 29757 34129 29795
rect 34083 29723 34089 29757
rect 34123 29723 34129 29757
rect 34083 29685 34129 29723
rect 34083 29651 34089 29685
rect 34123 29651 34129 29685
rect 34083 29613 34129 29651
rect 34083 29579 34089 29613
rect 34123 29579 34129 29613
rect 34083 29541 34129 29579
rect 34083 29507 34089 29541
rect 34123 29507 34129 29541
rect 34083 29469 34129 29507
rect 34083 29435 34089 29469
rect 34123 29435 34129 29469
rect 34083 29397 34129 29435
rect 34083 29363 34089 29397
rect 34123 29363 34129 29397
rect 34083 29325 34129 29363
rect 34083 29291 34089 29325
rect 34123 29291 34129 29325
rect 34083 29253 34129 29291
rect 34083 29219 34089 29253
rect 34123 29219 34129 29253
rect 34083 29181 34129 29219
rect 34083 29147 34089 29181
rect 34123 29147 34129 29181
rect 34083 29109 34129 29147
rect 34083 29075 34089 29109
rect 34123 29075 34129 29109
rect 34083 29037 34129 29075
rect 34083 29003 34089 29037
rect 34123 29003 34129 29037
rect 34083 28965 34129 29003
rect 34083 28931 34089 28965
rect 34123 28931 34129 28965
rect 34083 28893 34129 28931
rect 34083 28859 34089 28893
rect 34123 28859 34129 28893
rect 34083 28821 34129 28859
rect 34083 28787 34089 28821
rect 34123 28787 34129 28821
rect 34083 28749 34129 28787
rect 34083 28715 34089 28749
rect 34123 28715 34129 28749
rect 34083 28677 34129 28715
rect 34083 28676 34089 28677
rect 33535 28627 33581 28643
rect 33612 28648 34089 28676
rect 26510 28500 26516 28552
rect 26568 28540 26574 28552
rect 33612 28540 33640 28648
rect 34083 28643 34089 28648
rect 34123 28643 34129 28677
rect 34083 28627 34129 28643
rect 34541 29901 34587 29917
rect 34541 29867 34547 29901
rect 34581 29867 34587 29901
rect 34541 29829 34587 29867
rect 34541 29795 34547 29829
rect 34581 29795 34587 29829
rect 34541 29757 34587 29795
rect 34541 29723 34547 29757
rect 34581 29723 34587 29757
rect 34541 29685 34587 29723
rect 34541 29651 34547 29685
rect 34581 29651 34587 29685
rect 34541 29613 34587 29651
rect 34541 29579 34547 29613
rect 34581 29579 34587 29613
rect 34541 29541 34587 29579
rect 34541 29507 34547 29541
rect 34581 29507 34587 29541
rect 34541 29469 34587 29507
rect 34541 29435 34547 29469
rect 34581 29435 34587 29469
rect 34541 29397 34587 29435
rect 34541 29363 34547 29397
rect 34581 29363 34587 29397
rect 34541 29325 34587 29363
rect 34541 29291 34547 29325
rect 34581 29291 34587 29325
rect 34541 29253 34587 29291
rect 34541 29219 34547 29253
rect 34581 29219 34587 29253
rect 34541 29181 34587 29219
rect 34541 29147 34547 29181
rect 34581 29147 34587 29181
rect 34541 29109 34587 29147
rect 34541 29075 34547 29109
rect 34581 29075 34587 29109
rect 34541 29037 34587 29075
rect 34541 29003 34547 29037
rect 34581 29003 34587 29037
rect 34541 28965 34587 29003
rect 34541 28931 34547 28965
rect 34581 28931 34587 28965
rect 34541 28893 34587 28931
rect 34541 28859 34547 28893
rect 34581 28859 34587 28893
rect 34541 28821 34587 28859
rect 34541 28787 34547 28821
rect 34581 28787 34587 28821
rect 34541 28749 34587 28787
rect 34541 28715 34547 28749
rect 34581 28715 34587 28749
rect 34541 28677 34587 28715
rect 34541 28643 34547 28677
rect 34581 28643 34587 28677
rect 34541 28627 34587 28643
rect 34999 29901 35045 29917
rect 34999 29867 35005 29901
rect 35039 29867 35045 29901
rect 35360 29900 35388 30092
rect 38028 30008 39896 30036
rect 35457 29901 35503 29917
rect 35457 29900 35463 29901
rect 35360 29872 35463 29900
rect 34999 29829 35045 29867
rect 34999 29795 35005 29829
rect 35039 29795 35045 29829
rect 34999 29757 35045 29795
rect 34999 29723 35005 29757
rect 35039 29723 35045 29757
rect 34999 29685 35045 29723
rect 34999 29651 35005 29685
rect 35039 29651 35045 29685
rect 34999 29613 35045 29651
rect 34999 29579 35005 29613
rect 35039 29579 35045 29613
rect 34999 29541 35045 29579
rect 34999 29507 35005 29541
rect 35039 29507 35045 29541
rect 34999 29469 35045 29507
rect 34999 29435 35005 29469
rect 35039 29435 35045 29469
rect 34999 29397 35045 29435
rect 34999 29363 35005 29397
rect 35039 29363 35045 29397
rect 34999 29325 35045 29363
rect 34999 29291 35005 29325
rect 35039 29291 35045 29325
rect 34999 29253 35045 29291
rect 34999 29219 35005 29253
rect 35039 29219 35045 29253
rect 34999 29181 35045 29219
rect 34999 29147 35005 29181
rect 35039 29147 35045 29181
rect 34999 29109 35045 29147
rect 34999 29075 35005 29109
rect 35039 29075 35045 29109
rect 34999 29037 35045 29075
rect 34999 29003 35005 29037
rect 35039 29003 35045 29037
rect 34999 28965 35045 29003
rect 34999 28931 35005 28965
rect 35039 28931 35045 28965
rect 34999 28893 35045 28931
rect 34999 28859 35005 28893
rect 35039 28859 35045 28893
rect 34999 28821 35045 28859
rect 34999 28787 35005 28821
rect 35039 28787 35045 28821
rect 34999 28749 35045 28787
rect 34999 28715 35005 28749
rect 35039 28715 35045 28749
rect 34999 28677 35045 28715
rect 34999 28643 35005 28677
rect 35039 28643 35045 28677
rect 34999 28627 35045 28643
rect 35457 29867 35463 29872
rect 35497 29867 35503 29901
rect 35457 29829 35503 29867
rect 35457 29795 35463 29829
rect 35497 29795 35503 29829
rect 35457 29757 35503 29795
rect 35457 29723 35463 29757
rect 35497 29723 35503 29757
rect 35457 29685 35503 29723
rect 35457 29651 35463 29685
rect 35497 29651 35503 29685
rect 35457 29613 35503 29651
rect 35457 29579 35463 29613
rect 35497 29579 35503 29613
rect 35457 29541 35503 29579
rect 35457 29507 35463 29541
rect 35497 29507 35503 29541
rect 35457 29469 35503 29507
rect 35457 29435 35463 29469
rect 35497 29435 35503 29469
rect 35457 29397 35503 29435
rect 35457 29363 35463 29397
rect 35497 29363 35503 29397
rect 35457 29325 35503 29363
rect 35457 29291 35463 29325
rect 35497 29291 35503 29325
rect 35457 29253 35503 29291
rect 35457 29219 35463 29253
rect 35497 29219 35503 29253
rect 35457 29181 35503 29219
rect 35457 29147 35463 29181
rect 35497 29147 35503 29181
rect 35457 29109 35503 29147
rect 35457 29075 35463 29109
rect 35497 29075 35503 29109
rect 35457 29037 35503 29075
rect 35457 29003 35463 29037
rect 35497 29003 35503 29037
rect 35457 28965 35503 29003
rect 35457 28931 35463 28965
rect 35497 28931 35503 28965
rect 35457 28893 35503 28931
rect 35457 28859 35463 28893
rect 35497 28859 35503 28893
rect 35457 28821 35503 28859
rect 35457 28787 35463 28821
rect 35497 28787 35503 28821
rect 35457 28749 35503 28787
rect 35457 28715 35463 28749
rect 35497 28715 35503 28749
rect 35457 28677 35503 28715
rect 35457 28643 35463 28677
rect 35497 28643 35503 28677
rect 35457 28627 35503 28643
rect 35915 29901 35961 29917
rect 35915 29867 35921 29901
rect 35955 29867 35961 29901
rect 35915 29829 35961 29867
rect 35915 29795 35921 29829
rect 35955 29795 35961 29829
rect 35915 29757 35961 29795
rect 35915 29723 35921 29757
rect 35955 29723 35961 29757
rect 35915 29685 35961 29723
rect 35915 29651 35921 29685
rect 35955 29651 35961 29685
rect 35915 29613 35961 29651
rect 35915 29579 35921 29613
rect 35955 29579 35961 29613
rect 35915 29541 35961 29579
rect 35915 29507 35921 29541
rect 35955 29507 35961 29541
rect 35915 29469 35961 29507
rect 35915 29435 35921 29469
rect 35955 29435 35961 29469
rect 35915 29397 35961 29435
rect 35915 29363 35921 29397
rect 35955 29363 35961 29397
rect 35915 29325 35961 29363
rect 35915 29291 35921 29325
rect 35955 29291 35961 29325
rect 35915 29253 35961 29291
rect 35915 29219 35921 29253
rect 35955 29219 35961 29253
rect 35915 29181 35961 29219
rect 35915 29147 35921 29181
rect 35955 29147 35961 29181
rect 35915 29109 35961 29147
rect 35915 29075 35921 29109
rect 35955 29075 35961 29109
rect 35915 29037 35961 29075
rect 35915 29003 35921 29037
rect 35955 29003 35961 29037
rect 35915 28965 35961 29003
rect 35915 28931 35921 28965
rect 35955 28931 35961 28965
rect 35915 28893 35961 28931
rect 35915 28859 35921 28893
rect 35955 28859 35961 28893
rect 35915 28821 35961 28859
rect 35915 28787 35921 28821
rect 35955 28787 35961 28821
rect 35915 28749 35961 28787
rect 35915 28715 35921 28749
rect 35955 28715 35961 28749
rect 35915 28677 35961 28715
rect 35915 28643 35921 28677
rect 35955 28643 35961 28677
rect 35915 28627 35961 28643
rect 36373 29901 36419 29917
rect 36373 29867 36379 29901
rect 36413 29867 36419 29901
rect 36373 29829 36419 29867
rect 36373 29795 36379 29829
rect 36413 29795 36419 29829
rect 36373 29757 36419 29795
rect 36373 29723 36379 29757
rect 36413 29723 36419 29757
rect 36373 29685 36419 29723
rect 36373 29651 36379 29685
rect 36413 29651 36419 29685
rect 36373 29613 36419 29651
rect 36373 29579 36379 29613
rect 36413 29579 36419 29613
rect 36373 29541 36419 29579
rect 36373 29507 36379 29541
rect 36413 29507 36419 29541
rect 36373 29469 36419 29507
rect 36373 29435 36379 29469
rect 36413 29435 36419 29469
rect 36373 29397 36419 29435
rect 36373 29363 36379 29397
rect 36413 29363 36419 29397
rect 36373 29325 36419 29363
rect 36373 29291 36379 29325
rect 36413 29291 36419 29325
rect 36373 29253 36419 29291
rect 36373 29219 36379 29253
rect 36413 29219 36419 29253
rect 36373 29181 36419 29219
rect 36373 29147 36379 29181
rect 36413 29147 36419 29181
rect 36373 29109 36419 29147
rect 36373 29075 36379 29109
rect 36413 29075 36419 29109
rect 36373 29037 36419 29075
rect 36373 29003 36379 29037
rect 36413 29003 36419 29037
rect 36373 28965 36419 29003
rect 36373 28931 36379 28965
rect 36413 28931 36419 28965
rect 36373 28893 36419 28931
rect 36373 28859 36379 28893
rect 36413 28859 36419 28893
rect 36373 28821 36419 28859
rect 36373 28787 36379 28821
rect 36413 28787 36419 28821
rect 36373 28749 36419 28787
rect 36373 28715 36379 28749
rect 36413 28715 36419 28749
rect 36373 28677 36419 28715
rect 36373 28643 36379 28677
rect 36413 28643 36419 28677
rect 36373 28627 36419 28643
rect 36831 29901 36877 29917
rect 36831 29867 36837 29901
rect 36871 29867 36877 29901
rect 36831 29829 36877 29867
rect 36831 29795 36837 29829
rect 36871 29795 36877 29829
rect 36831 29757 36877 29795
rect 36831 29723 36837 29757
rect 36871 29723 36877 29757
rect 36831 29685 36877 29723
rect 36831 29651 36837 29685
rect 36871 29651 36877 29685
rect 36831 29613 36877 29651
rect 36831 29579 36837 29613
rect 36871 29579 36877 29613
rect 36831 29541 36877 29579
rect 36831 29507 36837 29541
rect 36871 29507 36877 29541
rect 36831 29469 36877 29507
rect 36831 29435 36837 29469
rect 36871 29435 36877 29469
rect 36831 29397 36877 29435
rect 36831 29363 36837 29397
rect 36871 29363 36877 29397
rect 36831 29325 36877 29363
rect 37405 29901 37815 29913
rect 37405 29363 37413 29901
rect 37807 29900 37815 29901
rect 38028 29900 38056 30008
rect 37807 29872 38056 29900
rect 39413 29901 39823 29913
rect 37807 29363 37815 29872
rect 37405 29351 37815 29363
rect 39413 29363 39420 29901
rect 39814 29363 39823 29901
rect 39868 29900 39896 30008
rect 40034 29900 40040 29912
rect 39868 29872 40040 29900
rect 40034 29860 40040 29872
rect 40092 29900 40098 29912
rect 40149 29901 40559 29913
rect 40149 29900 40157 29901
rect 40092 29872 40157 29900
rect 40092 29860 40098 29872
rect 39413 29351 39823 29363
rect 40149 29363 40157 29872
rect 40551 29363 40559 29901
rect 40149 29351 40559 29363
rect 42157 29901 42567 29913
rect 42157 29363 42164 29901
rect 42558 29363 42567 29901
rect 42157 29351 42567 29363
rect 36831 29291 36837 29325
rect 36871 29291 36877 29325
rect 36831 29253 36877 29291
rect 36831 29219 36837 29253
rect 36871 29219 36877 29253
rect 36831 29181 36877 29219
rect 36831 29147 36837 29181
rect 36871 29147 36877 29181
rect 36831 29109 36877 29147
rect 36831 29075 36837 29109
rect 36871 29075 36877 29109
rect 36831 29037 36877 29075
rect 36831 29003 36837 29037
rect 36871 29003 36877 29037
rect 36831 28965 36877 29003
rect 36831 28931 36837 28965
rect 36871 28931 36877 28965
rect 36831 28893 36877 28931
rect 36831 28859 36837 28893
rect 36871 28859 36877 28893
rect 36831 28821 36877 28859
rect 36831 28787 36837 28821
rect 36871 28787 36877 28821
rect 36831 28749 36877 28787
rect 36831 28715 36837 28749
rect 36871 28715 36877 28749
rect 36831 28677 36877 28715
rect 36831 28643 36837 28677
rect 36871 28643 36877 28677
rect 36831 28627 36877 28643
rect 37405 28948 37815 28953
rect 39298 28948 39304 28960
rect 37405 28941 39304 28948
rect 26568 28512 34100 28540
rect 26568 28500 26574 28512
rect 12526 28404 12532 28416
rect 12471 28376 12532 28404
rect 12526 28364 12532 28376
rect 12584 28364 12590 28416
rect 14182 28404 14188 28416
rect 14127 28376 14188 28404
rect 14182 28364 14188 28376
rect 14240 28364 14246 28416
rect 23382 28404 23388 28416
rect 23327 28376 23388 28404
rect 23382 28364 23388 28376
rect 23440 28364 23446 28416
rect 34072 28413 34100 28512
rect 34057 28407 34115 28413
rect 34057 28373 34069 28407
rect 34103 28373 34115 28407
rect 37405 28403 37413 28941
rect 37807 28920 39304 28941
rect 37807 28403 37815 28920
rect 39298 28908 39304 28920
rect 39356 28908 39362 28960
rect 39402 28941 39834 29351
rect 37405 28391 37815 28403
rect 39402 28403 39420 28941
rect 39814 28403 39834 28941
rect 40149 28941 40559 28953
rect 40034 28432 40040 28484
rect 40092 28472 40098 28484
rect 40149 28472 40157 28941
rect 40092 28444 40157 28472
rect 40092 28432 40098 28444
rect 39402 28387 39834 28403
rect 40149 28403 40157 28444
rect 40551 28403 40559 28941
rect 40149 28391 40559 28403
rect 42146 28941 42578 29351
rect 42146 28403 42164 28941
rect 42558 28403 42578 28941
rect 42146 28387 42578 28403
rect 34057 28367 34115 28373
rect 900 28330 47736 28332
rect 900 28214 922 28330
rect 2510 28289 46126 28330
rect 2510 28255 6197 28289
rect 6231 28255 6597 28289
rect 6631 28255 6997 28289
rect 7031 28255 7397 28289
rect 7431 28255 7797 28289
rect 7831 28255 8197 28289
rect 8231 28255 8597 28289
rect 8631 28255 8997 28289
rect 9031 28255 9397 28289
rect 9431 28255 9797 28289
rect 9831 28255 10197 28289
rect 10231 28255 10597 28289
rect 10631 28255 10997 28289
rect 11031 28255 11397 28289
rect 11431 28255 11797 28289
rect 11831 28255 12197 28289
rect 12231 28255 12597 28289
rect 12631 28255 12997 28289
rect 13031 28255 13397 28289
rect 13431 28255 13797 28289
rect 13831 28255 14197 28289
rect 14231 28255 14597 28289
rect 14631 28255 14997 28289
rect 15031 28255 15397 28289
rect 15431 28255 15797 28289
rect 15831 28255 16197 28289
rect 16231 28255 16597 28289
rect 16631 28255 16997 28289
rect 17031 28255 17397 28289
rect 17431 28255 17797 28289
rect 17831 28255 18197 28289
rect 18231 28255 18597 28289
rect 18631 28255 18997 28289
rect 19031 28255 19397 28289
rect 19431 28255 19797 28289
rect 19831 28255 20197 28289
rect 20231 28255 20597 28289
rect 20631 28255 20997 28289
rect 21031 28255 21397 28289
rect 21431 28255 21797 28289
rect 21831 28255 22197 28289
rect 22231 28255 22597 28289
rect 22631 28255 22997 28289
rect 23031 28255 23397 28289
rect 23431 28255 23797 28289
rect 23831 28255 24197 28289
rect 24231 28255 24597 28289
rect 24631 28255 24997 28289
rect 25031 28255 25397 28289
rect 25431 28255 25797 28289
rect 25831 28255 26197 28289
rect 26231 28255 26597 28289
rect 26631 28255 26997 28289
rect 27031 28255 27397 28289
rect 27431 28255 27797 28289
rect 27831 28255 28197 28289
rect 28231 28255 28597 28289
rect 28631 28255 28997 28289
rect 29031 28255 29397 28289
rect 29431 28255 29797 28289
rect 29831 28255 30197 28289
rect 30231 28255 30597 28289
rect 30631 28255 30997 28289
rect 31031 28255 31397 28289
rect 31431 28255 31797 28289
rect 31831 28255 32197 28289
rect 32231 28255 32597 28289
rect 32631 28255 32997 28289
rect 33031 28255 33397 28289
rect 33431 28255 34225 28289
rect 34259 28255 34625 28289
rect 34659 28255 35025 28289
rect 35059 28255 35425 28289
rect 35459 28255 35825 28289
rect 35859 28255 36225 28289
rect 36259 28255 36625 28289
rect 36659 28255 37577 28289
rect 37611 28255 37777 28289
rect 37811 28255 37977 28289
rect 38011 28255 38177 28289
rect 38211 28255 38377 28289
rect 38411 28255 38577 28289
rect 38611 28255 38777 28289
rect 38811 28255 38977 28289
rect 39011 28255 39177 28289
rect 39211 28255 39377 28289
rect 39411 28255 39577 28289
rect 39611 28255 40321 28289
rect 40355 28255 40521 28289
rect 40555 28255 40721 28289
rect 40755 28255 40921 28289
rect 40955 28255 41121 28289
rect 41155 28255 41321 28289
rect 41355 28255 41521 28289
rect 41555 28255 41721 28289
rect 41755 28255 41921 28289
rect 41955 28255 42121 28289
rect 42155 28255 42321 28289
rect 42355 28255 46126 28289
rect 2510 28214 46126 28255
rect 47714 28214 47736 28330
rect 900 28212 47736 28214
rect 3348 26450 45288 26452
rect 3348 26334 3370 26450
rect 4958 26409 43678 26450
rect 4958 26375 6903 26409
rect 6937 26375 7103 26409
rect 7137 26375 7303 26409
rect 7337 26375 7503 26409
rect 7537 26375 7703 26409
rect 7737 26375 7903 26409
rect 7937 26375 8103 26409
rect 8137 26375 8303 26409
rect 8337 26375 8503 26409
rect 8537 26375 8703 26409
rect 8737 26375 8903 26409
rect 8937 26375 9725 26409
rect 9759 26375 10125 26409
rect 10159 26375 10525 26409
rect 10559 26375 10925 26409
rect 10959 26375 11325 26409
rect 11359 26375 11725 26409
rect 11759 26375 12125 26409
rect 12159 26375 12525 26409
rect 12559 26375 12925 26409
rect 12959 26375 13325 26409
rect 13359 26375 13725 26409
rect 13759 26375 14125 26409
rect 14159 26375 14525 26409
rect 14559 26375 14925 26409
rect 14959 26375 15607 26409
rect 15641 26375 16007 26409
rect 16041 26375 16407 26409
rect 16441 26375 16807 26409
rect 16841 26375 17207 26409
rect 17241 26375 17607 26409
rect 17641 26375 18007 26409
rect 18041 26375 18407 26409
rect 18441 26375 18807 26409
rect 18841 26375 19207 26409
rect 19241 26375 19607 26409
rect 19641 26375 20007 26409
rect 20041 26375 20407 26409
rect 20441 26375 20807 26409
rect 20841 26375 21207 26409
rect 21241 26375 21607 26409
rect 21641 26375 22007 26409
rect 22041 26375 22407 26409
rect 22441 26375 23151 26409
rect 23185 26375 23551 26409
rect 23585 26375 23951 26409
rect 23985 26375 24351 26409
rect 24385 26375 24751 26409
rect 24785 26375 25151 26409
rect 25185 26375 25551 26409
rect 25585 26375 25951 26409
rect 25985 26375 26351 26409
rect 26385 26375 26751 26409
rect 26785 26375 28443 26409
rect 28477 26375 28643 26409
rect 28677 26375 28843 26409
rect 28877 26375 29043 26409
rect 29077 26375 29243 26409
rect 29277 26375 29443 26409
rect 29477 26375 29643 26409
rect 29677 26375 29843 26409
rect 29877 26375 30043 26409
rect 30077 26375 30243 26409
rect 30277 26375 30443 26409
rect 30477 26375 30643 26409
rect 30677 26375 30843 26409
rect 30877 26375 31043 26409
rect 31077 26375 31243 26409
rect 31277 26375 31443 26409
rect 31477 26375 31643 26409
rect 31677 26375 31843 26409
rect 31877 26375 32043 26409
rect 32077 26375 32243 26409
rect 32277 26375 32443 26409
rect 32477 26375 32643 26409
rect 32677 26375 32843 26409
rect 32877 26375 33043 26409
rect 33077 26375 33243 26409
rect 33277 26375 33443 26409
rect 33477 26375 33643 26409
rect 33677 26375 33843 26409
rect 33877 26375 34043 26409
rect 34077 26375 34243 26409
rect 34277 26375 34443 26409
rect 34477 26375 34643 26409
rect 34677 26375 34843 26409
rect 34877 26375 35043 26409
rect 35077 26375 35243 26409
rect 35277 26375 35443 26409
rect 35477 26375 35643 26409
rect 35677 26375 35843 26409
rect 35877 26375 36043 26409
rect 36077 26375 36243 26409
rect 36277 26375 36443 26409
rect 36477 26375 36643 26409
rect 36677 26375 36843 26409
rect 36877 26375 37043 26409
rect 37077 26375 37243 26409
rect 37277 26375 37443 26409
rect 37477 26375 37643 26409
rect 37677 26375 37843 26409
rect 37877 26375 38043 26409
rect 38077 26375 38243 26409
rect 38277 26375 38443 26409
rect 38477 26375 38643 26409
rect 38677 26375 38843 26409
rect 38877 26375 39929 26409
rect 39963 26375 40129 26409
rect 40163 26375 40329 26409
rect 40363 26375 40529 26409
rect 40563 26375 40729 26409
rect 40763 26375 40929 26409
rect 40963 26375 41129 26409
rect 41163 26375 41329 26409
rect 41363 26375 41529 26409
rect 41563 26375 41729 26409
rect 41763 26375 41929 26409
rect 41963 26375 43678 26409
rect 4958 26334 43678 26375
rect 45266 26334 45288 26450
rect 3348 26332 45288 26334
rect 6731 26141 7141 26153
rect 6731 25603 6739 26141
rect 7133 25628 7141 26141
rect 8739 26141 9149 26153
rect 6731 25591 7104 25603
rect 7098 25576 7104 25591
rect 7156 25576 7162 25628
rect 8739 25603 8746 26141
rect 9140 25603 9149 26141
rect 9582 26120 9588 26172
rect 9640 26120 9646 26172
rect 8739 25591 9149 25603
rect 9583 26107 9589 26120
rect 9623 26107 9629 26120
rect 9583 26069 9629 26107
rect 9583 26035 9589 26069
rect 9623 26035 9629 26069
rect 9968 26092 9996 26332
rect 26145 26231 26203 26237
rect 26145 26197 26157 26231
rect 26191 26228 26203 26231
rect 26234 26228 26240 26240
rect 26191 26200 26240 26228
rect 26191 26197 26203 26200
rect 26145 26191 26203 26197
rect 26234 26188 26240 26200
rect 26292 26188 26298 26240
rect 10041 26141 10087 26157
rect 10041 26107 10047 26141
rect 10081 26107 10087 26141
rect 10041 26092 10087 26107
rect 9968 26069 10087 26092
rect 9968 26064 10047 26069
rect 9583 25997 9629 26035
rect 9583 25963 9589 25997
rect 9623 25963 9629 25997
rect 9583 25925 9629 25963
rect 9583 25891 9589 25925
rect 9623 25891 9629 25925
rect 9583 25853 9629 25891
rect 9583 25819 9589 25853
rect 9623 25819 9629 25853
rect 9583 25781 9629 25819
rect 9583 25747 9589 25781
rect 9623 25747 9629 25781
rect 9583 25709 9629 25747
rect 9583 25675 9589 25709
rect 9623 25675 9629 25709
rect 9583 25637 9629 25675
rect 9583 25603 9589 25637
rect 9623 25603 9629 25637
rect 6731 25181 7141 25193
rect 6731 24643 6739 25181
rect 7133 24664 7141 25181
rect 8728 25181 9160 25591
rect 7190 24664 7196 24676
rect 7133 24643 7196 24664
rect 6731 24636 7196 24643
rect 6731 24631 7141 24636
rect 7190 24624 7196 24636
rect 7248 24624 7254 24676
rect 8728 24643 8746 25181
rect 9140 24643 9160 25181
rect 9583 25565 9629 25603
rect 9583 25531 9589 25565
rect 9623 25531 9629 25565
rect 9583 25493 9629 25531
rect 9583 25459 9589 25493
rect 9623 25459 9629 25493
rect 9583 25421 9629 25459
rect 9583 25387 9589 25421
rect 9623 25387 9629 25421
rect 9583 25349 9629 25387
rect 9583 25315 9589 25349
rect 9623 25315 9629 25349
rect 9583 25277 9629 25315
rect 9583 25243 9589 25277
rect 9623 25243 9629 25277
rect 9583 25205 9629 25243
rect 9583 25171 9589 25205
rect 9623 25171 9629 25205
rect 9583 25133 9629 25171
rect 9583 25099 9589 25133
rect 9623 25099 9629 25133
rect 9583 25061 9629 25099
rect 9583 25027 9589 25061
rect 9623 25027 9629 25061
rect 9583 24989 9629 25027
rect 9583 24955 9589 24989
rect 9623 24955 9629 24989
rect 9583 24917 9629 24955
rect 9583 24883 9589 24917
rect 9623 24883 9629 24917
rect 9583 24867 9629 24883
rect 10041 26035 10047 26064
rect 10081 26035 10087 26069
rect 10041 25997 10087 26035
rect 10041 25963 10047 25997
rect 10081 25963 10087 25997
rect 10041 25925 10087 25963
rect 10041 25891 10047 25925
rect 10081 25891 10087 25925
rect 10041 25853 10087 25891
rect 10041 25819 10047 25853
rect 10081 25819 10087 25853
rect 10041 25781 10087 25819
rect 10041 25747 10047 25781
rect 10081 25747 10087 25781
rect 10041 25709 10087 25747
rect 10041 25675 10047 25709
rect 10081 25675 10087 25709
rect 10041 25637 10087 25675
rect 10041 25603 10047 25637
rect 10081 25603 10087 25637
rect 10041 25565 10087 25603
rect 10041 25531 10047 25565
rect 10081 25531 10087 25565
rect 10041 25493 10087 25531
rect 10041 25459 10047 25493
rect 10081 25459 10087 25493
rect 10041 25421 10087 25459
rect 10041 25387 10047 25421
rect 10081 25387 10087 25421
rect 10041 25349 10087 25387
rect 10041 25315 10047 25349
rect 10081 25315 10087 25349
rect 10041 25277 10087 25315
rect 10041 25243 10047 25277
rect 10081 25243 10087 25277
rect 10041 25205 10087 25243
rect 10041 25171 10047 25205
rect 10081 25171 10087 25205
rect 10041 25133 10087 25171
rect 10041 25099 10047 25133
rect 10081 25099 10087 25133
rect 10041 25061 10087 25099
rect 10041 25027 10047 25061
rect 10081 25027 10087 25061
rect 10041 24989 10087 25027
rect 10041 24955 10047 24989
rect 10081 24955 10087 24989
rect 10041 24917 10087 24955
rect 10041 24883 10047 24917
rect 10081 24883 10087 24917
rect 10041 24867 10087 24883
rect 10499 26141 10545 26157
rect 10499 26107 10505 26141
rect 10539 26107 10545 26141
rect 10499 26069 10545 26107
rect 10499 26035 10505 26069
rect 10539 26035 10545 26069
rect 10499 25997 10545 26035
rect 10499 25963 10505 25997
rect 10539 25963 10545 25997
rect 10499 25925 10545 25963
rect 10499 25891 10505 25925
rect 10539 25891 10545 25925
rect 10499 25853 10545 25891
rect 10499 25819 10505 25853
rect 10539 25819 10545 25853
rect 10499 25781 10545 25819
rect 10499 25747 10505 25781
rect 10539 25747 10545 25781
rect 10499 25709 10545 25747
rect 10499 25675 10505 25709
rect 10539 25675 10545 25709
rect 10499 25637 10545 25675
rect 10499 25603 10505 25637
rect 10539 25603 10545 25637
rect 10499 25565 10545 25603
rect 10499 25531 10505 25565
rect 10539 25531 10545 25565
rect 10499 25493 10545 25531
rect 10499 25459 10505 25493
rect 10539 25459 10545 25493
rect 10499 25421 10545 25459
rect 10499 25387 10505 25421
rect 10539 25387 10545 25421
rect 10499 25349 10545 25387
rect 10499 25315 10505 25349
rect 10539 25315 10545 25349
rect 10499 25277 10545 25315
rect 10499 25243 10505 25277
rect 10539 25243 10545 25277
rect 10499 25205 10545 25243
rect 10499 25171 10505 25205
rect 10539 25171 10545 25205
rect 10499 25133 10545 25171
rect 10499 25099 10505 25133
rect 10539 25099 10545 25133
rect 10499 25061 10545 25099
rect 10499 25027 10505 25061
rect 10539 25027 10545 25061
rect 10499 24989 10545 25027
rect 10499 24955 10505 24989
rect 10539 24955 10545 24989
rect 10499 24917 10545 24955
rect 10499 24883 10505 24917
rect 10539 24883 10545 24917
rect 10499 24867 10545 24883
rect 10957 26141 11003 26157
rect 10957 26107 10963 26141
rect 10997 26107 11003 26141
rect 10957 26069 11003 26107
rect 10957 26035 10963 26069
rect 10997 26035 11003 26069
rect 10957 25997 11003 26035
rect 10957 25963 10963 25997
rect 10997 25963 11003 25997
rect 10957 25925 11003 25963
rect 10957 25891 10963 25925
rect 10997 25891 11003 25925
rect 10957 25853 11003 25891
rect 10957 25819 10963 25853
rect 10997 25819 11003 25853
rect 10957 25781 11003 25819
rect 10957 25747 10963 25781
rect 10997 25747 11003 25781
rect 10957 25709 11003 25747
rect 10957 25675 10963 25709
rect 10997 25675 11003 25709
rect 10957 25637 11003 25675
rect 10957 25603 10963 25637
rect 10997 25603 11003 25637
rect 10957 25565 11003 25603
rect 10957 25531 10963 25565
rect 10997 25531 11003 25565
rect 10957 25493 11003 25531
rect 10957 25459 10963 25493
rect 10997 25459 11003 25493
rect 10957 25421 11003 25459
rect 10957 25387 10963 25421
rect 10997 25387 11003 25421
rect 10957 25349 11003 25387
rect 10957 25315 10963 25349
rect 10997 25315 11003 25349
rect 10957 25277 11003 25315
rect 10957 25243 10963 25277
rect 10997 25243 11003 25277
rect 10957 25205 11003 25243
rect 10957 25171 10963 25205
rect 10997 25171 11003 25205
rect 10957 25133 11003 25171
rect 10957 25099 10963 25133
rect 10997 25099 11003 25133
rect 10957 25061 11003 25099
rect 10957 25027 10963 25061
rect 10997 25027 11003 25061
rect 10957 24989 11003 25027
rect 10957 24955 10963 24989
rect 10997 24955 11003 24989
rect 10957 24917 11003 24955
rect 10957 24883 10963 24917
rect 10997 24883 11003 24917
rect 10957 24867 11003 24883
rect 11415 26141 11461 26157
rect 11415 26107 11421 26141
rect 11455 26107 11461 26141
rect 11415 26069 11461 26107
rect 11415 26035 11421 26069
rect 11455 26035 11461 26069
rect 11415 25997 11461 26035
rect 11415 25963 11421 25997
rect 11455 25963 11461 25997
rect 11415 25925 11461 25963
rect 11415 25891 11421 25925
rect 11455 25891 11461 25925
rect 11415 25853 11461 25891
rect 11415 25819 11421 25853
rect 11455 25819 11461 25853
rect 11415 25781 11461 25819
rect 11415 25747 11421 25781
rect 11455 25747 11461 25781
rect 11415 25709 11461 25747
rect 11415 25675 11421 25709
rect 11455 25675 11461 25709
rect 11415 25637 11461 25675
rect 11415 25603 11421 25637
rect 11455 25603 11461 25637
rect 11415 25565 11461 25603
rect 11415 25531 11421 25565
rect 11455 25531 11461 25565
rect 11415 25493 11461 25531
rect 11415 25459 11421 25493
rect 11455 25459 11461 25493
rect 11415 25421 11461 25459
rect 11415 25387 11421 25421
rect 11455 25387 11461 25421
rect 11415 25349 11461 25387
rect 11415 25315 11421 25349
rect 11455 25315 11461 25349
rect 11415 25277 11461 25315
rect 11415 25243 11421 25277
rect 11455 25243 11461 25277
rect 11415 25205 11461 25243
rect 11415 25171 11421 25205
rect 11455 25171 11461 25205
rect 11415 25133 11461 25171
rect 11415 25099 11421 25133
rect 11455 25099 11461 25133
rect 11415 25061 11461 25099
rect 11415 25027 11421 25061
rect 11455 25027 11461 25061
rect 11415 24989 11461 25027
rect 11415 24955 11421 24989
rect 11455 24955 11461 24989
rect 11415 24917 11461 24955
rect 11415 24883 11421 24917
rect 11455 24883 11461 24917
rect 11415 24867 11461 24883
rect 11873 26141 11919 26157
rect 11873 26107 11879 26141
rect 11913 26107 11919 26141
rect 11873 26069 11919 26107
rect 11873 26035 11879 26069
rect 11913 26035 11919 26069
rect 11873 25997 11919 26035
rect 11873 25963 11879 25997
rect 11913 25963 11919 25997
rect 11873 25925 11919 25963
rect 11873 25891 11879 25925
rect 11913 25891 11919 25925
rect 11873 25853 11919 25891
rect 11873 25819 11879 25853
rect 11913 25819 11919 25853
rect 11873 25781 11919 25819
rect 11873 25747 11879 25781
rect 11913 25747 11919 25781
rect 11873 25709 11919 25747
rect 11873 25675 11879 25709
rect 11913 25675 11919 25709
rect 11873 25637 11919 25675
rect 11873 25603 11879 25637
rect 11913 25603 11919 25637
rect 11873 25565 11919 25603
rect 11873 25531 11879 25565
rect 11913 25531 11919 25565
rect 11873 25493 11919 25531
rect 11873 25459 11879 25493
rect 11913 25459 11919 25493
rect 11873 25421 11919 25459
rect 11873 25387 11879 25421
rect 11913 25387 11919 25421
rect 11873 25349 11919 25387
rect 11873 25315 11879 25349
rect 11913 25315 11919 25349
rect 11873 25277 11919 25315
rect 11873 25243 11879 25277
rect 11913 25243 11919 25277
rect 11873 25205 11919 25243
rect 11873 25171 11879 25205
rect 11913 25171 11919 25205
rect 11873 25133 11919 25171
rect 11873 25099 11879 25133
rect 11913 25099 11919 25133
rect 11873 25061 11919 25099
rect 11873 25027 11879 25061
rect 11913 25027 11919 25061
rect 11873 24989 11919 25027
rect 11873 24955 11879 24989
rect 11913 24955 11919 24989
rect 11873 24917 11919 24955
rect 11873 24883 11879 24917
rect 11913 24883 11919 24917
rect 11873 24867 11919 24883
rect 12331 26141 12377 26157
rect 12331 26107 12337 26141
rect 12371 26107 12377 26141
rect 12331 26069 12377 26107
rect 12331 26035 12337 26069
rect 12371 26035 12377 26069
rect 12331 25997 12377 26035
rect 12331 25963 12337 25997
rect 12371 25963 12377 25997
rect 12331 25925 12377 25963
rect 12331 25891 12337 25925
rect 12371 25891 12377 25925
rect 12331 25853 12377 25891
rect 12331 25819 12337 25853
rect 12371 25819 12377 25853
rect 12331 25781 12377 25819
rect 12331 25747 12337 25781
rect 12371 25747 12377 25781
rect 12331 25709 12377 25747
rect 12331 25675 12337 25709
rect 12371 25675 12377 25709
rect 12331 25637 12377 25675
rect 12331 25603 12337 25637
rect 12371 25603 12377 25637
rect 12331 25565 12377 25603
rect 12331 25531 12337 25565
rect 12371 25531 12377 25565
rect 12331 25493 12377 25531
rect 12331 25459 12337 25493
rect 12371 25459 12377 25493
rect 12331 25421 12377 25459
rect 12331 25387 12337 25421
rect 12371 25387 12377 25421
rect 12331 25349 12377 25387
rect 12331 25315 12337 25349
rect 12371 25315 12377 25349
rect 12331 25277 12377 25315
rect 12331 25243 12337 25277
rect 12371 25243 12377 25277
rect 12331 25205 12377 25243
rect 12331 25171 12337 25205
rect 12371 25171 12377 25205
rect 12331 25133 12377 25171
rect 12331 25099 12337 25133
rect 12371 25099 12377 25133
rect 12331 25061 12377 25099
rect 12331 25027 12337 25061
rect 12371 25027 12377 25061
rect 12331 24989 12377 25027
rect 12331 24955 12337 24989
rect 12371 24955 12377 24989
rect 12331 24917 12377 24955
rect 12331 24883 12337 24917
rect 12371 24883 12377 24917
rect 12331 24867 12377 24883
rect 12789 26141 12835 26157
rect 12789 26107 12795 26141
rect 12829 26107 12835 26141
rect 12789 26069 12835 26107
rect 12789 26035 12795 26069
rect 12829 26035 12835 26069
rect 12789 25997 12835 26035
rect 12789 25963 12795 25997
rect 12829 25963 12835 25997
rect 12789 25925 12835 25963
rect 12789 25891 12795 25925
rect 12829 25891 12835 25925
rect 12789 25853 12835 25891
rect 12789 25819 12795 25853
rect 12829 25819 12835 25853
rect 12789 25781 12835 25819
rect 12789 25747 12795 25781
rect 12829 25747 12835 25781
rect 12789 25709 12835 25747
rect 12789 25675 12795 25709
rect 12829 25675 12835 25709
rect 12789 25637 12835 25675
rect 12789 25603 12795 25637
rect 12829 25603 12835 25637
rect 12789 25565 12835 25603
rect 12789 25531 12795 25565
rect 12829 25531 12835 25565
rect 12789 25493 12835 25531
rect 12789 25459 12795 25493
rect 12829 25459 12835 25493
rect 12789 25421 12835 25459
rect 12789 25387 12795 25421
rect 12829 25387 12835 25421
rect 12789 25349 12835 25387
rect 12789 25315 12795 25349
rect 12829 25315 12835 25349
rect 12789 25277 12835 25315
rect 12789 25243 12795 25277
rect 12829 25243 12835 25277
rect 12789 25205 12835 25243
rect 12789 25171 12795 25205
rect 12829 25171 12835 25205
rect 12789 25133 12835 25171
rect 12789 25099 12795 25133
rect 12829 25099 12835 25133
rect 12789 25061 12835 25099
rect 12789 25027 12795 25061
rect 12829 25027 12835 25061
rect 12789 24989 12835 25027
rect 12789 24955 12795 24989
rect 12829 24955 12835 24989
rect 12789 24917 12835 24955
rect 12789 24883 12795 24917
rect 12829 24883 12835 24917
rect 12789 24867 12835 24883
rect 13247 26141 13293 26157
rect 13247 26107 13253 26141
rect 13287 26107 13293 26141
rect 13247 26069 13293 26107
rect 13247 26035 13253 26069
rect 13287 26035 13293 26069
rect 13247 25997 13293 26035
rect 13247 25963 13253 25997
rect 13287 25963 13293 25997
rect 13247 25925 13293 25963
rect 13247 25891 13253 25925
rect 13287 25891 13293 25925
rect 13247 25853 13293 25891
rect 13247 25819 13253 25853
rect 13287 25819 13293 25853
rect 13247 25781 13293 25819
rect 13247 25747 13253 25781
rect 13287 25747 13293 25781
rect 13247 25709 13293 25747
rect 13247 25675 13253 25709
rect 13287 25675 13293 25709
rect 13247 25637 13293 25675
rect 13247 25603 13253 25637
rect 13287 25603 13293 25637
rect 13247 25565 13293 25603
rect 13247 25531 13253 25565
rect 13287 25531 13293 25565
rect 13247 25493 13293 25531
rect 13247 25459 13253 25493
rect 13287 25459 13293 25493
rect 13247 25421 13293 25459
rect 13247 25387 13253 25421
rect 13287 25387 13293 25421
rect 13247 25349 13293 25387
rect 13247 25315 13253 25349
rect 13287 25315 13293 25349
rect 13247 25277 13293 25315
rect 13247 25243 13253 25277
rect 13287 25243 13293 25277
rect 13247 25205 13293 25243
rect 13247 25171 13253 25205
rect 13287 25171 13293 25205
rect 13247 25133 13293 25171
rect 13247 25099 13253 25133
rect 13287 25099 13293 25133
rect 13247 25061 13293 25099
rect 13247 25027 13253 25061
rect 13287 25027 13293 25061
rect 13247 24989 13293 25027
rect 13247 24955 13253 24989
rect 13287 24955 13293 24989
rect 13247 24917 13293 24955
rect 13247 24883 13253 24917
rect 13287 24883 13293 24917
rect 13247 24867 13293 24883
rect 13705 26141 13751 26157
rect 13705 26107 13711 26141
rect 13745 26107 13751 26141
rect 13705 26069 13751 26107
rect 13705 26035 13711 26069
rect 13745 26035 13751 26069
rect 13705 25997 13751 26035
rect 13705 25963 13711 25997
rect 13745 25963 13751 25997
rect 13705 25925 13751 25963
rect 13705 25891 13711 25925
rect 13745 25891 13751 25925
rect 13705 25853 13751 25891
rect 13705 25819 13711 25853
rect 13745 25819 13751 25853
rect 13705 25781 13751 25819
rect 13705 25747 13711 25781
rect 13745 25747 13751 25781
rect 13705 25709 13751 25747
rect 13705 25675 13711 25709
rect 13745 25675 13751 25709
rect 13705 25637 13751 25675
rect 13705 25603 13711 25637
rect 13745 25603 13751 25637
rect 13705 25565 13751 25603
rect 13705 25531 13711 25565
rect 13745 25531 13751 25565
rect 13705 25493 13751 25531
rect 13705 25459 13711 25493
rect 13745 25459 13751 25493
rect 13705 25421 13751 25459
rect 13705 25387 13711 25421
rect 13745 25387 13751 25421
rect 13705 25349 13751 25387
rect 13705 25315 13711 25349
rect 13745 25315 13751 25349
rect 13705 25277 13751 25315
rect 13705 25243 13711 25277
rect 13745 25243 13751 25277
rect 13705 25205 13751 25243
rect 13705 25171 13711 25205
rect 13745 25171 13751 25205
rect 13705 25133 13751 25171
rect 13705 25099 13711 25133
rect 13745 25099 13751 25133
rect 13705 25061 13751 25099
rect 13705 25027 13711 25061
rect 13745 25027 13751 25061
rect 13705 24989 13751 25027
rect 13705 24955 13711 24989
rect 13745 24955 13751 24989
rect 13705 24917 13751 24955
rect 13705 24883 13711 24917
rect 13745 24883 13751 24917
rect 13705 24867 13751 24883
rect 14163 26141 14209 26157
rect 14163 26107 14169 26141
rect 14203 26107 14209 26141
rect 14163 26069 14209 26107
rect 14163 26035 14169 26069
rect 14203 26035 14209 26069
rect 14163 25997 14209 26035
rect 14163 25963 14169 25997
rect 14203 25963 14209 25997
rect 14163 25925 14209 25963
rect 14163 25891 14169 25925
rect 14203 25891 14209 25925
rect 14163 25853 14209 25891
rect 14163 25819 14169 25853
rect 14203 25819 14209 25853
rect 14163 25781 14209 25819
rect 14163 25747 14169 25781
rect 14203 25747 14209 25781
rect 14163 25709 14209 25747
rect 14163 25675 14169 25709
rect 14203 25675 14209 25709
rect 14163 25637 14209 25675
rect 14163 25603 14169 25637
rect 14203 25603 14209 25637
rect 14163 25565 14209 25603
rect 14163 25531 14169 25565
rect 14203 25531 14209 25565
rect 14163 25493 14209 25531
rect 14163 25459 14169 25493
rect 14203 25459 14209 25493
rect 14163 25421 14209 25459
rect 14163 25387 14169 25421
rect 14203 25387 14209 25421
rect 14163 25349 14209 25387
rect 14163 25315 14169 25349
rect 14203 25315 14209 25349
rect 14163 25277 14209 25315
rect 14163 25243 14169 25277
rect 14203 25243 14209 25277
rect 14163 25205 14209 25243
rect 14163 25171 14169 25205
rect 14203 25171 14209 25205
rect 14163 25133 14209 25171
rect 14163 25099 14169 25133
rect 14203 25099 14209 25133
rect 14163 25061 14209 25099
rect 14163 25027 14169 25061
rect 14203 25027 14209 25061
rect 14163 24989 14209 25027
rect 14163 24955 14169 24989
rect 14203 24955 14209 24989
rect 14163 24917 14209 24955
rect 14163 24883 14169 24917
rect 14203 24883 14209 24917
rect 14163 24867 14209 24883
rect 14621 26141 14667 26157
rect 14621 26107 14627 26141
rect 14661 26107 14667 26141
rect 14621 26069 14667 26107
rect 14621 26035 14627 26069
rect 14661 26035 14667 26069
rect 14621 25997 14667 26035
rect 14621 25963 14627 25997
rect 14661 25963 14667 25997
rect 14621 25925 14667 25963
rect 14621 25891 14627 25925
rect 14661 25891 14667 25925
rect 14621 25853 14667 25891
rect 14621 25819 14627 25853
rect 14661 25819 14667 25853
rect 14621 25781 14667 25819
rect 14621 25747 14627 25781
rect 14661 25747 14667 25781
rect 14621 25709 14667 25747
rect 14621 25675 14627 25709
rect 14661 25675 14667 25709
rect 14621 25637 14667 25675
rect 14621 25603 14627 25637
rect 14661 25603 14667 25637
rect 14621 25565 14667 25603
rect 14621 25531 14627 25565
rect 14661 25531 14667 25565
rect 14621 25493 14667 25531
rect 14621 25459 14627 25493
rect 14661 25459 14667 25493
rect 14621 25421 14667 25459
rect 14621 25387 14627 25421
rect 14661 25387 14667 25421
rect 14621 25349 14667 25387
rect 14621 25315 14627 25349
rect 14661 25315 14667 25349
rect 14621 25277 14667 25315
rect 14621 25243 14627 25277
rect 14661 25243 14667 25277
rect 14621 25205 14667 25243
rect 14621 25171 14627 25205
rect 14661 25171 14667 25205
rect 14621 25133 14667 25171
rect 14621 25099 14627 25133
rect 14661 25099 14667 25133
rect 14621 25061 14667 25099
rect 14621 25027 14627 25061
rect 14661 25027 14667 25061
rect 14621 24989 14667 25027
rect 14621 24955 14627 24989
rect 14661 24955 14667 24989
rect 14621 24917 14667 24955
rect 14621 24883 14627 24917
rect 14661 24883 14667 24917
rect 14621 24867 14667 24883
rect 15079 26141 15125 26157
rect 15079 26107 15085 26141
rect 15119 26107 15125 26141
rect 15079 26069 15125 26107
rect 39757 26141 40167 26153
rect 15079 26035 15085 26069
rect 15119 26035 15125 26069
rect 15079 25997 15125 26035
rect 28286 26076 38954 26082
rect 28286 26042 28306 26076
rect 28340 26042 28396 26076
rect 28430 26042 28486 26076
rect 28520 26042 28576 26076
rect 28610 26042 28666 26076
rect 28700 26042 28756 26076
rect 28790 26042 28846 26076
rect 28880 26042 28936 26076
rect 28970 26042 29026 26076
rect 29060 26042 29116 26076
rect 29150 26042 29206 26076
rect 29240 26042 29296 26076
rect 29330 26042 29386 26076
rect 29420 26042 29476 26076
rect 29510 26042 29646 26076
rect 29680 26042 29736 26076
rect 29770 26042 29826 26076
rect 29860 26042 29916 26076
rect 29950 26042 30006 26076
rect 30040 26042 30096 26076
rect 30130 26042 30186 26076
rect 30220 26042 30276 26076
rect 30310 26042 30366 26076
rect 30400 26042 30456 26076
rect 30490 26042 30546 26076
rect 30580 26042 30636 26076
rect 30670 26042 30726 26076
rect 30760 26042 30816 26076
rect 30850 26042 30986 26076
rect 31020 26042 31076 26076
rect 31110 26042 31166 26076
rect 31200 26042 31256 26076
rect 31290 26042 31346 26076
rect 31380 26042 31436 26076
rect 31470 26042 31526 26076
rect 31560 26042 31616 26076
rect 31650 26042 31706 26076
rect 31740 26042 31796 26076
rect 31830 26042 31886 26076
rect 31920 26042 31976 26076
rect 32010 26042 32066 26076
rect 32100 26042 32156 26076
rect 32190 26042 32326 26076
rect 32360 26042 32416 26076
rect 32450 26042 32506 26076
rect 32540 26042 32596 26076
rect 32630 26042 32686 26076
rect 32720 26042 32776 26076
rect 32810 26042 32866 26076
rect 32900 26042 32956 26076
rect 32990 26042 33046 26076
rect 33080 26042 33136 26076
rect 33170 26042 33226 26076
rect 33260 26042 33316 26076
rect 33350 26042 33406 26076
rect 33440 26042 33496 26076
rect 33530 26042 33666 26076
rect 33700 26042 33756 26076
rect 33790 26042 33846 26076
rect 33880 26042 33936 26076
rect 33970 26042 34026 26076
rect 34060 26042 34116 26076
rect 34150 26042 34206 26076
rect 34240 26042 34296 26076
rect 34330 26042 34386 26076
rect 34420 26042 34476 26076
rect 34510 26042 34566 26076
rect 34600 26042 34656 26076
rect 34690 26042 34746 26076
rect 34780 26042 34836 26076
rect 34870 26042 35006 26076
rect 35040 26042 35096 26076
rect 35130 26042 35186 26076
rect 35220 26042 35276 26076
rect 35310 26042 35366 26076
rect 35400 26042 35456 26076
rect 35490 26042 35546 26076
rect 35580 26042 35636 26076
rect 35670 26042 35726 26076
rect 35760 26042 35816 26076
rect 35850 26042 35906 26076
rect 35940 26042 35996 26076
rect 36030 26042 36086 26076
rect 36120 26042 36176 26076
rect 36210 26042 36346 26076
rect 36380 26042 36436 26076
rect 36470 26042 36526 26076
rect 36560 26042 36616 26076
rect 36650 26042 36706 26076
rect 36740 26042 36796 26076
rect 36830 26042 36886 26076
rect 36920 26042 36976 26076
rect 37010 26042 37066 26076
rect 37100 26042 37156 26076
rect 37190 26042 37246 26076
rect 37280 26042 37336 26076
rect 37370 26042 37426 26076
rect 37460 26042 37516 26076
rect 37550 26042 37686 26076
rect 37720 26042 37776 26076
rect 37810 26042 37866 26076
rect 37900 26042 37956 26076
rect 37990 26042 38046 26076
rect 38080 26042 38136 26076
rect 38170 26042 38226 26076
rect 38260 26042 38316 26076
rect 38350 26042 38406 26076
rect 38440 26042 38496 26076
rect 38530 26042 38586 26076
rect 38620 26042 38676 26076
rect 38710 26042 38766 26076
rect 38800 26042 38856 26076
rect 38890 26042 38954 26076
rect 28286 26012 38954 26042
rect 15079 25963 15085 25997
rect 15119 25963 15125 25997
rect 15079 25925 15125 25963
rect 28460 25932 28488 26012
rect 15079 25891 15085 25925
rect 15119 25891 15125 25925
rect 28450 25916 38790 25932
rect 15079 25853 15125 25891
rect 15079 25819 15085 25853
rect 15119 25819 15125 25853
rect 15079 25781 15125 25819
rect 15079 25747 15085 25781
rect 15119 25747 15125 25781
rect 15079 25709 15125 25747
rect 15079 25675 15085 25709
rect 15119 25675 15125 25709
rect 15079 25637 15125 25675
rect 15079 25603 15085 25637
rect 15119 25603 15125 25637
rect 15079 25565 15125 25603
rect 15079 25531 15085 25565
rect 15119 25531 15125 25565
rect 15079 25493 15125 25531
rect 15079 25459 15085 25493
rect 15119 25459 15125 25493
rect 15079 25421 15125 25459
rect 15079 25387 15085 25421
rect 15119 25387 15125 25421
rect 15079 25349 15125 25387
rect 15079 25315 15085 25349
rect 15119 25315 15125 25349
rect 15079 25277 15125 25315
rect 15079 25243 15085 25277
rect 15119 25243 15125 25277
rect 15079 25205 15125 25243
rect 15079 25171 15085 25205
rect 15119 25171 15125 25205
rect 15079 25133 15125 25171
rect 15079 25099 15085 25133
rect 15119 25099 15125 25133
rect 22974 25889 23020 25912
rect 22974 25855 22980 25889
rect 23014 25855 23020 25889
rect 22974 25817 23020 25855
rect 22974 25783 22980 25817
rect 23014 25783 23020 25817
rect 22974 25745 23020 25783
rect 22974 25711 22980 25745
rect 23014 25711 23020 25745
rect 22974 25673 23020 25711
rect 22974 25639 22980 25673
rect 23014 25639 23020 25673
rect 22974 25601 23020 25639
rect 22974 25567 22980 25601
rect 23014 25567 23020 25601
rect 22974 25529 23020 25567
rect 22974 25495 22980 25529
rect 23014 25495 23020 25529
rect 22974 25457 23020 25495
rect 22974 25423 22980 25457
rect 23014 25423 23020 25457
rect 22974 25385 23020 25423
rect 22974 25351 22980 25385
rect 23014 25351 23020 25385
rect 22974 25313 23020 25351
rect 22974 25279 22980 25313
rect 23014 25279 23020 25313
rect 22974 25241 23020 25279
rect 22974 25207 22980 25241
rect 23014 25207 23020 25241
rect 22974 25169 23020 25207
rect 22974 25135 22980 25169
rect 23014 25135 23020 25169
rect 22974 25112 23020 25135
rect 23432 25889 23478 25912
rect 23432 25855 23438 25889
rect 23472 25855 23478 25889
rect 23432 25817 23478 25855
rect 23432 25783 23438 25817
rect 23472 25783 23478 25817
rect 23432 25745 23478 25783
rect 23432 25711 23438 25745
rect 23472 25711 23478 25745
rect 23432 25673 23478 25711
rect 23432 25639 23438 25673
rect 23472 25639 23478 25673
rect 23432 25601 23478 25639
rect 23432 25567 23438 25601
rect 23472 25567 23478 25601
rect 23432 25529 23478 25567
rect 23432 25495 23438 25529
rect 23472 25495 23478 25529
rect 23432 25457 23478 25495
rect 23432 25423 23438 25457
rect 23472 25423 23478 25457
rect 23432 25385 23478 25423
rect 23432 25351 23438 25385
rect 23472 25351 23478 25385
rect 23432 25313 23478 25351
rect 23432 25279 23438 25313
rect 23472 25279 23478 25313
rect 23432 25241 23478 25279
rect 23432 25207 23438 25241
rect 23472 25207 23478 25241
rect 23432 25169 23478 25207
rect 23432 25135 23438 25169
rect 23472 25135 23478 25169
rect 23432 25112 23478 25135
rect 23890 25889 23936 25912
rect 23890 25855 23896 25889
rect 23930 25855 23936 25889
rect 23890 25817 23936 25855
rect 23890 25783 23896 25817
rect 23930 25783 23936 25817
rect 23890 25745 23936 25783
rect 23890 25711 23896 25745
rect 23930 25711 23936 25745
rect 23890 25673 23936 25711
rect 23890 25639 23896 25673
rect 23930 25639 23936 25673
rect 23890 25601 23936 25639
rect 23890 25567 23896 25601
rect 23930 25567 23936 25601
rect 23890 25529 23936 25567
rect 23890 25495 23896 25529
rect 23930 25495 23936 25529
rect 23890 25457 23936 25495
rect 23890 25423 23896 25457
rect 23930 25423 23936 25457
rect 23890 25385 23936 25423
rect 23890 25351 23896 25385
rect 23930 25351 23936 25385
rect 23890 25313 23936 25351
rect 23890 25279 23896 25313
rect 23930 25279 23936 25313
rect 23890 25241 23936 25279
rect 23890 25207 23896 25241
rect 23930 25207 23936 25241
rect 23890 25169 23936 25207
rect 23890 25135 23896 25169
rect 23930 25135 23936 25169
rect 23890 25112 23936 25135
rect 24348 25889 24394 25912
rect 24348 25855 24354 25889
rect 24388 25855 24394 25889
rect 24348 25817 24394 25855
rect 24348 25783 24354 25817
rect 24388 25783 24394 25817
rect 24348 25745 24394 25783
rect 24348 25711 24354 25745
rect 24388 25711 24394 25745
rect 24348 25673 24394 25711
rect 24348 25639 24354 25673
rect 24388 25639 24394 25673
rect 24348 25601 24394 25639
rect 24348 25567 24354 25601
rect 24388 25567 24394 25601
rect 24348 25529 24394 25567
rect 24348 25495 24354 25529
rect 24388 25495 24394 25529
rect 24348 25457 24394 25495
rect 24348 25423 24354 25457
rect 24388 25423 24394 25457
rect 24348 25385 24394 25423
rect 24348 25351 24354 25385
rect 24388 25351 24394 25385
rect 24348 25313 24394 25351
rect 24348 25279 24354 25313
rect 24388 25279 24394 25313
rect 24348 25241 24394 25279
rect 24348 25207 24354 25241
rect 24388 25207 24394 25241
rect 24348 25169 24394 25207
rect 24348 25135 24354 25169
rect 24388 25135 24394 25169
rect 24348 25112 24394 25135
rect 24806 25889 24852 25912
rect 24806 25855 24812 25889
rect 24846 25855 24852 25889
rect 24806 25817 24852 25855
rect 24806 25783 24812 25817
rect 24846 25783 24852 25817
rect 24806 25745 24852 25783
rect 24806 25711 24812 25745
rect 24846 25711 24852 25745
rect 24806 25673 24852 25711
rect 24806 25639 24812 25673
rect 24846 25639 24852 25673
rect 24806 25601 24852 25639
rect 24806 25567 24812 25601
rect 24846 25567 24852 25601
rect 24806 25529 24852 25567
rect 24806 25495 24812 25529
rect 24846 25495 24852 25529
rect 24806 25457 24852 25495
rect 24806 25423 24812 25457
rect 24846 25423 24852 25457
rect 24806 25385 24852 25423
rect 24806 25351 24812 25385
rect 24846 25351 24852 25385
rect 24806 25313 24852 25351
rect 24806 25279 24812 25313
rect 24846 25279 24852 25313
rect 24806 25241 24852 25279
rect 24806 25207 24812 25241
rect 24846 25207 24852 25241
rect 24806 25169 24852 25207
rect 24806 25135 24812 25169
rect 24846 25135 24852 25169
rect 24806 25112 24852 25135
rect 25264 25889 25310 25912
rect 25264 25855 25270 25889
rect 25304 25855 25310 25889
rect 25264 25817 25310 25855
rect 25264 25783 25270 25817
rect 25304 25783 25310 25817
rect 25264 25745 25310 25783
rect 25264 25711 25270 25745
rect 25304 25711 25310 25745
rect 25264 25673 25310 25711
rect 25264 25639 25270 25673
rect 25304 25639 25310 25673
rect 25264 25601 25310 25639
rect 25264 25567 25270 25601
rect 25304 25567 25310 25601
rect 25264 25529 25310 25567
rect 25264 25495 25270 25529
rect 25304 25495 25310 25529
rect 25264 25457 25310 25495
rect 25264 25423 25270 25457
rect 25304 25423 25310 25457
rect 25264 25385 25310 25423
rect 25264 25351 25270 25385
rect 25304 25351 25310 25385
rect 25264 25313 25310 25351
rect 25264 25279 25270 25313
rect 25304 25279 25310 25313
rect 25264 25241 25310 25279
rect 25264 25207 25270 25241
rect 25304 25207 25310 25241
rect 25264 25169 25310 25207
rect 25264 25135 25270 25169
rect 25304 25135 25310 25169
rect 25264 25112 25310 25135
rect 25722 25889 25768 25912
rect 25722 25855 25728 25889
rect 25762 25855 25768 25889
rect 25722 25817 25768 25855
rect 25722 25783 25728 25817
rect 25762 25783 25768 25817
rect 25722 25745 25768 25783
rect 25722 25711 25728 25745
rect 25762 25711 25768 25745
rect 25722 25673 25768 25711
rect 25722 25639 25728 25673
rect 25762 25639 25768 25673
rect 25722 25601 25768 25639
rect 25722 25567 25728 25601
rect 25762 25567 25768 25601
rect 25722 25529 25768 25567
rect 25722 25495 25728 25529
rect 25762 25495 25768 25529
rect 25722 25457 25768 25495
rect 25722 25423 25728 25457
rect 25762 25423 25768 25457
rect 25722 25385 25768 25423
rect 25722 25351 25728 25385
rect 25762 25351 25768 25385
rect 25722 25313 25768 25351
rect 25722 25279 25728 25313
rect 25762 25279 25768 25313
rect 25722 25241 25768 25279
rect 25722 25207 25728 25241
rect 25762 25207 25768 25241
rect 25722 25169 25768 25207
rect 25722 25135 25728 25169
rect 25762 25135 25768 25169
rect 25722 25112 25768 25135
rect 26180 25889 26226 25912
rect 26180 25855 26186 25889
rect 26220 25855 26226 25889
rect 26180 25817 26226 25855
rect 26180 25783 26186 25817
rect 26220 25783 26226 25817
rect 26180 25745 26226 25783
rect 26180 25711 26186 25745
rect 26220 25711 26226 25745
rect 26180 25673 26226 25711
rect 26180 25639 26186 25673
rect 26220 25639 26226 25673
rect 26180 25601 26226 25639
rect 26180 25567 26186 25601
rect 26220 25567 26226 25601
rect 26180 25529 26226 25567
rect 26180 25495 26186 25529
rect 26220 25495 26226 25529
rect 26180 25457 26226 25495
rect 26180 25423 26186 25457
rect 26220 25423 26226 25457
rect 26180 25385 26226 25423
rect 26180 25351 26186 25385
rect 26220 25351 26226 25385
rect 26180 25313 26226 25351
rect 26180 25279 26186 25313
rect 26220 25279 26226 25313
rect 26180 25241 26226 25279
rect 26180 25207 26186 25241
rect 26220 25207 26226 25241
rect 26180 25169 26226 25207
rect 26180 25135 26186 25169
rect 26220 25135 26226 25169
rect 26180 25112 26226 25135
rect 26638 25889 26684 25912
rect 26638 25855 26644 25889
rect 26678 25855 26684 25889
rect 26638 25817 26684 25855
rect 26638 25783 26644 25817
rect 26678 25783 26684 25817
rect 26638 25745 26684 25783
rect 26638 25711 26644 25745
rect 26678 25711 26684 25745
rect 26638 25673 26684 25711
rect 26638 25639 26644 25673
rect 26678 25639 26684 25673
rect 26638 25601 26684 25639
rect 26638 25567 26644 25601
rect 26678 25567 26684 25601
rect 26638 25529 26684 25567
rect 26638 25495 26644 25529
rect 26678 25495 26684 25529
rect 26638 25457 26684 25495
rect 26638 25423 26644 25457
rect 26678 25423 26684 25457
rect 26638 25385 26684 25423
rect 26638 25351 26644 25385
rect 26678 25351 26684 25385
rect 26638 25313 26684 25351
rect 26638 25279 26644 25313
rect 26678 25279 26684 25313
rect 26638 25241 26684 25279
rect 26638 25207 26644 25241
rect 26678 25207 26684 25241
rect 26638 25169 26684 25207
rect 26638 25135 26644 25169
rect 26678 25135 26684 25169
rect 26638 25112 26684 25135
rect 27096 25889 27142 25912
rect 27096 25855 27102 25889
rect 27136 25855 27142 25889
rect 28450 25882 28470 25916
rect 28504 25882 28560 25916
rect 28594 25882 28650 25916
rect 28684 25882 28740 25916
rect 28774 25882 28830 25916
rect 28864 25882 28920 25916
rect 28954 25882 29010 25916
rect 29044 25882 29100 25916
rect 29134 25882 29190 25916
rect 29224 25882 29280 25916
rect 29314 25882 29370 25916
rect 29404 25882 29810 25916
rect 29844 25882 29900 25916
rect 29934 25882 29990 25916
rect 30024 25882 30080 25916
rect 30114 25882 30170 25916
rect 30204 25882 30260 25916
rect 30294 25882 30350 25916
rect 30384 25882 30440 25916
rect 30474 25882 30530 25916
rect 30564 25882 30620 25916
rect 30654 25882 30710 25916
rect 30744 25882 31150 25916
rect 31184 25882 31240 25916
rect 31274 25882 31330 25916
rect 31364 25882 31420 25916
rect 31454 25882 31510 25916
rect 31544 25882 31600 25916
rect 31634 25882 31690 25916
rect 31724 25882 31780 25916
rect 31814 25882 31870 25916
rect 31904 25882 31960 25916
rect 31994 25882 32050 25916
rect 32084 25882 32490 25916
rect 32524 25882 32580 25916
rect 32614 25882 32670 25916
rect 32704 25882 32760 25916
rect 32794 25882 32850 25916
rect 32884 25882 32940 25916
rect 32974 25882 33030 25916
rect 33064 25882 33120 25916
rect 33154 25882 33210 25916
rect 33244 25882 33300 25916
rect 33334 25882 33390 25916
rect 33424 25882 33830 25916
rect 33864 25882 33920 25916
rect 33954 25882 34010 25916
rect 34044 25882 34100 25916
rect 34134 25882 34190 25916
rect 34224 25882 34280 25916
rect 34314 25882 34370 25916
rect 34404 25882 34460 25916
rect 34494 25882 34550 25916
rect 34584 25882 34640 25916
rect 34674 25882 34730 25916
rect 34764 25882 35170 25916
rect 35204 25882 35260 25916
rect 35294 25882 35350 25916
rect 35384 25882 35440 25916
rect 35474 25882 35530 25916
rect 35564 25882 35620 25916
rect 35654 25882 35710 25916
rect 35744 25882 35800 25916
rect 35834 25882 35890 25916
rect 35924 25882 35980 25916
rect 36014 25882 36070 25916
rect 36104 25882 36510 25916
rect 36544 25882 36600 25916
rect 36634 25882 36690 25916
rect 36724 25882 36780 25916
rect 36814 25882 36870 25916
rect 36904 25882 36960 25916
rect 36994 25882 37050 25916
rect 37084 25882 37140 25916
rect 37174 25882 37230 25916
rect 37264 25882 37320 25916
rect 37354 25882 37410 25916
rect 37444 25882 37850 25916
rect 37884 25882 37940 25916
rect 37974 25882 38030 25916
rect 38064 25882 38120 25916
rect 38154 25882 38210 25916
rect 38244 25882 38300 25916
rect 38334 25882 38390 25916
rect 38424 25882 38480 25916
rect 38514 25882 38570 25916
rect 38604 25882 38660 25916
rect 38694 25882 38750 25916
rect 38784 25882 38790 25916
rect 28450 25862 38790 25882
rect 27096 25817 27142 25855
rect 27096 25783 27102 25817
rect 27136 25783 27142 25817
rect 27096 25745 27142 25783
rect 31662 25758 31668 25764
rect 27096 25711 27102 25745
rect 27136 25711 27142 25745
rect 27096 25673 27142 25711
rect 27096 25639 27102 25673
rect 27136 25639 27142 25673
rect 27096 25601 27142 25639
rect 27096 25567 27102 25601
rect 27136 25567 27142 25601
rect 27096 25529 27142 25567
rect 27096 25495 27102 25529
rect 27136 25495 27142 25529
rect 27096 25457 27142 25495
rect 27096 25423 27102 25457
rect 27136 25423 27142 25457
rect 27096 25385 27142 25423
rect 27096 25351 27102 25385
rect 27136 25351 27142 25385
rect 27096 25313 27142 25351
rect 27096 25279 27102 25313
rect 27136 25279 27142 25313
rect 27096 25241 27142 25279
rect 27096 25207 27102 25241
rect 27136 25207 27142 25241
rect 27096 25169 27142 25207
rect 27096 25135 27102 25169
rect 27136 25135 27142 25169
rect 28624 25712 31668 25758
rect 31720 25758 31726 25764
rect 31720 25712 38616 25758
rect 28624 25678 28656 25712
rect 28690 25678 28756 25712
rect 28790 25678 28856 25712
rect 28890 25678 28956 25712
rect 28990 25678 29056 25712
rect 29090 25678 29156 25712
rect 29190 25678 29996 25712
rect 30030 25678 30096 25712
rect 30130 25678 30196 25712
rect 30230 25678 30296 25712
rect 30330 25678 30396 25712
rect 30430 25678 30496 25712
rect 30530 25678 31336 25712
rect 31370 25678 31436 25712
rect 31470 25678 31536 25712
rect 31570 25678 31636 25712
rect 31670 25678 31736 25712
rect 31770 25678 31836 25712
rect 31870 25678 32676 25712
rect 32710 25678 32776 25712
rect 32810 25678 32876 25712
rect 32910 25678 32976 25712
rect 33010 25678 33076 25712
rect 33110 25678 33176 25712
rect 33210 25678 34016 25712
rect 34050 25678 34116 25712
rect 34150 25678 34216 25712
rect 34250 25678 34316 25712
rect 34350 25678 34416 25712
rect 34450 25678 34516 25712
rect 34550 25678 35356 25712
rect 35390 25678 35456 25712
rect 35490 25678 35556 25712
rect 35590 25678 35656 25712
rect 35690 25678 35756 25712
rect 35790 25678 35856 25712
rect 35890 25678 36696 25712
rect 36730 25678 36796 25712
rect 36830 25678 36896 25712
rect 36930 25678 36996 25712
rect 37030 25678 37096 25712
rect 37130 25678 37196 25712
rect 37230 25678 38036 25712
rect 38070 25678 38136 25712
rect 38170 25678 38236 25712
rect 38270 25678 38336 25712
rect 38370 25678 38436 25712
rect 38470 25678 38536 25712
rect 38570 25678 38616 25712
rect 28624 25612 38616 25678
rect 28624 25578 28656 25612
rect 28690 25578 28756 25612
rect 28790 25578 28856 25612
rect 28890 25578 28956 25612
rect 28990 25578 29056 25612
rect 29090 25578 29156 25612
rect 29190 25578 29996 25612
rect 30030 25578 30096 25612
rect 30130 25578 30196 25612
rect 30230 25578 30296 25612
rect 30330 25578 30396 25612
rect 30430 25578 30496 25612
rect 30530 25578 31336 25612
rect 31370 25578 31436 25612
rect 31470 25578 31536 25612
rect 31570 25578 31636 25612
rect 31670 25578 31736 25612
rect 31770 25578 31836 25612
rect 31870 25578 32676 25612
rect 32710 25578 32776 25612
rect 32810 25578 32876 25612
rect 32910 25578 32976 25612
rect 33010 25578 33076 25612
rect 33110 25578 33176 25612
rect 33210 25578 34016 25612
rect 34050 25578 34116 25612
rect 34150 25578 34216 25612
rect 34250 25578 34316 25612
rect 34350 25578 34416 25612
rect 34450 25578 34516 25612
rect 34550 25578 35356 25612
rect 35390 25578 35456 25612
rect 35490 25578 35556 25612
rect 35590 25578 35656 25612
rect 35690 25578 35756 25612
rect 35790 25578 35856 25612
rect 35890 25578 36696 25612
rect 36730 25578 36796 25612
rect 36830 25578 36896 25612
rect 36930 25578 36996 25612
rect 37030 25578 37096 25612
rect 37130 25578 37196 25612
rect 37230 25578 38036 25612
rect 38070 25578 38136 25612
rect 38170 25578 38236 25612
rect 38270 25578 38336 25612
rect 38370 25578 38436 25612
rect 38470 25578 38536 25612
rect 38570 25578 38616 25612
rect 28624 25512 38616 25578
rect 28624 25478 28656 25512
rect 28690 25478 28756 25512
rect 28790 25478 28856 25512
rect 28890 25478 28956 25512
rect 28990 25478 29056 25512
rect 29090 25478 29156 25512
rect 29190 25478 29996 25512
rect 30030 25478 30096 25512
rect 30130 25478 30196 25512
rect 30230 25478 30296 25512
rect 30330 25478 30396 25512
rect 30430 25478 30496 25512
rect 30530 25478 31336 25512
rect 31370 25478 31436 25512
rect 31470 25478 31536 25512
rect 31570 25478 31636 25512
rect 31670 25478 31736 25512
rect 31770 25478 31836 25512
rect 31870 25478 32676 25512
rect 32710 25478 32776 25512
rect 32810 25478 32876 25512
rect 32910 25478 32976 25512
rect 33010 25478 33076 25512
rect 33110 25478 33176 25512
rect 33210 25478 34016 25512
rect 34050 25478 34116 25512
rect 34150 25478 34216 25512
rect 34250 25478 34316 25512
rect 34350 25478 34416 25512
rect 34450 25478 34516 25512
rect 34550 25478 35356 25512
rect 35390 25478 35456 25512
rect 35490 25478 35556 25512
rect 35590 25478 35656 25512
rect 35690 25478 35756 25512
rect 35790 25478 35856 25512
rect 35890 25478 36696 25512
rect 36730 25478 36796 25512
rect 36830 25478 36896 25512
rect 36930 25478 36996 25512
rect 37030 25478 37096 25512
rect 37130 25478 37196 25512
rect 37230 25478 38036 25512
rect 38070 25478 38136 25512
rect 38170 25478 38236 25512
rect 38270 25478 38336 25512
rect 38370 25478 38436 25512
rect 38470 25478 38536 25512
rect 38570 25478 38616 25512
rect 28624 25412 38616 25478
rect 28624 25378 28656 25412
rect 28690 25378 28756 25412
rect 28790 25378 28856 25412
rect 28890 25378 28956 25412
rect 28990 25378 29056 25412
rect 29090 25378 29156 25412
rect 29190 25378 29996 25412
rect 30030 25378 30096 25412
rect 30130 25378 30196 25412
rect 30230 25378 30296 25412
rect 30330 25378 30396 25412
rect 30430 25378 30496 25412
rect 30530 25378 31336 25412
rect 31370 25378 31436 25412
rect 31470 25378 31536 25412
rect 31570 25378 31636 25412
rect 31670 25378 31736 25412
rect 31770 25378 31836 25412
rect 31870 25378 32676 25412
rect 32710 25378 32776 25412
rect 32810 25378 32876 25412
rect 32910 25378 32976 25412
rect 33010 25378 33076 25412
rect 33110 25378 33176 25412
rect 33210 25378 34016 25412
rect 34050 25378 34116 25412
rect 34150 25378 34216 25412
rect 34250 25378 34316 25412
rect 34350 25378 34416 25412
rect 34450 25378 34516 25412
rect 34550 25378 35356 25412
rect 35390 25378 35456 25412
rect 35490 25378 35556 25412
rect 35590 25378 35656 25412
rect 35690 25378 35756 25412
rect 35790 25378 35856 25412
rect 35890 25378 36696 25412
rect 36730 25378 36796 25412
rect 36830 25378 36896 25412
rect 36930 25378 36996 25412
rect 37030 25378 37096 25412
rect 37130 25378 37196 25412
rect 37230 25378 38036 25412
rect 38070 25378 38136 25412
rect 38170 25378 38236 25412
rect 38270 25378 38336 25412
rect 38370 25378 38436 25412
rect 38470 25378 38536 25412
rect 38570 25378 38616 25412
rect 28624 25312 38616 25378
rect 28624 25278 28656 25312
rect 28690 25278 28756 25312
rect 28790 25278 28856 25312
rect 28890 25278 28956 25312
rect 28990 25278 29056 25312
rect 29090 25278 29156 25312
rect 29190 25278 29996 25312
rect 30030 25278 30096 25312
rect 30130 25278 30196 25312
rect 30230 25278 30296 25312
rect 30330 25278 30396 25312
rect 30430 25278 30496 25312
rect 30530 25278 31336 25312
rect 31370 25278 31436 25312
rect 31470 25278 31536 25312
rect 31570 25278 31636 25312
rect 31670 25278 31736 25312
rect 31770 25278 31836 25312
rect 31870 25278 32676 25312
rect 32710 25278 32776 25312
rect 32810 25278 32876 25312
rect 32910 25278 32976 25312
rect 33010 25278 33076 25312
rect 33110 25278 33176 25312
rect 33210 25278 34016 25312
rect 34050 25278 34116 25312
rect 34150 25278 34216 25312
rect 34250 25278 34316 25312
rect 34350 25278 34416 25312
rect 34450 25278 34516 25312
rect 34550 25278 35356 25312
rect 35390 25278 35456 25312
rect 35490 25278 35556 25312
rect 35590 25278 35656 25312
rect 35690 25278 35756 25312
rect 35790 25278 35856 25312
rect 35890 25278 36696 25312
rect 36730 25278 36796 25312
rect 36830 25278 36896 25312
rect 36930 25278 36996 25312
rect 37030 25278 37096 25312
rect 37130 25278 37196 25312
rect 37230 25278 38036 25312
rect 38070 25278 38136 25312
rect 38170 25278 38236 25312
rect 38270 25278 38336 25312
rect 38370 25278 38436 25312
rect 38470 25278 38536 25312
rect 38570 25278 38616 25312
rect 28624 25220 38616 25278
rect 28624 25168 28632 25220
rect 28684 25212 38616 25220
rect 28690 25178 28756 25212
rect 28790 25178 28856 25212
rect 28890 25178 28956 25212
rect 28990 25178 29056 25212
rect 29090 25178 29156 25212
rect 29190 25178 29996 25212
rect 30030 25178 30096 25212
rect 30130 25178 30196 25212
rect 30230 25178 30296 25212
rect 30330 25178 30396 25212
rect 30430 25178 30496 25212
rect 30530 25178 31336 25212
rect 31370 25178 31436 25212
rect 31470 25178 31536 25212
rect 31570 25178 31636 25212
rect 31670 25178 31736 25212
rect 31770 25178 31836 25212
rect 31870 25178 32676 25212
rect 32710 25178 32776 25212
rect 32810 25178 32876 25212
rect 32910 25178 32976 25212
rect 33010 25178 33076 25212
rect 33110 25178 33176 25212
rect 33210 25178 34016 25212
rect 34050 25178 34116 25212
rect 34150 25178 34216 25212
rect 34250 25178 34316 25212
rect 34350 25178 34416 25212
rect 34450 25178 34516 25212
rect 34550 25178 35356 25212
rect 35390 25178 35456 25212
rect 35490 25178 35556 25212
rect 35590 25178 35656 25212
rect 35690 25178 35756 25212
rect 35790 25178 35856 25212
rect 35890 25178 36696 25212
rect 36730 25178 36796 25212
rect 36830 25178 36896 25212
rect 36930 25178 36996 25212
rect 37030 25178 37096 25212
rect 37130 25178 37196 25212
rect 37230 25178 38036 25212
rect 38070 25178 38136 25212
rect 38170 25178 38236 25212
rect 38270 25178 38336 25212
rect 38370 25178 38436 25212
rect 38470 25178 38536 25212
rect 38570 25178 38616 25212
rect 28684 25168 38616 25178
rect 28624 25146 38616 25168
rect 27096 25112 27142 25135
rect 38672 25140 38700 25862
rect 39390 25644 39396 25696
rect 39448 25684 39454 25696
rect 39757 25684 39765 26141
rect 39448 25656 39765 25684
rect 39448 25644 39454 25656
rect 39757 25603 39765 25656
rect 40159 25603 40167 26141
rect 39757 25591 40167 25603
rect 41765 26141 42175 26153
rect 41765 25603 41772 26141
rect 42166 25603 42175 26141
rect 41765 25591 42175 25603
rect 39757 25181 40167 25193
rect 39757 25140 39765 25181
rect 38672 25112 39765 25140
rect 15079 25061 15125 25099
rect 15079 25027 15085 25061
rect 15119 25027 15125 25061
rect 15079 24989 15125 25027
rect 23382 25004 23388 25016
rect 15079 24955 15085 24989
rect 15119 24955 15125 24989
rect 23327 24976 23388 25004
rect 23382 24964 23388 24976
rect 23440 24964 23446 25016
rect 15079 24917 15125 24955
rect 39390 24936 39396 24948
rect 15079 24883 15085 24917
rect 15119 24883 15125 24917
rect 15079 24867 15125 24883
rect 27632 24908 39396 24936
rect 27632 24880 27660 24908
rect 39390 24896 39396 24908
rect 39448 24896 39454 24948
rect 23290 24868 23296 24880
rect 23235 24840 23296 24868
rect 23290 24828 23296 24840
rect 23348 24828 23354 24880
rect 27614 24828 27620 24880
rect 27672 24828 27678 24880
rect 9674 24664 9680 24676
rect 8728 24627 9160 24643
rect 9619 24636 9680 24664
rect 9674 24624 9680 24636
rect 9732 24624 9738 24676
rect 12526 24664 12532 24676
rect 12471 24636 12532 24664
rect 12526 24624 12532 24636
rect 12584 24624 12590 24676
rect 39757 24643 39765 25112
rect 40159 24643 40167 25181
rect 39757 24631 40167 24643
rect 41754 25181 42186 25591
rect 41754 24643 41772 25181
rect 42166 24643 42186 25181
rect 40052 24572 40080 24631
rect 41754 24627 42186 24643
rect 900 24570 47736 24572
rect 900 24454 922 24570
rect 2510 24540 46126 24570
rect 2510 24529 15476 24540
rect 2510 24495 6903 24529
rect 6937 24495 7103 24529
rect 7137 24495 7303 24529
rect 7337 24495 7503 24529
rect 7537 24495 7703 24529
rect 7737 24495 7903 24529
rect 7937 24495 8103 24529
rect 8137 24495 8303 24529
rect 8337 24495 8503 24529
rect 8537 24495 8703 24529
rect 8737 24495 8903 24529
rect 8937 24495 9725 24529
rect 9759 24495 10125 24529
rect 10159 24495 10525 24529
rect 10559 24495 10925 24529
rect 10959 24495 11325 24529
rect 11359 24495 11725 24529
rect 11759 24495 12125 24529
rect 12159 24495 12525 24529
rect 12559 24495 12925 24529
rect 12959 24495 13325 24529
rect 13359 24495 13725 24529
rect 13759 24495 14125 24529
rect 14159 24495 14525 24529
rect 14559 24495 14925 24529
rect 14959 24495 15476 24529
rect 2510 24488 15476 24495
rect 15528 24529 46126 24540
rect 15528 24495 15607 24529
rect 15641 24495 16007 24529
rect 16041 24495 16407 24529
rect 16441 24495 16807 24529
rect 16841 24495 17207 24529
rect 17241 24495 17607 24529
rect 17641 24495 18007 24529
rect 18041 24495 18407 24529
rect 18441 24495 18807 24529
rect 18841 24495 19207 24529
rect 19241 24495 19607 24529
rect 19641 24495 20007 24529
rect 20041 24495 20407 24529
rect 20441 24495 20807 24529
rect 20841 24495 21207 24529
rect 21241 24495 21607 24529
rect 21641 24495 22007 24529
rect 22041 24495 22407 24529
rect 22441 24495 23151 24529
rect 23185 24495 23551 24529
rect 23585 24495 23951 24529
rect 23985 24495 24351 24529
rect 24385 24495 24751 24529
rect 24785 24495 25151 24529
rect 25185 24495 25551 24529
rect 25585 24495 25951 24529
rect 25985 24495 26351 24529
rect 26385 24495 26751 24529
rect 26785 24495 28443 24529
rect 28477 24495 28643 24529
rect 28677 24495 28843 24529
rect 28877 24495 29043 24529
rect 29077 24495 29243 24529
rect 29277 24495 29443 24529
rect 29477 24495 29643 24529
rect 29677 24495 29843 24529
rect 29877 24495 30043 24529
rect 30077 24495 30243 24529
rect 30277 24495 30443 24529
rect 30477 24495 30643 24529
rect 30677 24495 30843 24529
rect 30877 24495 31043 24529
rect 31077 24495 31243 24529
rect 31277 24495 31443 24529
rect 31477 24495 31643 24529
rect 31677 24495 31843 24529
rect 31877 24495 32043 24529
rect 32077 24495 32243 24529
rect 32277 24495 32443 24529
rect 32477 24495 32643 24529
rect 32677 24495 32843 24529
rect 32877 24495 33043 24529
rect 33077 24495 33243 24529
rect 33277 24495 33443 24529
rect 33477 24495 33643 24529
rect 33677 24495 33843 24529
rect 33877 24495 34043 24529
rect 34077 24495 34243 24529
rect 34277 24495 34443 24529
rect 34477 24495 34643 24529
rect 34677 24495 34843 24529
rect 34877 24495 35043 24529
rect 35077 24495 35243 24529
rect 35277 24495 35443 24529
rect 35477 24495 35643 24529
rect 35677 24495 35843 24529
rect 35877 24495 36043 24529
rect 36077 24495 36243 24529
rect 36277 24495 36443 24529
rect 36477 24495 36643 24529
rect 36677 24495 36843 24529
rect 36877 24495 37043 24529
rect 37077 24495 37243 24529
rect 37277 24495 37443 24529
rect 37477 24495 37643 24529
rect 37677 24495 37843 24529
rect 37877 24495 38043 24529
rect 38077 24495 38243 24529
rect 38277 24495 38443 24529
rect 38477 24495 38643 24529
rect 38677 24495 38843 24529
rect 38877 24495 39929 24529
rect 39963 24495 40129 24529
rect 40163 24495 40329 24529
rect 40363 24495 40529 24529
rect 40563 24495 40729 24529
rect 40763 24495 40929 24529
rect 40963 24495 41129 24529
rect 41163 24495 41329 24529
rect 41363 24495 41529 24529
rect 41563 24495 41729 24529
rect 41763 24495 41929 24529
rect 41963 24495 46126 24529
rect 15528 24488 46126 24495
rect 2510 24454 46126 24488
rect 47714 24454 47736 24570
rect 900 24452 47736 24454
rect 7190 24216 7196 24268
rect 7248 24256 7254 24268
rect 13354 24256 13360 24268
rect 7248 24228 13360 24256
rect 7248 24216 7254 24228
rect 13354 24216 13360 24228
rect 13412 24216 13418 24268
rect 7098 23468 7104 23520
rect 7156 23508 7162 23520
rect 30098 23508 30104 23520
rect 7156 23480 30104 23508
rect 7156 23468 7162 23480
rect 30098 23468 30104 23480
rect 30156 23468 30162 23520
rect 3348 22690 45288 22692
rect 3348 22574 3370 22690
rect 4958 22649 43678 22690
rect 4958 22615 7863 22649
rect 7897 22615 8263 22649
rect 8297 22615 8663 22649
rect 8697 22615 9063 22649
rect 9097 22615 9463 22649
rect 9497 22615 9863 22649
rect 9897 22615 10263 22649
rect 10297 22615 10663 22649
rect 10697 22615 11063 22649
rect 11097 22615 11463 22649
rect 11497 22615 11863 22649
rect 11897 22615 12263 22649
rect 12297 22615 12663 22649
rect 12697 22615 13063 22649
rect 13097 22615 13745 22649
rect 13779 22615 14145 22649
rect 14179 22615 14545 22649
rect 14579 22615 14945 22649
rect 14979 22615 15345 22649
rect 15379 22615 15745 22649
rect 15779 22615 16145 22649
rect 16179 22615 16545 22649
rect 16579 22615 16945 22649
rect 16979 22615 17345 22649
rect 17379 22615 17745 22649
rect 17779 22615 18145 22649
rect 18179 22615 18545 22649
rect 18579 22615 18945 22649
rect 18979 22615 19345 22649
rect 19379 22615 19745 22649
rect 19779 22615 20145 22649
rect 20179 22615 20545 22649
rect 20579 22615 21191 22649
rect 21225 22615 21391 22649
rect 21425 22615 21591 22649
rect 21625 22615 21791 22649
rect 21825 22615 21991 22649
rect 22025 22615 22191 22649
rect 22225 22615 23151 22649
rect 23185 22615 23551 22649
rect 23585 22615 23951 22649
rect 23985 22615 24351 22649
rect 24385 22615 24751 22649
rect 24785 22615 25151 22649
rect 25185 22615 25551 22649
rect 25585 22615 25951 22649
rect 25985 22615 26351 22649
rect 26385 22615 26751 22649
rect 26785 22615 28443 22649
rect 28477 22615 28643 22649
rect 28677 22615 28843 22649
rect 28877 22615 29043 22649
rect 29077 22615 29243 22649
rect 29277 22615 29443 22649
rect 29477 22615 29643 22649
rect 29677 22615 29843 22649
rect 29877 22615 30043 22649
rect 30077 22615 30243 22649
rect 30277 22615 30443 22649
rect 30477 22615 30643 22649
rect 30677 22615 30843 22649
rect 30877 22615 31043 22649
rect 31077 22615 31243 22649
rect 31277 22615 31443 22649
rect 31477 22615 31643 22649
rect 31677 22615 31843 22649
rect 31877 22615 32043 22649
rect 32077 22615 32243 22649
rect 32277 22615 32443 22649
rect 32477 22615 32643 22649
rect 32677 22615 32843 22649
rect 32877 22615 33043 22649
rect 33077 22615 33243 22649
rect 33277 22615 33443 22649
rect 33477 22615 33643 22649
rect 33677 22615 33843 22649
rect 33877 22615 34043 22649
rect 34077 22615 34243 22649
rect 34277 22615 34443 22649
rect 34477 22615 34643 22649
rect 34677 22615 34843 22649
rect 34877 22615 35043 22649
rect 35077 22615 35243 22649
rect 35277 22615 35443 22649
rect 35477 22615 35643 22649
rect 35677 22615 35843 22649
rect 35877 22615 36043 22649
rect 36077 22615 36243 22649
rect 36277 22615 36443 22649
rect 36477 22615 36643 22649
rect 36677 22615 36843 22649
rect 36877 22615 37043 22649
rect 37077 22615 37243 22649
rect 37277 22615 37443 22649
rect 37477 22615 37643 22649
rect 37677 22615 37843 22649
rect 37877 22615 38043 22649
rect 38077 22615 38243 22649
rect 38277 22615 38443 22649
rect 38477 22615 38643 22649
rect 38677 22615 38843 22649
rect 38877 22615 39929 22649
rect 39963 22615 40129 22649
rect 40163 22615 40329 22649
rect 40363 22615 40529 22649
rect 40563 22615 40729 22649
rect 40763 22615 40929 22649
rect 40963 22615 41129 22649
rect 41163 22615 41329 22649
rect 41363 22615 41529 22649
rect 41563 22615 41729 22649
rect 41763 22615 41929 22649
rect 41963 22615 43678 22649
rect 4958 22574 43678 22615
rect 45266 22574 45288 22690
rect 3348 22572 45288 22574
rect 8312 22500 8340 22572
rect 8294 22448 8300 22500
rect 8352 22448 8358 22500
rect 26418 22488 26424 22500
rect 26363 22460 26424 22488
rect 26418 22448 26424 22460
rect 26476 22448 26482 22500
rect 7721 22381 7767 22397
rect 7721 22347 7727 22381
rect 7761 22347 7767 22381
rect 7721 22309 7767 22347
rect 7721 22275 7727 22309
rect 7761 22275 7767 22309
rect 7721 22237 7767 22275
rect 7721 22203 7727 22237
rect 7761 22203 7767 22237
rect 7721 22165 7767 22203
rect 7721 22131 7727 22165
rect 7761 22131 7767 22165
rect 7721 22093 7767 22131
rect 7721 22059 7727 22093
rect 7761 22059 7767 22093
rect 7721 22021 7767 22059
rect 7721 21987 7727 22021
rect 7761 21987 7767 22021
rect 7721 21949 7767 21987
rect 7721 21915 7727 21949
rect 7761 21915 7767 21949
rect 7721 21877 7767 21915
rect 7721 21843 7727 21877
rect 7761 21843 7767 21877
rect 7721 21805 7767 21843
rect 7721 21771 7727 21805
rect 7761 21771 7767 21805
rect 7721 21733 7767 21771
rect 7721 21699 7727 21733
rect 7761 21699 7767 21733
rect 7721 21661 7767 21699
rect 7721 21627 7727 21661
rect 7761 21627 7767 21661
rect 7721 21589 7767 21627
rect 7721 21555 7727 21589
rect 7761 21555 7767 21589
rect 7721 21517 7767 21555
rect 7721 21483 7727 21517
rect 7761 21483 7767 21517
rect 7721 21445 7767 21483
rect 7721 21411 7727 21445
rect 7761 21411 7767 21445
rect 7721 21373 7767 21411
rect 7721 21339 7727 21373
rect 7761 21339 7767 21373
rect 7721 21301 7767 21339
rect 7721 21267 7727 21301
rect 7761 21267 7767 21301
rect 7721 21229 7767 21267
rect 7721 21195 7727 21229
rect 7761 21195 7767 21229
rect 7721 21157 7767 21195
rect 7721 21123 7727 21157
rect 7761 21123 7767 21157
rect 7721 21107 7767 21123
rect 8179 22381 8225 22397
rect 8179 22347 8185 22381
rect 8219 22347 8225 22381
rect 8179 22309 8225 22347
rect 8179 22275 8185 22309
rect 8219 22275 8225 22309
rect 8179 22237 8225 22275
rect 8179 22203 8185 22237
rect 8219 22203 8225 22237
rect 8179 22165 8225 22203
rect 8179 22131 8185 22165
rect 8219 22131 8225 22165
rect 8179 22093 8225 22131
rect 8179 22059 8185 22093
rect 8219 22059 8225 22093
rect 8179 22021 8225 22059
rect 8179 21987 8185 22021
rect 8219 21987 8225 22021
rect 8179 21949 8225 21987
rect 8179 21915 8185 21949
rect 8219 21915 8225 21949
rect 8179 21877 8225 21915
rect 8179 21843 8185 21877
rect 8219 21843 8225 21877
rect 8179 21805 8225 21843
rect 8179 21771 8185 21805
rect 8219 21771 8225 21805
rect 8179 21733 8225 21771
rect 8179 21699 8185 21733
rect 8219 21699 8225 21733
rect 8179 21661 8225 21699
rect 8179 21627 8185 21661
rect 8219 21627 8225 21661
rect 8179 21589 8225 21627
rect 8179 21555 8185 21589
rect 8219 21555 8225 21589
rect 8179 21517 8225 21555
rect 8179 21483 8185 21517
rect 8219 21483 8225 21517
rect 8179 21445 8225 21483
rect 8179 21411 8185 21445
rect 8219 21411 8225 21445
rect 8179 21373 8225 21411
rect 8179 21339 8185 21373
rect 8219 21339 8225 21373
rect 8179 21301 8225 21339
rect 8179 21267 8185 21301
rect 8219 21267 8225 21301
rect 8179 21229 8225 21267
rect 8179 21195 8185 21229
rect 8219 21195 8225 21229
rect 8179 21157 8225 21195
rect 8179 21123 8185 21157
rect 8219 21123 8225 21157
rect 8179 21107 8225 21123
rect 8637 22381 8683 22397
rect 8637 22347 8643 22381
rect 8677 22347 8683 22381
rect 8637 22309 8683 22347
rect 8637 22275 8643 22309
rect 8677 22275 8683 22309
rect 8637 22237 8683 22275
rect 8637 22203 8643 22237
rect 8677 22203 8683 22237
rect 8637 22165 8683 22203
rect 8637 22131 8643 22165
rect 8677 22131 8683 22165
rect 8637 22093 8683 22131
rect 8637 22059 8643 22093
rect 8677 22059 8683 22093
rect 8637 22021 8683 22059
rect 8637 21987 8643 22021
rect 8677 21987 8683 22021
rect 8637 21949 8683 21987
rect 8637 21915 8643 21949
rect 8677 21915 8683 21949
rect 8637 21877 8683 21915
rect 8637 21843 8643 21877
rect 8677 21843 8683 21877
rect 8637 21805 8683 21843
rect 8637 21771 8643 21805
rect 8677 21771 8683 21805
rect 8637 21733 8683 21771
rect 8637 21699 8643 21733
rect 8677 21699 8683 21733
rect 8637 21661 8683 21699
rect 8637 21627 8643 21661
rect 8677 21627 8683 21661
rect 8637 21589 8683 21627
rect 8637 21555 8643 21589
rect 8677 21555 8683 21589
rect 8637 21517 8683 21555
rect 8637 21483 8643 21517
rect 8677 21483 8683 21517
rect 8637 21445 8683 21483
rect 8637 21411 8643 21445
rect 8677 21411 8683 21445
rect 8637 21373 8683 21411
rect 8637 21339 8643 21373
rect 8677 21339 8683 21373
rect 8637 21301 8683 21339
rect 8637 21267 8643 21301
rect 8677 21267 8683 21301
rect 8637 21229 8683 21267
rect 8637 21195 8643 21229
rect 8677 21195 8683 21229
rect 8637 21157 8683 21195
rect 8637 21123 8643 21157
rect 8677 21123 8683 21157
rect 8637 21107 8683 21123
rect 9095 22381 9141 22397
rect 9095 22347 9101 22381
rect 9135 22347 9141 22381
rect 9095 22309 9141 22347
rect 9095 22275 9101 22309
rect 9135 22275 9141 22309
rect 9095 22237 9141 22275
rect 9095 22203 9101 22237
rect 9135 22203 9141 22237
rect 9095 22165 9141 22203
rect 9095 22131 9101 22165
rect 9135 22131 9141 22165
rect 9095 22093 9141 22131
rect 9095 22059 9101 22093
rect 9135 22059 9141 22093
rect 9095 22021 9141 22059
rect 9095 21987 9101 22021
rect 9135 21987 9141 22021
rect 9095 21949 9141 21987
rect 9095 21915 9101 21949
rect 9135 21915 9141 21949
rect 9095 21877 9141 21915
rect 9095 21843 9101 21877
rect 9135 21843 9141 21877
rect 9095 21805 9141 21843
rect 9095 21771 9101 21805
rect 9135 21771 9141 21805
rect 9095 21733 9141 21771
rect 9095 21699 9101 21733
rect 9135 21699 9141 21733
rect 9095 21661 9141 21699
rect 9095 21627 9101 21661
rect 9135 21627 9141 21661
rect 9095 21589 9141 21627
rect 9095 21555 9101 21589
rect 9135 21555 9141 21589
rect 9095 21517 9141 21555
rect 9095 21483 9101 21517
rect 9135 21483 9141 21517
rect 9095 21445 9141 21483
rect 9095 21411 9101 21445
rect 9135 21411 9141 21445
rect 9095 21373 9141 21411
rect 9095 21339 9101 21373
rect 9135 21339 9141 21373
rect 9095 21301 9141 21339
rect 9095 21267 9101 21301
rect 9135 21267 9141 21301
rect 9095 21229 9141 21267
rect 9095 21195 9101 21229
rect 9135 21195 9141 21229
rect 9095 21157 9141 21195
rect 9095 21123 9101 21157
rect 9135 21123 9141 21157
rect 9095 21107 9141 21123
rect 9553 22381 9599 22397
rect 9553 22347 9559 22381
rect 9593 22347 9599 22381
rect 9553 22309 9599 22347
rect 9553 22275 9559 22309
rect 9593 22275 9599 22309
rect 9553 22237 9599 22275
rect 9553 22203 9559 22237
rect 9593 22203 9599 22237
rect 9553 22165 9599 22203
rect 9553 22131 9559 22165
rect 9593 22131 9599 22165
rect 9553 22093 9599 22131
rect 9553 22059 9559 22093
rect 9593 22059 9599 22093
rect 9553 22021 9599 22059
rect 9553 21987 9559 22021
rect 9593 21987 9599 22021
rect 9553 21949 9599 21987
rect 9553 21915 9559 21949
rect 9593 21915 9599 21949
rect 9553 21877 9599 21915
rect 9553 21843 9559 21877
rect 9593 21843 9599 21877
rect 9553 21805 9599 21843
rect 9553 21771 9559 21805
rect 9593 21771 9599 21805
rect 9553 21733 9599 21771
rect 9553 21699 9559 21733
rect 9593 21699 9599 21733
rect 9553 21661 9599 21699
rect 9553 21627 9559 21661
rect 9593 21627 9599 21661
rect 9553 21589 9599 21627
rect 9553 21555 9559 21589
rect 9593 21555 9599 21589
rect 9553 21517 9599 21555
rect 9553 21483 9559 21517
rect 9593 21483 9599 21517
rect 9553 21445 9599 21483
rect 9553 21411 9559 21445
rect 9593 21411 9599 21445
rect 9553 21373 9599 21411
rect 9553 21339 9559 21373
rect 9593 21339 9599 21373
rect 9553 21301 9599 21339
rect 9553 21267 9559 21301
rect 9593 21267 9599 21301
rect 9553 21229 9599 21267
rect 9553 21195 9559 21229
rect 9593 21195 9599 21229
rect 9553 21157 9599 21195
rect 9553 21123 9559 21157
rect 9593 21123 9599 21157
rect 9553 21107 9599 21123
rect 10011 22381 10057 22397
rect 10011 22347 10017 22381
rect 10051 22347 10057 22381
rect 10011 22309 10057 22347
rect 10011 22275 10017 22309
rect 10051 22275 10057 22309
rect 10011 22237 10057 22275
rect 10011 22203 10017 22237
rect 10051 22203 10057 22237
rect 10011 22165 10057 22203
rect 10011 22131 10017 22165
rect 10051 22131 10057 22165
rect 10011 22093 10057 22131
rect 10011 22059 10017 22093
rect 10051 22059 10057 22093
rect 10011 22021 10057 22059
rect 10011 21987 10017 22021
rect 10051 21987 10057 22021
rect 10011 21949 10057 21987
rect 10011 21915 10017 21949
rect 10051 21915 10057 21949
rect 10011 21877 10057 21915
rect 10011 21843 10017 21877
rect 10051 21843 10057 21877
rect 10011 21805 10057 21843
rect 10011 21771 10017 21805
rect 10051 21771 10057 21805
rect 10011 21733 10057 21771
rect 10011 21699 10017 21733
rect 10051 21699 10057 21733
rect 10011 21661 10057 21699
rect 10011 21627 10017 21661
rect 10051 21627 10057 21661
rect 10011 21589 10057 21627
rect 10011 21555 10017 21589
rect 10051 21555 10057 21589
rect 10011 21517 10057 21555
rect 10011 21483 10017 21517
rect 10051 21483 10057 21517
rect 10011 21445 10057 21483
rect 10011 21411 10017 21445
rect 10051 21411 10057 21445
rect 10011 21373 10057 21411
rect 10011 21339 10017 21373
rect 10051 21339 10057 21373
rect 10011 21301 10057 21339
rect 10011 21267 10017 21301
rect 10051 21267 10057 21301
rect 10011 21229 10057 21267
rect 10011 21195 10017 21229
rect 10051 21195 10057 21229
rect 10011 21157 10057 21195
rect 10011 21123 10017 21157
rect 10051 21123 10057 21157
rect 10011 21107 10057 21123
rect 10469 22381 10515 22397
rect 10469 22347 10475 22381
rect 10509 22347 10515 22381
rect 10469 22309 10515 22347
rect 10469 22275 10475 22309
rect 10509 22275 10515 22309
rect 10469 22237 10515 22275
rect 10469 22203 10475 22237
rect 10509 22203 10515 22237
rect 10469 22165 10515 22203
rect 10469 22131 10475 22165
rect 10509 22131 10515 22165
rect 10469 22093 10515 22131
rect 10469 22059 10475 22093
rect 10509 22059 10515 22093
rect 10469 22021 10515 22059
rect 10469 21987 10475 22021
rect 10509 21987 10515 22021
rect 10469 21949 10515 21987
rect 10469 21915 10475 21949
rect 10509 21915 10515 21949
rect 10469 21877 10515 21915
rect 10469 21843 10475 21877
rect 10509 21843 10515 21877
rect 10469 21805 10515 21843
rect 10469 21771 10475 21805
rect 10509 21771 10515 21805
rect 10469 21733 10515 21771
rect 10469 21699 10475 21733
rect 10509 21699 10515 21733
rect 10469 21661 10515 21699
rect 10469 21627 10475 21661
rect 10509 21627 10515 21661
rect 10469 21589 10515 21627
rect 10469 21555 10475 21589
rect 10509 21555 10515 21589
rect 10469 21517 10515 21555
rect 10469 21483 10475 21517
rect 10509 21483 10515 21517
rect 10469 21445 10515 21483
rect 10469 21411 10475 21445
rect 10509 21411 10515 21445
rect 10469 21373 10515 21411
rect 10469 21339 10475 21373
rect 10509 21339 10515 21373
rect 10469 21301 10515 21339
rect 10469 21267 10475 21301
rect 10509 21267 10515 21301
rect 10469 21229 10515 21267
rect 10469 21195 10475 21229
rect 10509 21195 10515 21229
rect 10469 21157 10515 21195
rect 10469 21123 10475 21157
rect 10509 21123 10515 21157
rect 10469 21107 10515 21123
rect 10927 22381 10973 22397
rect 10927 22347 10933 22381
rect 10967 22347 10973 22381
rect 10927 22309 10973 22347
rect 10927 22275 10933 22309
rect 10967 22275 10973 22309
rect 10927 22237 10973 22275
rect 10927 22203 10933 22237
rect 10967 22203 10973 22237
rect 10927 22165 10973 22203
rect 10927 22131 10933 22165
rect 10967 22131 10973 22165
rect 10927 22093 10973 22131
rect 10927 22059 10933 22093
rect 10967 22059 10973 22093
rect 10927 22021 10973 22059
rect 10927 21987 10933 22021
rect 10967 21987 10973 22021
rect 10927 21949 10973 21987
rect 10927 21915 10933 21949
rect 10967 21915 10973 21949
rect 10927 21877 10973 21915
rect 10927 21843 10933 21877
rect 10967 21843 10973 21877
rect 10927 21805 10973 21843
rect 10927 21771 10933 21805
rect 10967 21771 10973 21805
rect 10927 21733 10973 21771
rect 10927 21699 10933 21733
rect 10967 21699 10973 21733
rect 10927 21661 10973 21699
rect 10927 21627 10933 21661
rect 10967 21627 10973 21661
rect 10927 21589 10973 21627
rect 10927 21555 10933 21589
rect 10967 21555 10973 21589
rect 10927 21517 10973 21555
rect 10927 21483 10933 21517
rect 10967 21483 10973 21517
rect 10927 21445 10973 21483
rect 10927 21411 10933 21445
rect 10967 21411 10973 21445
rect 10927 21373 10973 21411
rect 10927 21339 10933 21373
rect 10967 21339 10973 21373
rect 10927 21301 10973 21339
rect 10927 21267 10933 21301
rect 10967 21267 10973 21301
rect 10927 21229 10973 21267
rect 10927 21195 10933 21229
rect 10967 21195 10973 21229
rect 10927 21157 10973 21195
rect 10927 21123 10933 21157
rect 10967 21123 10973 21157
rect 10927 21107 10973 21123
rect 11385 22381 11431 22397
rect 11385 22347 11391 22381
rect 11425 22347 11431 22381
rect 11385 22309 11431 22347
rect 11385 22275 11391 22309
rect 11425 22275 11431 22309
rect 11385 22237 11431 22275
rect 11385 22203 11391 22237
rect 11425 22203 11431 22237
rect 11385 22165 11431 22203
rect 11385 22131 11391 22165
rect 11425 22131 11431 22165
rect 11385 22093 11431 22131
rect 11385 22059 11391 22093
rect 11425 22059 11431 22093
rect 11385 22021 11431 22059
rect 11385 21987 11391 22021
rect 11425 21987 11431 22021
rect 11385 21949 11431 21987
rect 11385 21915 11391 21949
rect 11425 21915 11431 21949
rect 11385 21877 11431 21915
rect 11385 21843 11391 21877
rect 11425 21843 11431 21877
rect 11385 21805 11431 21843
rect 11385 21771 11391 21805
rect 11425 21771 11431 21805
rect 11385 21733 11431 21771
rect 11385 21699 11391 21733
rect 11425 21699 11431 21733
rect 11385 21661 11431 21699
rect 11385 21627 11391 21661
rect 11425 21627 11431 21661
rect 11385 21589 11431 21627
rect 11385 21555 11391 21589
rect 11425 21555 11431 21589
rect 11385 21517 11431 21555
rect 11385 21483 11391 21517
rect 11425 21483 11431 21517
rect 11385 21445 11431 21483
rect 11385 21411 11391 21445
rect 11425 21411 11431 21445
rect 11385 21373 11431 21411
rect 11385 21339 11391 21373
rect 11425 21339 11431 21373
rect 11385 21301 11431 21339
rect 11385 21267 11391 21301
rect 11425 21267 11431 21301
rect 11385 21229 11431 21267
rect 11385 21195 11391 21229
rect 11425 21195 11431 21229
rect 11385 21157 11431 21195
rect 11385 21123 11391 21157
rect 11425 21123 11431 21157
rect 11385 21107 11431 21123
rect 11843 22381 11889 22397
rect 11843 22347 11849 22381
rect 11883 22347 11889 22381
rect 11843 22309 11889 22347
rect 11843 22275 11849 22309
rect 11883 22275 11889 22309
rect 11843 22237 11889 22275
rect 11843 22203 11849 22237
rect 11883 22203 11889 22237
rect 11843 22165 11889 22203
rect 11843 22131 11849 22165
rect 11883 22131 11889 22165
rect 11843 22093 11889 22131
rect 11843 22059 11849 22093
rect 11883 22059 11889 22093
rect 11843 22021 11889 22059
rect 11843 21987 11849 22021
rect 11883 21987 11889 22021
rect 11843 21949 11889 21987
rect 11843 21915 11849 21949
rect 11883 21915 11889 21949
rect 11843 21877 11889 21915
rect 11843 21843 11849 21877
rect 11883 21843 11889 21877
rect 11843 21805 11889 21843
rect 11843 21771 11849 21805
rect 11883 21771 11889 21805
rect 11843 21733 11889 21771
rect 11843 21699 11849 21733
rect 11883 21699 11889 21733
rect 11843 21661 11889 21699
rect 11843 21627 11849 21661
rect 11883 21627 11889 21661
rect 11843 21589 11889 21627
rect 11843 21555 11849 21589
rect 11883 21555 11889 21589
rect 11843 21517 11889 21555
rect 11843 21483 11849 21517
rect 11883 21483 11889 21517
rect 11843 21445 11889 21483
rect 11843 21411 11849 21445
rect 11883 21411 11889 21445
rect 11843 21373 11889 21411
rect 11843 21339 11849 21373
rect 11883 21339 11889 21373
rect 11843 21301 11889 21339
rect 11843 21267 11849 21301
rect 11883 21267 11889 21301
rect 11843 21229 11889 21267
rect 11843 21195 11849 21229
rect 11883 21195 11889 21229
rect 11843 21157 11889 21195
rect 11843 21123 11849 21157
rect 11883 21123 11889 21157
rect 11843 21107 11889 21123
rect 12301 22381 12347 22397
rect 12301 22347 12307 22381
rect 12341 22347 12347 22381
rect 12301 22309 12347 22347
rect 12301 22275 12307 22309
rect 12341 22275 12347 22309
rect 12301 22237 12347 22275
rect 12301 22203 12307 22237
rect 12341 22203 12347 22237
rect 12301 22165 12347 22203
rect 12301 22131 12307 22165
rect 12341 22131 12347 22165
rect 12301 22093 12347 22131
rect 12301 22059 12307 22093
rect 12341 22059 12347 22093
rect 12301 22021 12347 22059
rect 12301 21987 12307 22021
rect 12341 21987 12347 22021
rect 12301 21949 12347 21987
rect 12301 21915 12307 21949
rect 12341 21915 12347 21949
rect 12301 21877 12347 21915
rect 12301 21843 12307 21877
rect 12341 21843 12347 21877
rect 12301 21805 12347 21843
rect 12301 21771 12307 21805
rect 12341 21771 12347 21805
rect 12301 21733 12347 21771
rect 12301 21699 12307 21733
rect 12341 21699 12347 21733
rect 12301 21661 12347 21699
rect 12301 21627 12307 21661
rect 12341 21627 12347 21661
rect 12301 21589 12347 21627
rect 12301 21555 12307 21589
rect 12341 21555 12347 21589
rect 12301 21517 12347 21555
rect 12301 21483 12307 21517
rect 12341 21483 12347 21517
rect 12301 21445 12347 21483
rect 12301 21411 12307 21445
rect 12341 21411 12347 21445
rect 12301 21373 12347 21411
rect 12301 21339 12307 21373
rect 12341 21339 12347 21373
rect 12301 21301 12347 21339
rect 12301 21267 12307 21301
rect 12341 21267 12347 21301
rect 12301 21229 12347 21267
rect 12301 21195 12307 21229
rect 12341 21195 12347 21229
rect 12301 21157 12347 21195
rect 12301 21123 12307 21157
rect 12341 21123 12347 21157
rect 12301 21107 12347 21123
rect 12759 22381 12805 22397
rect 12759 22347 12765 22381
rect 12799 22347 12805 22381
rect 12759 22309 12805 22347
rect 12759 22275 12765 22309
rect 12799 22275 12805 22309
rect 12759 22237 12805 22275
rect 12759 22203 12765 22237
rect 12799 22203 12805 22237
rect 12759 22165 12805 22203
rect 12759 22131 12765 22165
rect 12799 22131 12805 22165
rect 12759 22093 12805 22131
rect 12759 22059 12765 22093
rect 12799 22059 12805 22093
rect 12759 22021 12805 22059
rect 12759 21987 12765 22021
rect 12799 21987 12805 22021
rect 12759 21949 12805 21987
rect 12759 21915 12765 21949
rect 12799 21915 12805 21949
rect 12759 21877 12805 21915
rect 12759 21843 12765 21877
rect 12799 21843 12805 21877
rect 12759 21805 12805 21843
rect 12759 21771 12765 21805
rect 12799 21771 12805 21805
rect 12759 21733 12805 21771
rect 12759 21699 12765 21733
rect 12799 21699 12805 21733
rect 12759 21661 12805 21699
rect 12759 21627 12765 21661
rect 12799 21627 12805 21661
rect 12759 21589 12805 21627
rect 12759 21555 12765 21589
rect 12799 21555 12805 21589
rect 12759 21517 12805 21555
rect 12759 21483 12765 21517
rect 12799 21483 12805 21517
rect 12759 21445 12805 21483
rect 12759 21411 12765 21445
rect 12799 21411 12805 21445
rect 12759 21373 12805 21411
rect 12759 21339 12765 21373
rect 12799 21339 12805 21373
rect 12759 21301 12805 21339
rect 12759 21267 12765 21301
rect 12799 21267 12805 21301
rect 12759 21229 12805 21267
rect 12759 21195 12765 21229
rect 12799 21195 12805 21229
rect 12759 21157 12805 21195
rect 12759 21123 12765 21157
rect 12799 21123 12805 21157
rect 12759 21107 12805 21123
rect 13217 22381 13263 22397
rect 13217 22347 13223 22381
rect 13257 22347 13263 22381
rect 38654 22380 38660 22432
rect 38712 22420 38718 22432
rect 38712 22392 39068 22420
rect 38712 22380 38718 22392
rect 13217 22309 13263 22347
rect 39040 22352 39068 22392
rect 39757 22381 40167 22393
rect 39757 22352 39765 22381
rect 39040 22324 39765 22352
rect 13217 22275 13223 22309
rect 13257 22275 13263 22309
rect 13217 22237 13263 22275
rect 28286 22316 38954 22322
rect 28286 22282 28306 22316
rect 28340 22282 28396 22316
rect 28430 22282 28486 22316
rect 28520 22282 28576 22316
rect 28610 22282 28666 22316
rect 28700 22282 28756 22316
rect 28790 22282 28846 22316
rect 28880 22282 28936 22316
rect 28970 22282 29026 22316
rect 29060 22282 29116 22316
rect 29150 22282 29206 22316
rect 29240 22282 29296 22316
rect 29330 22282 29386 22316
rect 29420 22282 29476 22316
rect 29510 22282 29646 22316
rect 29680 22282 29736 22316
rect 29770 22282 29826 22316
rect 29860 22282 29916 22316
rect 29950 22282 30006 22316
rect 30040 22282 30096 22316
rect 30130 22282 30186 22316
rect 30220 22282 30276 22316
rect 30310 22282 30366 22316
rect 30400 22282 30456 22316
rect 30490 22282 30546 22316
rect 30580 22282 30636 22316
rect 30670 22282 30726 22316
rect 30760 22282 30816 22316
rect 30850 22282 30986 22316
rect 31020 22282 31076 22316
rect 31110 22282 31166 22316
rect 31200 22282 31256 22316
rect 31290 22282 31346 22316
rect 31380 22282 31436 22316
rect 31470 22282 31526 22316
rect 31560 22282 31616 22316
rect 31650 22282 31706 22316
rect 31740 22282 31796 22316
rect 31830 22282 31886 22316
rect 31920 22282 31976 22316
rect 32010 22282 32066 22316
rect 32100 22282 32156 22316
rect 32190 22282 32326 22316
rect 32360 22282 32416 22316
rect 32450 22282 32506 22316
rect 32540 22282 32596 22316
rect 32630 22282 32686 22316
rect 32720 22282 32776 22316
rect 32810 22282 32866 22316
rect 32900 22282 32956 22316
rect 32990 22282 33046 22316
rect 33080 22282 33136 22316
rect 33170 22282 33226 22316
rect 33260 22282 33316 22316
rect 33350 22282 33406 22316
rect 33440 22282 33496 22316
rect 33530 22282 33666 22316
rect 33700 22282 33756 22316
rect 33790 22282 33846 22316
rect 33880 22282 33936 22316
rect 33970 22282 34026 22316
rect 34060 22282 34116 22316
rect 34150 22282 34206 22316
rect 34240 22282 34296 22316
rect 34330 22282 34386 22316
rect 34420 22282 34476 22316
rect 34510 22282 34566 22316
rect 34600 22282 34656 22316
rect 34690 22282 34746 22316
rect 34780 22282 34836 22316
rect 34870 22282 35006 22316
rect 35040 22282 35096 22316
rect 35130 22282 35186 22316
rect 35220 22282 35276 22316
rect 35310 22282 35366 22316
rect 35400 22282 35456 22316
rect 35490 22282 35546 22316
rect 35580 22282 35636 22316
rect 35670 22282 35726 22316
rect 35760 22282 35816 22316
rect 35850 22282 35906 22316
rect 35940 22282 35996 22316
rect 36030 22282 36086 22316
rect 36120 22282 36176 22316
rect 36210 22282 36346 22316
rect 36380 22282 36436 22316
rect 36470 22282 36526 22316
rect 36560 22282 36616 22316
rect 36650 22282 36706 22316
rect 36740 22282 36796 22316
rect 36830 22282 36886 22316
rect 36920 22282 36976 22316
rect 37010 22282 37066 22316
rect 37100 22282 37156 22316
rect 37190 22282 37246 22316
rect 37280 22282 37336 22316
rect 37370 22282 37426 22316
rect 37460 22282 37516 22316
rect 37550 22282 37686 22316
rect 37720 22282 37776 22316
rect 37810 22282 37866 22316
rect 37900 22282 37956 22316
rect 37990 22282 38046 22316
rect 38080 22282 38136 22316
rect 38170 22282 38226 22316
rect 38260 22282 38316 22316
rect 38350 22282 38406 22316
rect 38440 22282 38496 22316
rect 38530 22282 38586 22316
rect 38620 22282 38676 22316
rect 38710 22282 38766 22316
rect 38800 22282 38856 22316
rect 38890 22282 38954 22316
rect 28286 22252 38954 22282
rect 13217 22203 13223 22237
rect 13257 22203 13263 22237
rect 23290 22216 23296 22228
rect 13217 22165 13263 22203
rect 13217 22131 13223 22165
rect 13257 22131 13263 22165
rect 13217 22093 13263 22131
rect 13217 22059 13223 22093
rect 13257 22059 13263 22093
rect 13217 22021 13263 22059
rect 13217 21987 13223 22021
rect 13257 21987 13263 22021
rect 22848 22188 23296 22216
rect 13217 21949 13263 21987
rect 13217 21915 13223 21949
rect 13257 21915 13263 21949
rect 13217 21877 13263 21915
rect 13217 21843 13223 21877
rect 13257 21843 13263 21877
rect 13217 21805 13263 21843
rect 13217 21771 13223 21805
rect 13257 21771 13263 21805
rect 13217 21733 13263 21771
rect 13217 21699 13223 21733
rect 13257 21699 13263 21733
rect 13217 21661 13263 21699
rect 13217 21627 13223 21661
rect 13257 21627 13263 21661
rect 13217 21589 13263 21627
rect 21373 21952 21983 21997
rect 21373 21918 21404 21952
rect 21438 21918 21504 21952
rect 21538 21918 21604 21952
rect 21638 21918 21704 21952
rect 21738 21918 21804 21952
rect 21838 21918 21904 21952
rect 21938 21944 21983 21952
rect 22848 21944 22876 22188
rect 23290 22176 23296 22188
rect 23348 22176 23354 22228
rect 30576 22172 30604 22252
rect 28450 22160 38790 22172
rect 28450 22156 30564 22160
rect 21938 21918 22876 21944
rect 21373 21916 22876 21918
rect 22974 22129 23020 22152
rect 22974 22095 22980 22129
rect 23014 22095 23020 22129
rect 22974 22057 23020 22095
rect 22974 22023 22980 22057
rect 23014 22023 23020 22057
rect 22974 21985 23020 22023
rect 22974 21951 22980 21985
rect 23014 21951 23020 21985
rect 21373 21852 21983 21916
rect 21373 21818 21404 21852
rect 21438 21818 21504 21852
rect 21538 21818 21604 21852
rect 21638 21818 21704 21852
rect 21738 21818 21804 21852
rect 21838 21818 21904 21852
rect 21938 21818 21983 21852
rect 21373 21752 21983 21818
rect 21373 21718 21404 21752
rect 21438 21718 21504 21752
rect 21538 21718 21604 21752
rect 21638 21718 21704 21752
rect 21738 21718 21804 21752
rect 21838 21718 21904 21752
rect 21938 21718 21983 21752
rect 21373 21652 21983 21718
rect 21373 21618 21404 21652
rect 21438 21618 21504 21652
rect 21538 21618 21604 21652
rect 21638 21618 21704 21652
rect 21738 21618 21804 21652
rect 21838 21618 21904 21652
rect 21938 21618 21983 21652
rect 13217 21555 13223 21589
rect 13257 21555 13263 21589
rect 20898 21564 20904 21616
rect 20956 21604 20962 21616
rect 21373 21604 21983 21618
rect 20956 21576 21983 21604
rect 20956 21564 20962 21576
rect 13217 21517 13263 21555
rect 13217 21483 13223 21517
rect 13257 21483 13263 21517
rect 13217 21445 13263 21483
rect 13217 21411 13223 21445
rect 13257 21411 13263 21445
rect 13217 21373 13263 21411
rect 21373 21552 21983 21576
rect 21373 21518 21404 21552
rect 21438 21518 21504 21552
rect 21538 21518 21604 21552
rect 21638 21518 21704 21552
rect 21738 21518 21804 21552
rect 21838 21518 21904 21552
rect 21938 21518 21983 21552
rect 21373 21452 21983 21518
rect 21373 21418 21404 21452
rect 21438 21418 21504 21452
rect 21538 21418 21604 21452
rect 21638 21418 21704 21452
rect 21738 21418 21804 21452
rect 21838 21418 21904 21452
rect 21938 21418 21983 21452
rect 21373 21387 21983 21418
rect 22974 21913 23020 21951
rect 22974 21879 22980 21913
rect 23014 21879 23020 21913
rect 22974 21841 23020 21879
rect 22974 21807 22980 21841
rect 23014 21807 23020 21841
rect 22974 21769 23020 21807
rect 22974 21735 22980 21769
rect 23014 21735 23020 21769
rect 22974 21697 23020 21735
rect 22974 21663 22980 21697
rect 23014 21663 23020 21697
rect 22974 21625 23020 21663
rect 22974 21591 22980 21625
rect 23014 21591 23020 21625
rect 22974 21553 23020 21591
rect 22974 21519 22980 21553
rect 23014 21519 23020 21553
rect 22974 21481 23020 21519
rect 22974 21447 22980 21481
rect 23014 21447 23020 21481
rect 22974 21409 23020 21447
rect 13217 21339 13223 21373
rect 13257 21339 13263 21373
rect 22974 21375 22980 21409
rect 23014 21375 23020 21409
rect 22974 21352 23020 21375
rect 23432 22129 23478 22152
rect 23432 22095 23438 22129
rect 23472 22095 23478 22129
rect 23432 22057 23478 22095
rect 23432 22023 23438 22057
rect 23472 22023 23478 22057
rect 23432 21985 23478 22023
rect 23432 21951 23438 21985
rect 23472 21951 23478 21985
rect 23432 21913 23478 21951
rect 23432 21879 23438 21913
rect 23472 21879 23478 21913
rect 23432 21841 23478 21879
rect 23432 21807 23438 21841
rect 23472 21807 23478 21841
rect 23432 21769 23478 21807
rect 23432 21735 23438 21769
rect 23472 21735 23478 21769
rect 23432 21697 23478 21735
rect 23432 21663 23438 21697
rect 23472 21663 23478 21697
rect 23432 21625 23478 21663
rect 23432 21591 23438 21625
rect 23472 21591 23478 21625
rect 23432 21553 23478 21591
rect 23432 21519 23438 21553
rect 23472 21519 23478 21553
rect 23432 21481 23478 21519
rect 23432 21447 23438 21481
rect 23472 21447 23478 21481
rect 23432 21409 23478 21447
rect 23432 21375 23438 21409
rect 23472 21375 23478 21409
rect 23432 21352 23478 21375
rect 23890 22129 23936 22152
rect 23890 22095 23896 22129
rect 23930 22095 23936 22129
rect 23890 22057 23936 22095
rect 23890 22023 23896 22057
rect 23930 22023 23936 22057
rect 23890 21985 23936 22023
rect 23890 21951 23896 21985
rect 23930 21951 23936 21985
rect 23890 21913 23936 21951
rect 23890 21879 23896 21913
rect 23930 21879 23936 21913
rect 23890 21841 23936 21879
rect 23890 21807 23896 21841
rect 23930 21807 23936 21841
rect 23890 21769 23936 21807
rect 23890 21735 23896 21769
rect 23930 21735 23936 21769
rect 23890 21697 23936 21735
rect 23890 21663 23896 21697
rect 23930 21663 23936 21697
rect 23890 21625 23936 21663
rect 23890 21591 23896 21625
rect 23930 21591 23936 21625
rect 23890 21553 23936 21591
rect 23890 21519 23896 21553
rect 23930 21519 23936 21553
rect 23890 21481 23936 21519
rect 23890 21447 23896 21481
rect 23930 21447 23936 21481
rect 23890 21409 23936 21447
rect 23890 21375 23896 21409
rect 23930 21375 23936 21409
rect 23890 21352 23936 21375
rect 24348 22129 24394 22152
rect 24348 22095 24354 22129
rect 24388 22095 24394 22129
rect 24348 22057 24394 22095
rect 24348 22023 24354 22057
rect 24388 22023 24394 22057
rect 24348 21985 24394 22023
rect 24348 21951 24354 21985
rect 24388 21951 24394 21985
rect 24348 21913 24394 21951
rect 24348 21879 24354 21913
rect 24388 21879 24394 21913
rect 24348 21841 24394 21879
rect 24348 21807 24354 21841
rect 24388 21807 24394 21841
rect 24348 21769 24394 21807
rect 24348 21735 24354 21769
rect 24388 21735 24394 21769
rect 24348 21697 24394 21735
rect 24348 21663 24354 21697
rect 24388 21663 24394 21697
rect 24348 21625 24394 21663
rect 24348 21591 24354 21625
rect 24388 21591 24394 21625
rect 24348 21553 24394 21591
rect 24348 21519 24354 21553
rect 24388 21519 24394 21553
rect 24348 21481 24394 21519
rect 24348 21447 24354 21481
rect 24388 21447 24394 21481
rect 24348 21409 24394 21447
rect 24348 21375 24354 21409
rect 24388 21375 24394 21409
rect 24348 21352 24394 21375
rect 24806 22129 24852 22152
rect 24806 22095 24812 22129
rect 24846 22095 24852 22129
rect 24806 22057 24852 22095
rect 24806 22023 24812 22057
rect 24846 22023 24852 22057
rect 24806 21985 24852 22023
rect 24806 21951 24812 21985
rect 24846 21951 24852 21985
rect 24806 21913 24852 21951
rect 24806 21879 24812 21913
rect 24846 21879 24852 21913
rect 24806 21841 24852 21879
rect 24806 21807 24812 21841
rect 24846 21807 24852 21841
rect 24806 21769 24852 21807
rect 24806 21735 24812 21769
rect 24846 21735 24852 21769
rect 24806 21697 24852 21735
rect 24806 21663 24812 21697
rect 24846 21663 24852 21697
rect 24806 21625 24852 21663
rect 24806 21591 24812 21625
rect 24846 21591 24852 21625
rect 24806 21553 24852 21591
rect 24806 21519 24812 21553
rect 24846 21519 24852 21553
rect 24806 21481 24852 21519
rect 24806 21447 24812 21481
rect 24846 21447 24852 21481
rect 24806 21409 24852 21447
rect 24806 21375 24812 21409
rect 24846 21375 24852 21409
rect 24806 21352 24852 21375
rect 25264 22129 25310 22152
rect 25264 22095 25270 22129
rect 25304 22095 25310 22129
rect 25264 22057 25310 22095
rect 25264 22023 25270 22057
rect 25304 22023 25310 22057
rect 25264 21985 25310 22023
rect 25264 21951 25270 21985
rect 25304 21951 25310 21985
rect 25264 21913 25310 21951
rect 25264 21879 25270 21913
rect 25304 21879 25310 21913
rect 25264 21841 25310 21879
rect 25264 21807 25270 21841
rect 25304 21807 25310 21841
rect 25264 21769 25310 21807
rect 25264 21735 25270 21769
rect 25304 21735 25310 21769
rect 25264 21697 25310 21735
rect 25264 21663 25270 21697
rect 25304 21663 25310 21697
rect 25264 21625 25310 21663
rect 25264 21591 25270 21625
rect 25304 21591 25310 21625
rect 25264 21553 25310 21591
rect 25264 21519 25270 21553
rect 25304 21519 25310 21553
rect 25264 21481 25310 21519
rect 25264 21447 25270 21481
rect 25304 21447 25310 21481
rect 25264 21409 25310 21447
rect 25264 21375 25270 21409
rect 25304 21375 25310 21409
rect 25264 21352 25310 21375
rect 25722 22129 25768 22152
rect 25722 22095 25728 22129
rect 25762 22095 25768 22129
rect 25722 22057 25768 22095
rect 25722 22023 25728 22057
rect 25762 22023 25768 22057
rect 25722 21985 25768 22023
rect 25722 21951 25728 21985
rect 25762 21951 25768 21985
rect 25722 21913 25768 21951
rect 25722 21879 25728 21913
rect 25762 21879 25768 21913
rect 25722 21841 25768 21879
rect 25722 21807 25728 21841
rect 25762 21807 25768 21841
rect 25722 21769 25768 21807
rect 25722 21735 25728 21769
rect 25762 21735 25768 21769
rect 25722 21697 25768 21735
rect 25722 21663 25728 21697
rect 25762 21663 25768 21697
rect 25722 21625 25768 21663
rect 25722 21591 25728 21625
rect 25762 21591 25768 21625
rect 25722 21553 25768 21591
rect 25722 21519 25728 21553
rect 25762 21519 25768 21553
rect 25722 21481 25768 21519
rect 25722 21447 25728 21481
rect 25762 21447 25768 21481
rect 25722 21409 25768 21447
rect 25722 21375 25728 21409
rect 25762 21375 25768 21409
rect 25722 21352 25768 21375
rect 26180 22129 26226 22152
rect 26180 22095 26186 22129
rect 26220 22095 26226 22129
rect 26180 22057 26226 22095
rect 26180 22023 26186 22057
rect 26220 22023 26226 22057
rect 26180 21985 26226 22023
rect 26180 21951 26186 21985
rect 26220 21951 26226 21985
rect 26180 21913 26226 21951
rect 26180 21879 26186 21913
rect 26220 21879 26226 21913
rect 26180 21841 26226 21879
rect 26180 21807 26186 21841
rect 26220 21807 26226 21841
rect 26180 21769 26226 21807
rect 26180 21735 26186 21769
rect 26220 21735 26226 21769
rect 26180 21697 26226 21735
rect 26180 21663 26186 21697
rect 26220 21663 26226 21697
rect 26180 21625 26226 21663
rect 26180 21591 26186 21625
rect 26220 21591 26226 21625
rect 26180 21553 26226 21591
rect 26180 21519 26186 21553
rect 26220 21519 26226 21553
rect 26180 21481 26226 21519
rect 26180 21447 26186 21481
rect 26220 21447 26226 21481
rect 26180 21409 26226 21447
rect 26180 21375 26186 21409
rect 26220 21375 26226 21409
rect 26180 21352 26226 21375
rect 26638 22129 26684 22152
rect 26638 22095 26644 22129
rect 26678 22095 26684 22129
rect 26638 22057 26684 22095
rect 26638 22023 26644 22057
rect 26678 22023 26684 22057
rect 26638 21985 26684 22023
rect 26638 21951 26644 21985
rect 26678 21951 26684 21985
rect 26638 21913 26684 21951
rect 26638 21879 26644 21913
rect 26678 21879 26684 21913
rect 26638 21841 26684 21879
rect 26638 21807 26644 21841
rect 26678 21807 26684 21841
rect 26638 21769 26684 21807
rect 26638 21735 26644 21769
rect 26678 21735 26684 21769
rect 26638 21697 26684 21735
rect 26638 21663 26644 21697
rect 26678 21663 26684 21697
rect 26638 21625 26684 21663
rect 26638 21591 26644 21625
rect 26678 21591 26684 21625
rect 26638 21553 26684 21591
rect 26638 21519 26644 21553
rect 26678 21519 26684 21553
rect 26638 21481 26684 21519
rect 26638 21447 26644 21481
rect 26678 21447 26684 21481
rect 26638 21409 26684 21447
rect 26638 21375 26644 21409
rect 26678 21375 26684 21409
rect 26638 21352 26684 21375
rect 27096 22129 27142 22152
rect 27096 22095 27102 22129
rect 27136 22095 27142 22129
rect 28450 22122 28470 22156
rect 28504 22122 28560 22156
rect 28594 22122 28650 22156
rect 28684 22122 28740 22156
rect 28774 22122 28830 22156
rect 28864 22122 28920 22156
rect 28954 22122 29010 22156
rect 29044 22122 29100 22156
rect 29134 22122 29190 22156
rect 29224 22122 29280 22156
rect 29314 22122 29370 22156
rect 29404 22122 29810 22156
rect 29844 22122 29900 22156
rect 29934 22122 29990 22156
rect 30024 22122 30080 22156
rect 30114 22122 30170 22156
rect 30204 22122 30260 22156
rect 30294 22122 30350 22156
rect 30384 22122 30440 22156
rect 30474 22122 30530 22156
rect 28450 22108 30564 22122
rect 30616 22156 38790 22160
rect 30616 22122 30620 22156
rect 30654 22122 30710 22156
rect 30744 22122 31150 22156
rect 31184 22122 31240 22156
rect 31274 22122 31330 22156
rect 31364 22122 31420 22156
rect 31454 22122 31510 22156
rect 31544 22122 31600 22156
rect 31634 22122 31690 22156
rect 31724 22122 31780 22156
rect 31814 22122 31870 22156
rect 31904 22122 31960 22156
rect 31994 22122 32050 22156
rect 32084 22122 32490 22156
rect 32524 22122 32580 22156
rect 32614 22122 32670 22156
rect 32704 22122 32760 22156
rect 32794 22122 32850 22156
rect 32884 22122 32940 22156
rect 32974 22122 33030 22156
rect 33064 22122 33120 22156
rect 33154 22122 33210 22156
rect 33244 22122 33300 22156
rect 33334 22122 33390 22156
rect 33424 22122 33830 22156
rect 33864 22122 33920 22156
rect 33954 22122 34010 22156
rect 34044 22122 34100 22156
rect 34134 22122 34190 22156
rect 34224 22122 34280 22156
rect 34314 22122 34370 22156
rect 34404 22122 34460 22156
rect 34494 22122 34550 22156
rect 34584 22122 34640 22156
rect 34674 22122 34730 22156
rect 34764 22122 35170 22156
rect 35204 22122 35260 22156
rect 35294 22122 35350 22156
rect 35384 22122 35440 22156
rect 35474 22122 35530 22156
rect 35564 22122 35620 22156
rect 35654 22122 35710 22156
rect 35744 22122 35800 22156
rect 35834 22122 35890 22156
rect 35924 22122 35980 22156
rect 36014 22122 36070 22156
rect 36104 22122 36510 22156
rect 36544 22122 36600 22156
rect 36634 22122 36690 22156
rect 36724 22122 36780 22156
rect 36814 22122 36870 22156
rect 36904 22122 36960 22156
rect 36994 22122 37050 22156
rect 37084 22122 37140 22156
rect 37174 22122 37230 22156
rect 37264 22122 37320 22156
rect 37354 22122 37410 22156
rect 37444 22122 37850 22156
rect 37884 22122 37940 22156
rect 37974 22122 38030 22156
rect 38064 22122 38120 22156
rect 38154 22122 38210 22156
rect 38244 22122 38300 22156
rect 38334 22122 38390 22156
rect 38424 22122 38480 22156
rect 38514 22122 38570 22156
rect 38604 22122 38660 22156
rect 38694 22122 38750 22156
rect 38784 22122 38790 22156
rect 30616 22108 38790 22122
rect 28450 22102 38790 22108
rect 27096 22057 27142 22095
rect 27096 22023 27102 22057
rect 27136 22023 27142 22057
rect 27096 21985 27142 22023
rect 28626 21998 28632 22024
rect 27096 21951 27102 21985
rect 27136 21951 27142 21985
rect 27096 21913 27142 21951
rect 27096 21879 27102 21913
rect 27136 21879 27142 21913
rect 27096 21841 27142 21879
rect 27096 21807 27102 21841
rect 27136 21807 27142 21841
rect 27096 21769 27142 21807
rect 27096 21735 27102 21769
rect 27136 21735 27142 21769
rect 27096 21697 27142 21735
rect 27096 21663 27102 21697
rect 27136 21663 27142 21697
rect 27096 21625 27142 21663
rect 27096 21591 27102 21625
rect 27136 21591 27142 21625
rect 27096 21553 27142 21591
rect 27096 21519 27102 21553
rect 27136 21519 27142 21553
rect 27096 21481 27142 21519
rect 27096 21447 27102 21481
rect 27136 21447 27142 21481
rect 27096 21409 27142 21447
rect 27096 21375 27102 21409
rect 27136 21375 27142 21409
rect 28624 21972 28632 21998
rect 28684 21998 28690 22024
rect 28684 21972 38616 21998
rect 28624 21952 38616 21972
rect 28624 21918 28656 21952
rect 28690 21918 28756 21952
rect 28790 21918 28856 21952
rect 28890 21918 28956 21952
rect 28990 21918 29056 21952
rect 29090 21918 29156 21952
rect 29190 21918 29996 21952
rect 30030 21918 30096 21952
rect 30130 21918 30196 21952
rect 30230 21918 30296 21952
rect 30330 21918 30396 21952
rect 30430 21918 30496 21952
rect 30530 21918 31336 21952
rect 31370 21918 31436 21952
rect 31470 21918 31536 21952
rect 31570 21918 31636 21952
rect 31670 21918 31736 21952
rect 31770 21918 31836 21952
rect 31870 21918 32676 21952
rect 32710 21918 32776 21952
rect 32810 21918 32876 21952
rect 32910 21918 32976 21952
rect 33010 21918 33076 21952
rect 33110 21918 33176 21952
rect 33210 21918 34016 21952
rect 34050 21918 34116 21952
rect 34150 21918 34216 21952
rect 34250 21918 34316 21952
rect 34350 21918 34416 21952
rect 34450 21918 34516 21952
rect 34550 21918 35356 21952
rect 35390 21918 35456 21952
rect 35490 21918 35556 21952
rect 35590 21918 35656 21952
rect 35690 21918 35756 21952
rect 35790 21918 35856 21952
rect 35890 21918 36696 21952
rect 36730 21918 36796 21952
rect 36830 21918 36896 21952
rect 36930 21918 36996 21952
rect 37030 21918 37096 21952
rect 37130 21918 37196 21952
rect 37230 21918 38036 21952
rect 38070 21918 38136 21952
rect 38170 21918 38236 21952
rect 38270 21918 38336 21952
rect 38370 21918 38436 21952
rect 38470 21918 38536 21952
rect 38570 21918 38616 21952
rect 28624 21852 38616 21918
rect 28624 21818 28656 21852
rect 28690 21818 28756 21852
rect 28790 21818 28856 21852
rect 28890 21818 28956 21852
rect 28990 21818 29056 21852
rect 29090 21818 29156 21852
rect 29190 21818 29996 21852
rect 30030 21818 30096 21852
rect 30130 21818 30196 21852
rect 30230 21818 30296 21852
rect 30330 21818 30396 21852
rect 30430 21818 30496 21852
rect 30530 21818 31336 21852
rect 31370 21818 31436 21852
rect 31470 21818 31536 21852
rect 31570 21818 31636 21852
rect 31670 21818 31736 21852
rect 31770 21818 31836 21852
rect 31870 21818 32676 21852
rect 32710 21818 32776 21852
rect 32810 21818 32876 21852
rect 32910 21818 32976 21852
rect 33010 21818 33076 21852
rect 33110 21818 33176 21852
rect 33210 21818 34016 21852
rect 34050 21818 34116 21852
rect 34150 21818 34216 21852
rect 34250 21818 34316 21852
rect 34350 21818 34416 21852
rect 34450 21818 34516 21852
rect 34550 21818 35356 21852
rect 35390 21818 35456 21852
rect 35490 21818 35556 21852
rect 35590 21818 35656 21852
rect 35690 21818 35756 21852
rect 35790 21818 35856 21852
rect 35890 21818 36696 21852
rect 36730 21818 36796 21852
rect 36830 21818 36896 21852
rect 36930 21818 36996 21852
rect 37030 21818 37096 21852
rect 37130 21818 37196 21852
rect 37230 21818 38036 21852
rect 38070 21818 38136 21852
rect 38170 21818 38236 21852
rect 38270 21818 38336 21852
rect 38370 21818 38436 21852
rect 38470 21818 38536 21852
rect 38570 21818 38616 21852
rect 39757 21843 39765 22324
rect 40159 21843 40167 22381
rect 39757 21831 40167 21843
rect 41765 22381 42175 22393
rect 41765 21843 41772 22381
rect 42166 21843 42175 22381
rect 41765 21831 42175 21843
rect 28624 21752 38616 21818
rect 28624 21718 28656 21752
rect 28690 21718 28756 21752
rect 28790 21718 28856 21752
rect 28890 21718 28956 21752
rect 28990 21718 29056 21752
rect 29090 21718 29156 21752
rect 29190 21718 29996 21752
rect 30030 21718 30096 21752
rect 30130 21718 30196 21752
rect 30230 21718 30296 21752
rect 30330 21718 30396 21752
rect 30430 21718 30496 21752
rect 30530 21718 31336 21752
rect 31370 21718 31436 21752
rect 31470 21718 31536 21752
rect 31570 21718 31636 21752
rect 31670 21718 31736 21752
rect 31770 21718 31836 21752
rect 31870 21718 32676 21752
rect 32710 21718 32776 21752
rect 32810 21718 32876 21752
rect 32910 21718 32976 21752
rect 33010 21718 33076 21752
rect 33110 21718 33176 21752
rect 33210 21718 34016 21752
rect 34050 21718 34116 21752
rect 34150 21718 34216 21752
rect 34250 21718 34316 21752
rect 34350 21718 34416 21752
rect 34450 21718 34516 21752
rect 34550 21718 35356 21752
rect 35390 21718 35456 21752
rect 35490 21718 35556 21752
rect 35590 21718 35656 21752
rect 35690 21718 35756 21752
rect 35790 21718 35856 21752
rect 35890 21718 36696 21752
rect 36730 21718 36796 21752
rect 36830 21718 36896 21752
rect 36930 21718 36996 21752
rect 37030 21718 37096 21752
rect 37130 21718 37196 21752
rect 37230 21718 38036 21752
rect 38070 21718 38136 21752
rect 38170 21718 38236 21752
rect 38270 21718 38336 21752
rect 38370 21718 38436 21752
rect 38470 21718 38536 21752
rect 38570 21718 38616 21752
rect 28624 21652 38616 21718
rect 28624 21618 28656 21652
rect 28690 21618 28756 21652
rect 28790 21618 28856 21652
rect 28890 21618 28956 21652
rect 28990 21618 29056 21652
rect 29090 21618 29156 21652
rect 29190 21618 29996 21652
rect 30030 21618 30096 21652
rect 30130 21618 30196 21652
rect 30230 21618 30296 21652
rect 30330 21618 30396 21652
rect 30430 21618 30496 21652
rect 30530 21618 31336 21652
rect 31370 21618 31436 21652
rect 31470 21618 31536 21652
rect 31570 21618 31636 21652
rect 31670 21618 31736 21652
rect 31770 21618 31836 21652
rect 31870 21618 32676 21652
rect 32710 21618 32776 21652
rect 32810 21618 32876 21652
rect 32910 21618 32976 21652
rect 33010 21618 33076 21652
rect 33110 21618 33176 21652
rect 33210 21618 34016 21652
rect 34050 21618 34116 21652
rect 34150 21618 34216 21652
rect 34250 21618 34316 21652
rect 34350 21618 34416 21652
rect 34450 21618 34516 21652
rect 34550 21618 35356 21652
rect 35390 21618 35456 21652
rect 35490 21618 35556 21652
rect 35590 21618 35656 21652
rect 35690 21618 35756 21652
rect 35790 21618 35856 21652
rect 35890 21618 36696 21652
rect 36730 21618 36796 21652
rect 36830 21618 36896 21652
rect 36930 21618 36996 21652
rect 37030 21618 37096 21652
rect 37130 21618 37196 21652
rect 37230 21618 38036 21652
rect 38070 21618 38136 21652
rect 38170 21618 38236 21652
rect 38270 21618 38336 21652
rect 38370 21618 38436 21652
rect 38470 21618 38536 21652
rect 38570 21618 38616 21652
rect 28624 21552 38616 21618
rect 28624 21518 28656 21552
rect 28690 21518 28756 21552
rect 28790 21518 28856 21552
rect 28890 21518 28956 21552
rect 28990 21518 29056 21552
rect 29090 21518 29156 21552
rect 29190 21518 29996 21552
rect 30030 21518 30096 21552
rect 30130 21518 30196 21552
rect 30230 21518 30296 21552
rect 30330 21518 30396 21552
rect 30430 21518 30496 21552
rect 30530 21518 31336 21552
rect 31370 21518 31436 21552
rect 31470 21518 31536 21552
rect 31570 21518 31636 21552
rect 31670 21518 31736 21552
rect 31770 21518 31836 21552
rect 31870 21518 32676 21552
rect 32710 21518 32776 21552
rect 32810 21518 32876 21552
rect 32910 21518 32976 21552
rect 33010 21518 33076 21552
rect 33110 21518 33176 21552
rect 33210 21518 34016 21552
rect 34050 21518 34116 21552
rect 34150 21518 34216 21552
rect 34250 21518 34316 21552
rect 34350 21518 34416 21552
rect 34450 21518 34516 21552
rect 34550 21518 35356 21552
rect 35390 21518 35456 21552
rect 35490 21518 35556 21552
rect 35590 21518 35656 21552
rect 35690 21518 35756 21552
rect 35790 21518 35856 21552
rect 35890 21518 36696 21552
rect 36730 21518 36796 21552
rect 36830 21518 36896 21552
rect 36930 21518 36996 21552
rect 37030 21518 37096 21552
rect 37130 21518 37196 21552
rect 37230 21518 38036 21552
rect 38070 21518 38136 21552
rect 38170 21518 38236 21552
rect 38270 21518 38336 21552
rect 38370 21518 38436 21552
rect 38470 21518 38536 21552
rect 38570 21518 38616 21552
rect 28624 21452 38616 21518
rect 28624 21418 28656 21452
rect 28690 21418 28756 21452
rect 28790 21418 28856 21452
rect 28890 21418 28956 21452
rect 28990 21418 29056 21452
rect 29090 21418 29156 21452
rect 29190 21418 29996 21452
rect 30030 21418 30096 21452
rect 30130 21418 30196 21452
rect 30230 21418 30296 21452
rect 30330 21418 30396 21452
rect 30430 21418 30496 21452
rect 30530 21418 31336 21452
rect 31370 21418 31436 21452
rect 31470 21418 31536 21452
rect 31570 21418 31636 21452
rect 31670 21418 31736 21452
rect 31770 21418 31836 21452
rect 31870 21418 32676 21452
rect 32710 21418 32776 21452
rect 32810 21418 32876 21452
rect 32910 21418 32976 21452
rect 33010 21418 33076 21452
rect 33110 21418 33176 21452
rect 33210 21418 34016 21452
rect 34050 21418 34116 21452
rect 34150 21418 34216 21452
rect 34250 21418 34316 21452
rect 34350 21418 34416 21452
rect 34450 21418 34516 21452
rect 34550 21418 35356 21452
rect 35390 21418 35456 21452
rect 35490 21418 35556 21452
rect 35590 21418 35656 21452
rect 35690 21418 35756 21452
rect 35790 21418 35856 21452
rect 35890 21418 36696 21452
rect 36730 21418 36796 21452
rect 36830 21418 36896 21452
rect 36930 21418 36996 21452
rect 37030 21418 37096 21452
rect 37130 21418 37196 21452
rect 37230 21418 38036 21452
rect 38070 21418 38136 21452
rect 38170 21418 38236 21452
rect 38270 21418 38336 21452
rect 38370 21418 38436 21452
rect 38470 21418 38536 21452
rect 38570 21418 38616 21452
rect 28624 21412 38616 21418
rect 28624 21386 28724 21412
rect 27096 21352 27142 21375
rect 28718 21360 28724 21386
rect 28776 21386 38616 21412
rect 39757 21421 40167 21433
rect 28776 21360 28782 21386
rect 13217 21301 13263 21339
rect 13217 21267 13223 21301
rect 13257 21267 13263 21301
rect 13217 21229 13263 21267
rect 13217 21195 13223 21229
rect 13257 21195 13263 21229
rect 21177 21267 21235 21273
rect 21177 21233 21189 21267
rect 21223 21233 21235 21267
rect 26510 21264 26516 21276
rect 26455 21236 26516 21264
rect 21177 21227 21235 21233
rect 13217 21157 13263 21195
rect 13217 21123 13223 21157
rect 13257 21123 13263 21157
rect 13217 21107 13263 21123
rect 21085 21131 21143 21137
rect 21085 21097 21097 21131
rect 21131 21128 21143 21131
rect 21192 21128 21220 21227
rect 26510 21224 26516 21236
rect 26568 21224 26574 21276
rect 30098 21156 30104 21208
rect 30156 21196 30162 21208
rect 39757 21196 39765 21421
rect 30156 21168 39765 21196
rect 30156 21156 30162 21168
rect 26878 21128 26884 21140
rect 21131 21100 21220 21128
rect 26823 21100 26884 21128
rect 21131 21097 21143 21100
rect 21085 21091 21143 21097
rect 13262 20992 13268 21004
rect 13207 20964 13268 20992
rect 13262 20952 13268 20964
rect 13320 20952 13326 21004
rect 8294 20884 8300 20936
rect 8352 20924 8358 20936
rect 8352 20896 8413 20924
rect 8352 20884 8358 20896
rect 21100 20812 21128 21091
rect 26878 21088 26884 21100
rect 26936 21088 26942 21140
rect 39757 20883 39765 21168
rect 40159 20883 40167 21421
rect 39757 20871 40167 20883
rect 41754 21421 42186 21831
rect 41754 20883 41772 21421
rect 42166 20883 42186 21421
rect 41754 20867 42186 20883
rect 900 20810 47736 20812
rect 900 20694 922 20810
rect 2510 20800 46126 20810
rect 2510 20769 14096 20800
rect 14148 20769 30564 20800
rect 2510 20735 7863 20769
rect 7897 20735 8263 20769
rect 8297 20735 8663 20769
rect 8697 20735 9063 20769
rect 9097 20735 9463 20769
rect 9497 20735 9863 20769
rect 9897 20735 10263 20769
rect 10297 20735 10663 20769
rect 10697 20735 11063 20769
rect 11097 20735 11463 20769
rect 11497 20735 11863 20769
rect 11897 20735 12263 20769
rect 12297 20735 12663 20769
rect 12697 20735 13063 20769
rect 13097 20735 13745 20769
rect 13779 20748 14096 20769
rect 13779 20735 14145 20748
rect 14179 20735 14545 20769
rect 14579 20735 14945 20769
rect 14979 20735 15345 20769
rect 15379 20735 15745 20769
rect 15779 20735 16145 20769
rect 16179 20735 16545 20769
rect 16579 20735 16945 20769
rect 16979 20735 17345 20769
rect 17379 20735 17745 20769
rect 17779 20735 18145 20769
rect 18179 20735 18545 20769
rect 18579 20735 18945 20769
rect 18979 20735 19345 20769
rect 19379 20735 19745 20769
rect 19779 20735 20145 20769
rect 20179 20735 20545 20769
rect 20579 20735 21191 20769
rect 21225 20735 21391 20769
rect 21425 20735 21591 20769
rect 21625 20735 21791 20769
rect 21825 20735 21991 20769
rect 22025 20735 22191 20769
rect 22225 20735 23151 20769
rect 23185 20735 23551 20769
rect 23585 20735 23951 20769
rect 23985 20735 24351 20769
rect 24385 20735 24751 20769
rect 24785 20735 25151 20769
rect 25185 20735 25551 20769
rect 25585 20735 25951 20769
rect 25985 20735 26351 20769
rect 26385 20735 26751 20769
rect 26785 20735 28443 20769
rect 28477 20735 28643 20769
rect 28677 20735 28843 20769
rect 28877 20735 29043 20769
rect 29077 20735 29243 20769
rect 29277 20735 29443 20769
rect 29477 20735 29643 20769
rect 29677 20735 29843 20769
rect 29877 20735 30043 20769
rect 30077 20735 30243 20769
rect 30277 20735 30443 20769
rect 30477 20748 30564 20769
rect 30616 20769 46126 20800
rect 30616 20748 30643 20769
rect 30477 20735 30643 20748
rect 30677 20735 30843 20769
rect 30877 20735 31043 20769
rect 31077 20735 31243 20769
rect 31277 20735 31443 20769
rect 31477 20735 31643 20769
rect 31677 20735 31843 20769
rect 31877 20735 32043 20769
rect 32077 20735 32243 20769
rect 32277 20735 32443 20769
rect 32477 20735 32643 20769
rect 32677 20735 32843 20769
rect 32877 20735 33043 20769
rect 33077 20735 33243 20769
rect 33277 20735 33443 20769
rect 33477 20735 33643 20769
rect 33677 20735 33843 20769
rect 33877 20735 34043 20769
rect 34077 20735 34243 20769
rect 34277 20735 34443 20769
rect 34477 20735 34643 20769
rect 34677 20735 34843 20769
rect 34877 20735 35043 20769
rect 35077 20735 35243 20769
rect 35277 20735 35443 20769
rect 35477 20735 35643 20769
rect 35677 20735 35843 20769
rect 35877 20735 36043 20769
rect 36077 20735 36243 20769
rect 36277 20735 36443 20769
rect 36477 20735 36643 20769
rect 36677 20735 36843 20769
rect 36877 20735 37043 20769
rect 37077 20735 37243 20769
rect 37277 20735 37443 20769
rect 37477 20735 37643 20769
rect 37677 20735 37843 20769
rect 37877 20735 38043 20769
rect 38077 20735 38243 20769
rect 38277 20735 38443 20769
rect 38477 20735 38643 20769
rect 38677 20735 38843 20769
rect 38877 20735 39929 20769
rect 39963 20735 40129 20769
rect 40163 20735 40329 20769
rect 40363 20735 40529 20769
rect 40563 20735 40729 20769
rect 40763 20735 40929 20769
rect 40963 20735 41129 20769
rect 41163 20735 41329 20769
rect 41363 20735 41529 20769
rect 41563 20735 41729 20769
rect 41763 20735 41929 20769
rect 41963 20735 46126 20769
rect 2510 20694 46126 20735
rect 47714 20694 47736 20810
rect 900 20692 47736 20694
rect 3348 18930 45288 18932
rect 3348 18814 3370 18930
rect 4958 18889 43678 18930
rect 4958 18855 6197 18889
rect 6231 18855 6597 18889
rect 6631 18855 6997 18889
rect 7031 18855 7397 18889
rect 7431 18855 7797 18889
rect 7831 18855 8197 18889
rect 8231 18855 8597 18889
rect 8631 18855 8997 18889
rect 9031 18855 9397 18889
rect 9431 18855 9797 18889
rect 9831 18855 10823 18889
rect 10857 18855 11023 18889
rect 11057 18855 11223 18889
rect 11257 18855 11423 18889
rect 11457 18855 11623 18889
rect 11657 18855 11823 18889
rect 11857 18855 12023 18889
rect 12057 18855 12223 18889
rect 12257 18855 12423 18889
rect 12457 18855 12623 18889
rect 12657 18855 12823 18889
rect 12857 18855 13567 18889
rect 13601 18855 13767 18889
rect 13801 18855 13967 18889
rect 14001 18855 14167 18889
rect 14201 18855 14367 18889
rect 14401 18855 14567 18889
rect 14601 18855 14767 18889
rect 14801 18855 14967 18889
rect 15001 18855 15167 18889
rect 15201 18855 15367 18889
rect 15401 18855 15567 18889
rect 15601 18855 16293 18889
rect 16327 18855 16693 18889
rect 16727 18855 17093 18889
rect 17127 18855 17493 18889
rect 17527 18855 17893 18889
rect 17927 18855 18293 18889
rect 18327 18855 18693 18889
rect 18727 18855 19093 18889
rect 19127 18855 19493 18889
rect 19527 18855 19893 18889
rect 19927 18855 20293 18889
rect 20327 18855 20693 18889
rect 20727 18855 21093 18889
rect 21127 18855 21493 18889
rect 21527 18855 21893 18889
rect 21927 18855 22293 18889
rect 22327 18855 22693 18889
rect 22727 18855 23093 18889
rect 23127 18855 24131 18889
rect 24165 18855 24531 18889
rect 24565 18855 24931 18889
rect 24965 18855 25331 18889
rect 25365 18855 25731 18889
rect 25765 18855 26131 18889
rect 26165 18855 26531 18889
rect 26565 18855 28443 18889
rect 28477 18855 28643 18889
rect 28677 18855 28843 18889
rect 28877 18855 29043 18889
rect 29077 18855 29243 18889
rect 29277 18855 29443 18889
rect 29477 18855 29643 18889
rect 29677 18855 29843 18889
rect 29877 18855 30043 18889
rect 30077 18855 30243 18889
rect 30277 18855 30443 18889
rect 30477 18855 30643 18889
rect 30677 18855 30843 18889
rect 30877 18855 31043 18889
rect 31077 18855 31243 18889
rect 31277 18855 31443 18889
rect 31477 18855 31643 18889
rect 31677 18855 31843 18889
rect 31877 18855 32043 18889
rect 32077 18855 32243 18889
rect 32277 18855 32443 18889
rect 32477 18855 32643 18889
rect 32677 18855 32843 18889
rect 32877 18855 33043 18889
rect 33077 18855 33243 18889
rect 33277 18855 33443 18889
rect 33477 18855 33643 18889
rect 33677 18855 33843 18889
rect 33877 18855 34043 18889
rect 34077 18855 34243 18889
rect 34277 18855 34443 18889
rect 34477 18855 34643 18889
rect 34677 18855 34843 18889
rect 34877 18855 35043 18889
rect 35077 18855 35243 18889
rect 35277 18855 35443 18889
rect 35477 18855 35643 18889
rect 35677 18855 35843 18889
rect 35877 18855 36043 18889
rect 36077 18855 36243 18889
rect 36277 18855 36443 18889
rect 36477 18855 36643 18889
rect 36677 18855 36843 18889
rect 36877 18855 37043 18889
rect 37077 18855 37243 18889
rect 37277 18855 37443 18889
rect 37477 18855 37643 18889
rect 37677 18855 37843 18889
rect 37877 18855 38043 18889
rect 38077 18855 38243 18889
rect 38277 18855 38443 18889
rect 38477 18855 38643 18889
rect 38677 18855 38843 18889
rect 38877 18855 39439 18889
rect 39473 18855 39639 18889
rect 39673 18855 39839 18889
rect 39873 18855 40039 18889
rect 40073 18855 40239 18889
rect 40273 18855 40439 18889
rect 40473 18855 40639 18889
rect 40673 18855 40839 18889
rect 40873 18855 41039 18889
rect 41073 18855 41239 18889
rect 41273 18855 41439 18889
rect 41473 18855 43678 18889
rect 4958 18814 43678 18855
rect 45266 18814 45288 18930
rect 3348 18812 45288 18814
rect 26160 18723 26188 18812
rect 26145 18717 26203 18723
rect 26145 18683 26157 18717
rect 26191 18683 26203 18717
rect 26145 18677 26203 18683
rect 10651 18621 11061 18633
rect 6020 18369 6066 18392
rect 6020 18335 6026 18369
rect 6060 18335 6066 18369
rect 6020 18297 6066 18335
rect 6020 18263 6026 18297
rect 6060 18263 6066 18297
rect 6020 18225 6066 18263
rect 6020 18191 6026 18225
rect 6060 18191 6066 18225
rect 6020 18153 6066 18191
rect 6020 18119 6026 18153
rect 6060 18119 6066 18153
rect 6020 18081 6066 18119
rect 6020 18047 6026 18081
rect 6060 18047 6066 18081
rect 6020 18009 6066 18047
rect 6020 17975 6026 18009
rect 6060 17975 6066 18009
rect 6020 17937 6066 17975
rect 6020 17903 6026 17937
rect 6060 17903 6066 17937
rect 6020 17865 6066 17903
rect 6020 17831 6026 17865
rect 6060 17831 6066 17865
rect 6020 17793 6066 17831
rect 6020 17759 6026 17793
rect 6060 17759 6066 17793
rect 6020 17721 6066 17759
rect 6020 17687 6026 17721
rect 6060 17687 6066 17721
rect 6020 17649 6066 17687
rect 6020 17615 6026 17649
rect 6060 17615 6066 17649
rect 6020 17592 6066 17615
rect 6478 18369 6524 18392
rect 6478 18335 6484 18369
rect 6518 18335 6524 18369
rect 6478 18297 6524 18335
rect 6478 18263 6484 18297
rect 6518 18263 6524 18297
rect 6478 18225 6524 18263
rect 6478 18191 6484 18225
rect 6518 18191 6524 18225
rect 6478 18153 6524 18191
rect 6478 18119 6484 18153
rect 6518 18119 6524 18153
rect 6478 18081 6524 18119
rect 6478 18047 6484 18081
rect 6518 18047 6524 18081
rect 6478 18009 6524 18047
rect 6478 17975 6484 18009
rect 6518 17975 6524 18009
rect 6478 17937 6524 17975
rect 6478 17903 6484 17937
rect 6518 17903 6524 17937
rect 6478 17865 6524 17903
rect 6478 17831 6484 17865
rect 6518 17831 6524 17865
rect 6478 17793 6524 17831
rect 6478 17759 6484 17793
rect 6518 17759 6524 17793
rect 6478 17721 6524 17759
rect 6478 17687 6484 17721
rect 6518 17687 6524 17721
rect 6478 17649 6524 17687
rect 6478 17615 6484 17649
rect 6518 17615 6524 17649
rect 6478 17592 6524 17615
rect 6936 18369 6982 18392
rect 6936 18335 6942 18369
rect 6976 18335 6982 18369
rect 6936 18297 6982 18335
rect 6936 18263 6942 18297
rect 6976 18263 6982 18297
rect 6936 18225 6982 18263
rect 6936 18191 6942 18225
rect 6976 18191 6982 18225
rect 6936 18153 6982 18191
rect 6936 18119 6942 18153
rect 6976 18119 6982 18153
rect 6936 18081 6982 18119
rect 6936 18047 6942 18081
rect 6976 18047 6982 18081
rect 6936 18009 6982 18047
rect 6936 17975 6942 18009
rect 6976 17975 6982 18009
rect 6936 17937 6982 17975
rect 6936 17903 6942 17937
rect 6976 17903 6982 17937
rect 6936 17865 6982 17903
rect 6936 17831 6942 17865
rect 6976 17831 6982 17865
rect 6936 17793 6982 17831
rect 6936 17759 6942 17793
rect 6976 17759 6982 17793
rect 6936 17721 6982 17759
rect 6936 17687 6942 17721
rect 6976 17687 6982 17721
rect 6936 17649 6982 17687
rect 6936 17615 6942 17649
rect 6976 17615 6982 17649
rect 6936 17592 6982 17615
rect 7394 18369 7440 18392
rect 7394 18335 7400 18369
rect 7434 18335 7440 18369
rect 7394 18297 7440 18335
rect 7394 18263 7400 18297
rect 7434 18263 7440 18297
rect 7394 18225 7440 18263
rect 7394 18191 7400 18225
rect 7434 18191 7440 18225
rect 7394 18153 7440 18191
rect 7394 18119 7400 18153
rect 7434 18119 7440 18153
rect 7394 18081 7440 18119
rect 7394 18047 7400 18081
rect 7434 18047 7440 18081
rect 7394 18009 7440 18047
rect 7394 17975 7400 18009
rect 7434 17975 7440 18009
rect 7394 17937 7440 17975
rect 7394 17903 7400 17937
rect 7434 17903 7440 17937
rect 7394 17865 7440 17903
rect 7394 17831 7400 17865
rect 7434 17831 7440 17865
rect 7394 17793 7440 17831
rect 7394 17759 7400 17793
rect 7434 17759 7440 17793
rect 7394 17721 7440 17759
rect 7394 17687 7400 17721
rect 7434 17687 7440 17721
rect 7394 17649 7440 17687
rect 7394 17615 7400 17649
rect 7434 17615 7440 17649
rect 7394 17592 7440 17615
rect 7852 18369 7898 18392
rect 7852 18335 7858 18369
rect 7892 18335 7898 18369
rect 7852 18297 7898 18335
rect 7852 18263 7858 18297
rect 7892 18263 7898 18297
rect 7852 18225 7898 18263
rect 7852 18191 7858 18225
rect 7892 18191 7898 18225
rect 7852 18153 7898 18191
rect 7852 18119 7858 18153
rect 7892 18119 7898 18153
rect 7852 18081 7898 18119
rect 7852 18047 7858 18081
rect 7892 18047 7898 18081
rect 7852 18009 7898 18047
rect 7852 17975 7858 18009
rect 7892 17975 7898 18009
rect 7852 17937 7898 17975
rect 7852 17903 7858 17937
rect 7892 17903 7898 17937
rect 7852 17865 7898 17903
rect 7852 17831 7858 17865
rect 7892 17831 7898 17865
rect 7852 17793 7898 17831
rect 7852 17759 7858 17793
rect 7892 17759 7898 17793
rect 7852 17721 7898 17759
rect 7852 17687 7858 17721
rect 7892 17687 7898 17721
rect 7852 17649 7898 17687
rect 7852 17615 7858 17649
rect 7892 17615 7898 17649
rect 7852 17592 7898 17615
rect 8310 18369 8356 18392
rect 8310 18335 8316 18369
rect 8350 18335 8356 18369
rect 8310 18297 8356 18335
rect 8310 18263 8316 18297
rect 8350 18263 8356 18297
rect 8310 18225 8356 18263
rect 8310 18191 8316 18225
rect 8350 18191 8356 18225
rect 8310 18153 8356 18191
rect 8310 18119 8316 18153
rect 8350 18119 8356 18153
rect 8310 18081 8356 18119
rect 8310 18047 8316 18081
rect 8350 18047 8356 18081
rect 8310 18009 8356 18047
rect 8310 17975 8316 18009
rect 8350 17975 8356 18009
rect 8310 17937 8356 17975
rect 8310 17903 8316 17937
rect 8350 17903 8356 17937
rect 8310 17865 8356 17903
rect 8310 17831 8316 17865
rect 8350 17831 8356 17865
rect 8310 17793 8356 17831
rect 8310 17759 8316 17793
rect 8350 17759 8356 17793
rect 8310 17721 8356 17759
rect 8310 17687 8316 17721
rect 8350 17687 8356 17721
rect 8310 17649 8356 17687
rect 8310 17615 8316 17649
rect 8350 17615 8356 17649
rect 8310 17592 8356 17615
rect 8768 18369 8814 18392
rect 8768 18335 8774 18369
rect 8808 18335 8814 18369
rect 8768 18297 8814 18335
rect 8768 18263 8774 18297
rect 8808 18263 8814 18297
rect 8768 18225 8814 18263
rect 8768 18191 8774 18225
rect 8808 18191 8814 18225
rect 8768 18153 8814 18191
rect 8768 18119 8774 18153
rect 8808 18119 8814 18153
rect 8768 18081 8814 18119
rect 8768 18047 8774 18081
rect 8808 18047 8814 18081
rect 8768 18009 8814 18047
rect 8768 17975 8774 18009
rect 8808 17975 8814 18009
rect 8768 17937 8814 17975
rect 8768 17903 8774 17937
rect 8808 17903 8814 17937
rect 8768 17865 8814 17903
rect 8768 17831 8774 17865
rect 8808 17831 8814 17865
rect 8768 17793 8814 17831
rect 8768 17759 8774 17793
rect 8808 17759 8814 17793
rect 8768 17721 8814 17759
rect 8768 17687 8774 17721
rect 8808 17687 8814 17721
rect 8768 17649 8814 17687
rect 8768 17615 8774 17649
rect 8808 17615 8814 17649
rect 8768 17592 8814 17615
rect 9226 18369 9272 18392
rect 9226 18335 9232 18369
rect 9266 18335 9272 18369
rect 9684 18369 9730 18392
rect 9684 18352 9690 18369
rect 9724 18352 9730 18369
rect 10142 18369 10188 18392
rect 9226 18297 9272 18335
rect 9674 18300 9680 18352
rect 9732 18300 9738 18352
rect 10142 18335 10148 18369
rect 10182 18335 10188 18369
rect 9226 18263 9232 18297
rect 9266 18263 9272 18297
rect 9226 18225 9272 18263
rect 9226 18191 9232 18225
rect 9266 18191 9272 18225
rect 9226 18153 9272 18191
rect 9226 18119 9232 18153
rect 9266 18119 9272 18153
rect 9226 18081 9272 18119
rect 9226 18047 9232 18081
rect 9266 18047 9272 18081
rect 9226 18009 9272 18047
rect 9226 17975 9232 18009
rect 9266 17975 9272 18009
rect 9226 17937 9272 17975
rect 9226 17903 9232 17937
rect 9266 17903 9272 17937
rect 9226 17865 9272 17903
rect 9226 17831 9232 17865
rect 9266 17831 9272 17865
rect 9226 17793 9272 17831
rect 9226 17759 9232 17793
rect 9266 17759 9272 17793
rect 9226 17721 9272 17759
rect 9226 17687 9232 17721
rect 9266 17687 9272 17721
rect 9226 17649 9272 17687
rect 9226 17615 9232 17649
rect 9266 17615 9272 17649
rect 9226 17592 9272 17615
rect 9684 18297 9730 18300
rect 9684 18263 9690 18297
rect 9724 18263 9730 18297
rect 9684 18225 9730 18263
rect 9684 18191 9690 18225
rect 9724 18191 9730 18225
rect 9684 18153 9730 18191
rect 9684 18119 9690 18153
rect 9724 18119 9730 18153
rect 9684 18081 9730 18119
rect 9684 18047 9690 18081
rect 9724 18047 9730 18081
rect 9684 18009 9730 18047
rect 9684 17975 9690 18009
rect 9724 17975 9730 18009
rect 9684 17937 9730 17975
rect 9684 17903 9690 17937
rect 9724 17903 9730 17937
rect 9684 17865 9730 17903
rect 9684 17831 9690 17865
rect 9724 17831 9730 17865
rect 9684 17793 9730 17831
rect 9684 17759 9690 17793
rect 9724 17759 9730 17793
rect 9684 17721 9730 17759
rect 9684 17687 9690 17721
rect 9724 17687 9730 17721
rect 9684 17649 9730 17687
rect 9684 17615 9690 17649
rect 9724 17615 9730 17649
rect 9684 17592 9730 17615
rect 10142 18297 10188 18335
rect 10142 18263 10148 18297
rect 10182 18263 10188 18297
rect 10142 18225 10188 18263
rect 10142 18191 10148 18225
rect 10182 18191 10188 18225
rect 10142 18153 10188 18191
rect 10142 18119 10148 18153
rect 10182 18119 10188 18153
rect 10142 18081 10188 18119
rect 10142 18047 10148 18081
rect 10182 18047 10188 18081
rect 10651 18083 10659 18621
rect 11053 18136 11061 18621
rect 12659 18621 13069 18633
rect 13395 18624 13805 18633
rect 12526 18136 12532 18148
rect 11053 18108 12532 18136
rect 11053 18083 11061 18108
rect 12526 18096 12532 18108
rect 12584 18096 12590 18148
rect 10651 18071 11061 18083
rect 12659 18083 12666 18621
rect 13060 18083 13069 18621
rect 13354 18572 13360 18624
rect 13412 18621 13805 18624
rect 12659 18071 13069 18083
rect 13395 18083 13403 18572
rect 13797 18083 13805 18621
rect 13395 18071 13805 18083
rect 15403 18621 15813 18633
rect 15403 18083 15410 18621
rect 15804 18083 15813 18621
rect 15403 18071 15813 18083
rect 23989 18621 24035 18637
rect 23989 18587 23995 18621
rect 24029 18587 24035 18621
rect 23989 18549 24035 18587
rect 23989 18515 23995 18549
rect 24029 18515 24035 18549
rect 23989 18477 24035 18515
rect 23989 18443 23995 18477
rect 24029 18443 24035 18477
rect 23989 18405 24035 18443
rect 23989 18371 23995 18405
rect 24029 18371 24035 18405
rect 23989 18333 24035 18371
rect 23989 18299 23995 18333
rect 24029 18299 24035 18333
rect 23989 18261 24035 18299
rect 23989 18227 23995 18261
rect 24029 18227 24035 18261
rect 23989 18189 24035 18227
rect 23989 18155 23995 18189
rect 24029 18155 24035 18189
rect 23989 18117 24035 18155
rect 23989 18083 23995 18117
rect 24029 18083 24035 18117
rect 10142 18009 10188 18047
rect 10142 17975 10148 18009
rect 10182 17975 10188 18009
rect 10142 17937 10188 17975
rect 10142 17903 10148 17937
rect 10182 17903 10188 17937
rect 10142 17865 10188 17903
rect 10142 17831 10148 17865
rect 10182 17831 10188 17865
rect 10142 17793 10188 17831
rect 10142 17759 10148 17793
rect 10182 17759 10188 17793
rect 10142 17721 10188 17759
rect 10142 17687 10148 17721
rect 10182 17687 10188 17721
rect 10142 17649 10188 17687
rect 10142 17615 10148 17649
rect 10182 17615 10188 17649
rect 10142 17592 10188 17615
rect 10651 17661 11061 17673
rect 6089 17323 6147 17329
rect 6089 17320 6101 17323
rect 0 17292 6101 17320
rect 6089 17289 6101 17292
rect 6135 17289 6147 17323
rect 6089 17283 6147 17289
rect 8312 17052 8340 17592
rect 8754 17144 8760 17196
rect 8812 17184 8818 17196
rect 10651 17184 10659 17661
rect 8812 17156 10659 17184
rect 8812 17144 8818 17156
rect 10651 17123 10659 17156
rect 11053 17123 11061 17661
rect 10651 17111 11061 17123
rect 12648 17661 13080 18071
rect 12648 17123 12666 17661
rect 13060 17123 13080 17661
rect 13170 17620 13176 17672
rect 13228 17660 13234 17672
rect 13395 17661 13805 17673
rect 13395 17660 13403 17661
rect 13228 17632 13403 17660
rect 13228 17620 13234 17632
rect 12648 17107 13080 17123
rect 13395 17123 13403 17632
rect 13797 17123 13805 17661
rect 13395 17111 13805 17123
rect 15392 17661 15824 18071
rect 15392 17123 15410 17661
rect 15804 17123 15824 17661
rect 23989 18045 24035 18083
rect 23989 18011 23995 18045
rect 24029 18011 24035 18045
rect 23989 17973 24035 18011
rect 23989 17939 23995 17973
rect 24029 17939 24035 17973
rect 23989 17901 24035 17939
rect 23989 17867 23995 17901
rect 24029 17867 24035 17901
rect 23989 17829 24035 17867
rect 23989 17795 23995 17829
rect 24029 17795 24035 17829
rect 23989 17757 24035 17795
rect 23989 17723 23995 17757
rect 24029 17723 24035 17757
rect 23989 17685 24035 17723
rect 23989 17651 23995 17685
rect 24029 17651 24035 17685
rect 23989 17613 24035 17651
rect 23989 17579 23995 17613
rect 24029 17579 24035 17613
rect 23989 17541 24035 17579
rect 23989 17507 23995 17541
rect 24029 17507 24035 17541
rect 23989 17469 24035 17507
rect 23989 17435 23995 17469
rect 24029 17435 24035 17469
rect 23989 17397 24035 17435
rect 23989 17363 23995 17397
rect 24029 17363 24035 17397
rect 23989 17347 24035 17363
rect 24447 18621 24493 18637
rect 24447 18587 24453 18621
rect 24487 18587 24493 18621
rect 24447 18549 24493 18587
rect 24447 18515 24453 18549
rect 24487 18515 24493 18549
rect 24447 18477 24493 18515
rect 24447 18443 24453 18477
rect 24487 18443 24493 18477
rect 24447 18405 24493 18443
rect 24447 18371 24453 18405
rect 24487 18371 24493 18405
rect 24447 18333 24493 18371
rect 24447 18299 24453 18333
rect 24487 18299 24493 18333
rect 24447 18261 24493 18299
rect 24447 18227 24453 18261
rect 24487 18227 24493 18261
rect 24447 18189 24493 18227
rect 24447 18155 24453 18189
rect 24487 18155 24493 18189
rect 24447 18117 24493 18155
rect 24447 18083 24453 18117
rect 24487 18083 24493 18117
rect 24447 18045 24493 18083
rect 24447 18011 24453 18045
rect 24487 18011 24493 18045
rect 24447 17973 24493 18011
rect 24447 17939 24453 17973
rect 24487 17939 24493 17973
rect 24447 17901 24493 17939
rect 24447 17867 24453 17901
rect 24487 17867 24493 17901
rect 24447 17829 24493 17867
rect 24447 17795 24453 17829
rect 24487 17795 24493 17829
rect 24447 17757 24493 17795
rect 24447 17723 24453 17757
rect 24487 17723 24493 17757
rect 24447 17685 24493 17723
rect 24447 17651 24453 17685
rect 24487 17651 24493 17685
rect 24447 17613 24493 17651
rect 24447 17579 24453 17613
rect 24487 17579 24493 17613
rect 24447 17541 24493 17579
rect 24447 17507 24453 17541
rect 24487 17507 24493 17541
rect 24447 17469 24493 17507
rect 24447 17435 24453 17469
rect 24487 17435 24493 17469
rect 24447 17397 24493 17435
rect 24447 17363 24453 17397
rect 24487 17363 24493 17397
rect 24447 17347 24493 17363
rect 24905 18621 24951 18637
rect 24905 18587 24911 18621
rect 24945 18587 24951 18621
rect 24905 18549 24951 18587
rect 24905 18515 24911 18549
rect 24945 18515 24951 18549
rect 24905 18477 24951 18515
rect 24905 18443 24911 18477
rect 24945 18443 24951 18477
rect 24905 18405 24951 18443
rect 24905 18371 24911 18405
rect 24945 18371 24951 18405
rect 24905 18333 24951 18371
rect 24905 18299 24911 18333
rect 24945 18299 24951 18333
rect 24905 18261 24951 18299
rect 24905 18227 24911 18261
rect 24945 18227 24951 18261
rect 24905 18189 24951 18227
rect 24905 18155 24911 18189
rect 24945 18155 24951 18189
rect 24905 18117 24951 18155
rect 24905 18083 24911 18117
rect 24945 18083 24951 18117
rect 24905 18045 24951 18083
rect 24905 18011 24911 18045
rect 24945 18011 24951 18045
rect 24905 17973 24951 18011
rect 24905 17939 24911 17973
rect 24945 17939 24951 17973
rect 24905 17901 24951 17939
rect 24905 17867 24911 17901
rect 24945 17867 24951 17901
rect 24905 17829 24951 17867
rect 24905 17795 24911 17829
rect 24945 17795 24951 17829
rect 24905 17757 24951 17795
rect 24905 17723 24911 17757
rect 24945 17723 24951 17757
rect 24905 17685 24951 17723
rect 24905 17651 24911 17685
rect 24945 17651 24951 17685
rect 24905 17613 24951 17651
rect 24905 17579 24911 17613
rect 24945 17579 24951 17613
rect 24905 17541 24951 17579
rect 24905 17507 24911 17541
rect 24945 17507 24951 17541
rect 24905 17469 24951 17507
rect 24905 17435 24911 17469
rect 24945 17435 24951 17469
rect 24905 17397 24951 17435
rect 24905 17363 24911 17397
rect 24945 17363 24951 17397
rect 24905 17347 24951 17363
rect 25363 18621 25409 18637
rect 25363 18587 25369 18621
rect 25403 18587 25409 18621
rect 25363 18549 25409 18587
rect 25363 18515 25369 18549
rect 25403 18515 25409 18549
rect 25363 18477 25409 18515
rect 25363 18443 25369 18477
rect 25403 18443 25409 18477
rect 25363 18405 25409 18443
rect 25363 18371 25369 18405
rect 25403 18371 25409 18405
rect 25363 18333 25409 18371
rect 25363 18299 25369 18333
rect 25403 18299 25409 18333
rect 25363 18261 25409 18299
rect 25363 18227 25369 18261
rect 25403 18227 25409 18261
rect 25363 18189 25409 18227
rect 25363 18155 25369 18189
rect 25403 18155 25409 18189
rect 25363 18117 25409 18155
rect 25363 18083 25369 18117
rect 25403 18083 25409 18117
rect 25363 18045 25409 18083
rect 25363 18011 25369 18045
rect 25403 18011 25409 18045
rect 25363 17973 25409 18011
rect 25363 17939 25369 17973
rect 25403 17939 25409 17973
rect 25363 17901 25409 17939
rect 25363 17867 25369 17901
rect 25403 17867 25409 17901
rect 25363 17829 25409 17867
rect 25363 17795 25369 17829
rect 25403 17795 25409 17829
rect 25363 17757 25409 17795
rect 25363 17723 25369 17757
rect 25403 17723 25409 17757
rect 25363 17685 25409 17723
rect 25363 17651 25369 17685
rect 25403 17651 25409 17685
rect 25363 17613 25409 17651
rect 25363 17579 25369 17613
rect 25403 17579 25409 17613
rect 25363 17541 25409 17579
rect 25363 17507 25369 17541
rect 25403 17507 25409 17541
rect 25363 17469 25409 17507
rect 25363 17435 25369 17469
rect 25403 17435 25409 17469
rect 25363 17397 25409 17435
rect 25363 17363 25369 17397
rect 25403 17363 25409 17397
rect 25363 17347 25409 17363
rect 25821 18621 25867 18637
rect 25821 18587 25827 18621
rect 25861 18587 25867 18621
rect 25821 18549 25867 18587
rect 25821 18515 25827 18549
rect 25861 18515 25867 18549
rect 25821 18477 25867 18515
rect 25821 18443 25827 18477
rect 25861 18443 25867 18477
rect 25821 18405 25867 18443
rect 25821 18371 25827 18405
rect 25861 18371 25867 18405
rect 25821 18333 25867 18371
rect 25821 18299 25827 18333
rect 25861 18299 25867 18333
rect 25821 18261 25867 18299
rect 25821 18227 25827 18261
rect 25861 18227 25867 18261
rect 25821 18189 25867 18227
rect 25821 18155 25827 18189
rect 25861 18155 25867 18189
rect 25821 18117 25867 18155
rect 25821 18083 25827 18117
rect 25861 18083 25867 18117
rect 25821 18045 25867 18083
rect 25821 18011 25827 18045
rect 25861 18011 25867 18045
rect 25821 17973 25867 18011
rect 25821 17939 25827 17973
rect 25861 17939 25867 17973
rect 25821 17901 25867 17939
rect 25821 17867 25827 17901
rect 25861 17867 25867 17901
rect 25821 17829 25867 17867
rect 25821 17795 25827 17829
rect 25861 17795 25867 17829
rect 25821 17757 25867 17795
rect 25821 17723 25827 17757
rect 25861 17723 25867 17757
rect 25821 17685 25867 17723
rect 25821 17651 25827 17685
rect 25861 17651 25867 17685
rect 25821 17613 25867 17651
rect 25821 17579 25827 17613
rect 25861 17579 25867 17613
rect 25821 17541 25867 17579
rect 25821 17507 25827 17541
rect 25861 17507 25867 17541
rect 25821 17469 25867 17507
rect 25821 17435 25827 17469
rect 25861 17435 25867 17469
rect 25821 17397 25867 17435
rect 25821 17363 25827 17397
rect 25861 17363 25867 17397
rect 25821 17347 25867 17363
rect 26279 18621 26325 18637
rect 26279 18587 26285 18621
rect 26319 18587 26325 18621
rect 26279 18549 26325 18587
rect 26279 18515 26285 18549
rect 26319 18515 26325 18549
rect 26279 18477 26325 18515
rect 26279 18443 26285 18477
rect 26319 18443 26325 18477
rect 26279 18405 26325 18443
rect 26279 18371 26285 18405
rect 26319 18371 26325 18405
rect 26279 18333 26325 18371
rect 26279 18299 26285 18333
rect 26319 18299 26325 18333
rect 26279 18261 26325 18299
rect 26279 18227 26285 18261
rect 26319 18227 26325 18261
rect 26279 18189 26325 18227
rect 26279 18155 26285 18189
rect 26319 18155 26325 18189
rect 26279 18117 26325 18155
rect 26279 18083 26285 18117
rect 26319 18083 26325 18117
rect 26279 18045 26325 18083
rect 26279 18011 26285 18045
rect 26319 18011 26325 18045
rect 26279 17973 26325 18011
rect 26279 17939 26285 17973
rect 26319 17939 26325 17973
rect 26279 17901 26325 17939
rect 26279 17867 26285 17901
rect 26319 17867 26325 17901
rect 26279 17829 26325 17867
rect 26279 17795 26285 17829
rect 26319 17795 26325 17829
rect 26279 17757 26325 17795
rect 26279 17723 26285 17757
rect 26319 17723 26325 17757
rect 26279 17685 26325 17723
rect 26279 17651 26285 17685
rect 26319 17651 26325 17685
rect 26279 17613 26325 17651
rect 26279 17579 26285 17613
rect 26319 17579 26325 17613
rect 26279 17541 26325 17579
rect 26279 17507 26285 17541
rect 26319 17507 26325 17541
rect 26279 17469 26325 17507
rect 26279 17435 26285 17469
rect 26319 17435 26325 17469
rect 26279 17397 26325 17435
rect 26279 17363 26285 17397
rect 26319 17363 26325 17397
rect 26279 17347 26325 17363
rect 26737 18621 26783 18637
rect 26737 18587 26743 18621
rect 26777 18587 26783 18621
rect 26737 18549 26783 18587
rect 39267 18624 39677 18633
rect 39267 18621 39488 18624
rect 39540 18621 39677 18624
rect 26737 18515 26743 18549
rect 26777 18515 26783 18549
rect 26737 18477 26783 18515
rect 28286 18556 38954 18562
rect 28286 18522 28306 18556
rect 28340 18522 28396 18556
rect 28430 18522 28486 18556
rect 28520 18522 28576 18556
rect 28610 18522 28666 18556
rect 28700 18522 28756 18556
rect 28790 18522 28846 18556
rect 28880 18522 28936 18556
rect 28970 18522 29026 18556
rect 29060 18522 29116 18556
rect 29150 18522 29206 18556
rect 29240 18522 29296 18556
rect 29330 18522 29386 18556
rect 29420 18522 29476 18556
rect 29510 18522 29646 18556
rect 29680 18522 29736 18556
rect 29770 18522 29826 18556
rect 29860 18522 29916 18556
rect 29950 18522 30006 18556
rect 30040 18522 30096 18556
rect 30130 18522 30186 18556
rect 30220 18522 30276 18556
rect 30310 18522 30366 18556
rect 30400 18522 30456 18556
rect 30490 18522 30546 18556
rect 30580 18522 30636 18556
rect 30670 18522 30726 18556
rect 30760 18522 30816 18556
rect 30850 18522 30986 18556
rect 31020 18522 31076 18556
rect 31110 18522 31166 18556
rect 31200 18522 31256 18556
rect 31290 18522 31346 18556
rect 31380 18522 31436 18556
rect 31470 18522 31526 18556
rect 31560 18522 31616 18556
rect 31650 18522 31706 18556
rect 31740 18522 31796 18556
rect 31830 18522 31886 18556
rect 31920 18522 31976 18556
rect 32010 18522 32066 18556
rect 32100 18522 32156 18556
rect 32190 18522 32326 18556
rect 32360 18522 32416 18556
rect 32450 18522 32506 18556
rect 32540 18522 32596 18556
rect 32630 18522 32686 18556
rect 32720 18522 32776 18556
rect 32810 18522 32866 18556
rect 32900 18522 32956 18556
rect 32990 18522 33046 18556
rect 33080 18522 33136 18556
rect 33170 18522 33226 18556
rect 33260 18522 33316 18556
rect 33350 18522 33406 18556
rect 33440 18522 33496 18556
rect 33530 18522 33666 18556
rect 33700 18522 33756 18556
rect 33790 18522 33846 18556
rect 33880 18522 33936 18556
rect 33970 18522 34026 18556
rect 34060 18522 34116 18556
rect 34150 18522 34206 18556
rect 34240 18522 34296 18556
rect 34330 18522 34386 18556
rect 34420 18522 34476 18556
rect 34510 18522 34566 18556
rect 34600 18522 34656 18556
rect 34690 18522 34746 18556
rect 34780 18522 34836 18556
rect 34870 18522 35006 18556
rect 35040 18522 35096 18556
rect 35130 18522 35186 18556
rect 35220 18522 35276 18556
rect 35310 18522 35366 18556
rect 35400 18522 35456 18556
rect 35490 18522 35546 18556
rect 35580 18522 35636 18556
rect 35670 18522 35726 18556
rect 35760 18522 35816 18556
rect 35850 18522 35906 18556
rect 35940 18522 35996 18556
rect 36030 18522 36086 18556
rect 36120 18522 36176 18556
rect 36210 18522 36346 18556
rect 36380 18522 36436 18556
rect 36470 18522 36526 18556
rect 36560 18522 36616 18556
rect 36650 18522 36706 18556
rect 36740 18522 36796 18556
rect 36830 18522 36886 18556
rect 36920 18522 36976 18556
rect 37010 18522 37066 18556
rect 37100 18522 37156 18556
rect 37190 18522 37246 18556
rect 37280 18522 37336 18556
rect 37370 18522 37426 18556
rect 37460 18522 37516 18556
rect 37550 18522 37686 18556
rect 37720 18522 37776 18556
rect 37810 18522 37866 18556
rect 37900 18522 37956 18556
rect 37990 18522 38046 18556
rect 38080 18522 38136 18556
rect 38170 18522 38226 18556
rect 38260 18522 38316 18556
rect 38350 18522 38406 18556
rect 38440 18522 38496 18556
rect 38530 18522 38586 18556
rect 38620 18522 38676 18556
rect 38710 18522 38766 18556
rect 38800 18522 38856 18556
rect 38890 18522 38954 18556
rect 28286 18492 38954 18522
rect 26737 18443 26743 18477
rect 26777 18443 26783 18477
rect 26737 18405 26783 18443
rect 28626 18412 28632 18420
rect 26737 18371 26743 18405
rect 26777 18371 26783 18405
rect 26737 18333 26783 18371
rect 28450 18396 28632 18412
rect 28684 18412 28690 18420
rect 34440 18412 34468 18492
rect 28684 18396 38790 18412
rect 28450 18362 28470 18396
rect 28504 18362 28560 18396
rect 28594 18368 28632 18396
rect 28594 18362 28650 18368
rect 28684 18362 28740 18396
rect 28774 18362 28830 18396
rect 28864 18362 28920 18396
rect 28954 18362 29010 18396
rect 29044 18362 29100 18396
rect 29134 18362 29190 18396
rect 29224 18362 29280 18396
rect 29314 18362 29370 18396
rect 29404 18362 29810 18396
rect 29844 18362 29900 18396
rect 29934 18362 29990 18396
rect 30024 18362 30080 18396
rect 30114 18362 30170 18396
rect 30204 18362 30260 18396
rect 30294 18362 30350 18396
rect 30384 18362 30440 18396
rect 30474 18362 30530 18396
rect 30564 18362 30620 18396
rect 30654 18362 30710 18396
rect 30744 18362 31150 18396
rect 31184 18362 31240 18396
rect 31274 18362 31330 18396
rect 31364 18362 31420 18396
rect 31454 18362 31510 18396
rect 31544 18362 31600 18396
rect 31634 18362 31690 18396
rect 31724 18362 31780 18396
rect 31814 18362 31870 18396
rect 31904 18362 31960 18396
rect 31994 18362 32050 18396
rect 32084 18362 32490 18396
rect 32524 18362 32580 18396
rect 32614 18362 32670 18396
rect 32704 18362 32760 18396
rect 32794 18362 32850 18396
rect 32884 18362 32940 18396
rect 32974 18362 33030 18396
rect 33064 18362 33120 18396
rect 33154 18362 33210 18396
rect 33244 18362 33300 18396
rect 33334 18362 33390 18396
rect 33424 18362 33830 18396
rect 33864 18362 33920 18396
rect 33954 18362 34010 18396
rect 34044 18362 34100 18396
rect 34134 18362 34190 18396
rect 34224 18362 34280 18396
rect 34314 18362 34370 18396
rect 34404 18362 34460 18396
rect 34494 18362 34550 18396
rect 34584 18362 34640 18396
rect 34674 18362 34730 18396
rect 34764 18362 35170 18396
rect 35204 18362 35260 18396
rect 35294 18362 35350 18396
rect 35384 18362 35440 18396
rect 35474 18362 35530 18396
rect 35564 18362 35620 18396
rect 35654 18362 35710 18396
rect 35744 18362 35800 18396
rect 35834 18362 35890 18396
rect 35924 18362 35980 18396
rect 36014 18362 36070 18396
rect 36104 18362 36510 18396
rect 36544 18362 36600 18396
rect 36634 18362 36690 18396
rect 36724 18362 36780 18396
rect 36814 18362 36870 18396
rect 36904 18362 36960 18396
rect 36994 18362 37050 18396
rect 37084 18362 37140 18396
rect 37174 18362 37230 18396
rect 37264 18362 37320 18396
rect 37354 18362 37410 18396
rect 37444 18362 37850 18396
rect 37884 18362 37940 18396
rect 37974 18362 38030 18396
rect 38064 18362 38120 18396
rect 38154 18362 38210 18396
rect 38244 18362 38300 18396
rect 38334 18362 38390 18396
rect 38424 18362 38480 18396
rect 38514 18362 38570 18396
rect 38604 18362 38660 18396
rect 38694 18362 38750 18396
rect 38784 18362 38790 18396
rect 28450 18342 38790 18362
rect 26737 18299 26743 18333
rect 26777 18299 26783 18333
rect 26737 18261 26783 18299
rect 26737 18227 26743 18261
rect 26777 18227 26783 18261
rect 26737 18189 26783 18227
rect 26737 18155 26743 18189
rect 26777 18155 26783 18189
rect 26737 18117 26783 18155
rect 26737 18083 26743 18117
rect 26777 18083 26783 18117
rect 26737 18045 26783 18083
rect 26737 18011 26743 18045
rect 26777 18011 26783 18045
rect 26737 17973 26783 18011
rect 26737 17939 26743 17973
rect 26777 17939 26783 17973
rect 26737 17901 26783 17939
rect 26737 17867 26743 17901
rect 26777 17867 26783 17901
rect 26737 17829 26783 17867
rect 26737 17795 26743 17829
rect 26777 17795 26783 17829
rect 26737 17757 26783 17795
rect 26737 17723 26743 17757
rect 26777 17723 26783 17757
rect 26737 17685 26783 17723
rect 26737 17651 26743 17685
rect 26777 17651 26783 17685
rect 26737 17613 26783 17651
rect 28624 18216 38616 18238
rect 28624 18192 28724 18216
rect 28776 18192 38616 18216
rect 28624 18158 28656 18192
rect 28690 18164 28724 18192
rect 28690 18158 28756 18164
rect 28790 18158 28856 18192
rect 28890 18158 28956 18192
rect 28990 18158 29056 18192
rect 29090 18158 29156 18192
rect 29190 18158 29996 18192
rect 30030 18158 30096 18192
rect 30130 18158 30196 18192
rect 30230 18158 30296 18192
rect 30330 18158 30396 18192
rect 30430 18158 30496 18192
rect 30530 18158 31336 18192
rect 31370 18158 31436 18192
rect 31470 18158 31536 18192
rect 31570 18158 31636 18192
rect 31670 18158 31736 18192
rect 31770 18158 31836 18192
rect 31870 18158 32676 18192
rect 32710 18158 32776 18192
rect 32810 18158 32876 18192
rect 32910 18158 32976 18192
rect 33010 18158 33076 18192
rect 33110 18158 33176 18192
rect 33210 18158 34016 18192
rect 34050 18158 34116 18192
rect 34150 18158 34216 18192
rect 34250 18158 34316 18192
rect 34350 18158 34416 18192
rect 34450 18158 34516 18192
rect 34550 18158 35356 18192
rect 35390 18158 35456 18192
rect 35490 18158 35556 18192
rect 35590 18158 35656 18192
rect 35690 18158 35756 18192
rect 35790 18158 35856 18192
rect 35890 18158 36696 18192
rect 36730 18158 36796 18192
rect 36830 18158 36896 18192
rect 36930 18158 36996 18192
rect 37030 18158 37096 18192
rect 37130 18158 37196 18192
rect 37230 18158 38036 18192
rect 38070 18158 38136 18192
rect 38170 18158 38236 18192
rect 38270 18158 38336 18192
rect 38370 18158 38436 18192
rect 38470 18158 38536 18192
rect 38570 18158 38616 18192
rect 28624 18092 38616 18158
rect 28624 18058 28656 18092
rect 28690 18058 28756 18092
rect 28790 18058 28856 18092
rect 28890 18058 28956 18092
rect 28990 18058 29056 18092
rect 29090 18058 29156 18092
rect 29190 18058 29996 18092
rect 30030 18058 30096 18092
rect 30130 18058 30196 18092
rect 30230 18058 30296 18092
rect 30330 18058 30396 18092
rect 30430 18058 30496 18092
rect 30530 18058 31336 18092
rect 31370 18058 31436 18092
rect 31470 18058 31536 18092
rect 31570 18058 31636 18092
rect 31670 18058 31736 18092
rect 31770 18058 31836 18092
rect 31870 18058 32676 18092
rect 32710 18058 32776 18092
rect 32810 18058 32876 18092
rect 32910 18058 32976 18092
rect 33010 18058 33076 18092
rect 33110 18058 33176 18092
rect 33210 18058 34016 18092
rect 34050 18058 34116 18092
rect 34150 18058 34216 18092
rect 34250 18058 34316 18092
rect 34350 18058 34416 18092
rect 34450 18058 34516 18092
rect 34550 18058 35356 18092
rect 35390 18058 35456 18092
rect 35490 18058 35556 18092
rect 35590 18058 35656 18092
rect 35690 18058 35756 18092
rect 35790 18058 35856 18092
rect 35890 18058 36696 18092
rect 36730 18058 36796 18092
rect 36830 18058 36896 18092
rect 36930 18058 36996 18092
rect 37030 18058 37096 18092
rect 37130 18058 37196 18092
rect 37230 18058 38036 18092
rect 38070 18058 38136 18092
rect 38170 18058 38236 18092
rect 38270 18058 38336 18092
rect 38370 18058 38436 18092
rect 38470 18058 38536 18092
rect 38570 18058 38616 18092
rect 39267 18083 39275 18621
rect 39669 18083 39677 18621
rect 39267 18071 39677 18083
rect 41275 18621 41685 18633
rect 41275 18083 41282 18621
rect 41676 18083 41685 18621
rect 41275 18071 41685 18083
rect 28624 17992 38616 18058
rect 28624 17958 28656 17992
rect 28690 17958 28756 17992
rect 28790 17958 28856 17992
rect 28890 17958 28956 17992
rect 28990 17958 29056 17992
rect 29090 17958 29156 17992
rect 29190 17958 29996 17992
rect 30030 17958 30096 17992
rect 30130 17958 30196 17992
rect 30230 17958 30296 17992
rect 30330 17958 30396 17992
rect 30430 17958 30496 17992
rect 30530 17958 31336 17992
rect 31370 17958 31436 17992
rect 31470 17958 31536 17992
rect 31570 17958 31636 17992
rect 31670 17958 31736 17992
rect 31770 17958 31836 17992
rect 31870 17958 32676 17992
rect 32710 17958 32776 17992
rect 32810 17958 32876 17992
rect 32910 17958 32976 17992
rect 33010 17958 33076 17992
rect 33110 17958 33176 17992
rect 33210 17958 34016 17992
rect 34050 17958 34116 17992
rect 34150 17958 34216 17992
rect 34250 17958 34316 17992
rect 34350 17958 34416 17992
rect 34450 17958 34516 17992
rect 34550 17958 35356 17992
rect 35390 17958 35456 17992
rect 35490 17958 35556 17992
rect 35590 17958 35656 17992
rect 35690 17958 35756 17992
rect 35790 17958 35856 17992
rect 35890 17958 36696 17992
rect 36730 17958 36796 17992
rect 36830 17958 36896 17992
rect 36930 17958 36996 17992
rect 37030 17958 37096 17992
rect 37130 17958 37196 17992
rect 37230 17958 38036 17992
rect 38070 17958 38136 17992
rect 38170 17958 38236 17992
rect 38270 17958 38336 17992
rect 38370 17958 38436 17992
rect 38470 17958 38536 17992
rect 38570 17958 38616 17992
rect 28624 17892 38616 17958
rect 28624 17858 28656 17892
rect 28690 17858 28756 17892
rect 28790 17858 28856 17892
rect 28890 17858 28956 17892
rect 28990 17858 29056 17892
rect 29090 17858 29156 17892
rect 29190 17858 29996 17892
rect 30030 17858 30096 17892
rect 30130 17858 30196 17892
rect 30230 17858 30296 17892
rect 30330 17858 30396 17892
rect 30430 17858 30496 17892
rect 30530 17858 31336 17892
rect 31370 17858 31436 17892
rect 31470 17858 31536 17892
rect 31570 17858 31636 17892
rect 31670 17858 31736 17892
rect 31770 17858 31836 17892
rect 31870 17858 32676 17892
rect 32710 17858 32776 17892
rect 32810 17858 32876 17892
rect 32910 17858 32976 17892
rect 33010 17858 33076 17892
rect 33110 17858 33176 17892
rect 33210 17858 34016 17892
rect 34050 17858 34116 17892
rect 34150 17858 34216 17892
rect 34250 17858 34316 17892
rect 34350 17858 34416 17892
rect 34450 17858 34516 17892
rect 34550 17858 35356 17892
rect 35390 17858 35456 17892
rect 35490 17858 35556 17892
rect 35590 17858 35656 17892
rect 35690 17858 35756 17892
rect 35790 17858 35856 17892
rect 35890 17858 36696 17892
rect 36730 17858 36796 17892
rect 36830 17858 36896 17892
rect 36930 17858 36996 17892
rect 37030 17858 37096 17892
rect 37130 17858 37196 17892
rect 37230 17858 38036 17892
rect 38070 17858 38136 17892
rect 38170 17858 38236 17892
rect 38270 17858 38336 17892
rect 38370 17858 38436 17892
rect 38470 17858 38536 17892
rect 38570 17858 38616 17892
rect 28624 17792 38616 17858
rect 28624 17758 28656 17792
rect 28690 17758 28756 17792
rect 28790 17758 28856 17792
rect 28890 17758 28956 17792
rect 28990 17758 29056 17792
rect 29090 17758 29156 17792
rect 29190 17758 29996 17792
rect 30030 17758 30096 17792
rect 30130 17758 30196 17792
rect 30230 17758 30296 17792
rect 30330 17758 30396 17792
rect 30430 17758 30496 17792
rect 30530 17758 31336 17792
rect 31370 17758 31436 17792
rect 31470 17758 31536 17792
rect 31570 17758 31636 17792
rect 31670 17758 31736 17792
rect 31770 17758 31836 17792
rect 31870 17758 32676 17792
rect 32710 17758 32776 17792
rect 32810 17758 32876 17792
rect 32910 17758 32976 17792
rect 33010 17758 33076 17792
rect 33110 17758 33176 17792
rect 33210 17758 34016 17792
rect 34050 17758 34116 17792
rect 34150 17758 34216 17792
rect 34250 17758 34316 17792
rect 34350 17758 34416 17792
rect 34450 17758 34516 17792
rect 34550 17758 35356 17792
rect 35390 17758 35456 17792
rect 35490 17758 35556 17792
rect 35590 17758 35656 17792
rect 35690 17758 35756 17792
rect 35790 17758 35856 17792
rect 35890 17758 36696 17792
rect 36730 17758 36796 17792
rect 36830 17758 36896 17792
rect 36930 17758 36996 17792
rect 37030 17758 37096 17792
rect 37130 17758 37196 17792
rect 37230 17758 38036 17792
rect 38070 17758 38136 17792
rect 38170 17758 38236 17792
rect 38270 17758 38336 17792
rect 38370 17758 38436 17792
rect 38470 17758 38536 17792
rect 38570 17758 38616 17792
rect 28624 17692 38616 17758
rect 28624 17658 28656 17692
rect 28690 17672 28756 17692
rect 28690 17658 28724 17672
rect 28790 17658 28856 17692
rect 28890 17658 28956 17692
rect 28990 17658 29056 17692
rect 29090 17658 29156 17692
rect 29190 17658 29996 17692
rect 30030 17658 30096 17692
rect 30130 17658 30196 17692
rect 30230 17658 30296 17692
rect 30330 17658 30396 17692
rect 30430 17658 30496 17692
rect 30530 17658 31336 17692
rect 31370 17658 31436 17692
rect 31470 17658 31536 17692
rect 31570 17658 31636 17692
rect 31670 17658 31736 17692
rect 31770 17658 31836 17692
rect 31870 17658 32676 17692
rect 32710 17658 32776 17692
rect 32810 17658 32876 17692
rect 32910 17658 32976 17692
rect 33010 17658 33076 17692
rect 33110 17658 33176 17692
rect 33210 17658 34016 17692
rect 34050 17658 34116 17692
rect 34150 17658 34216 17692
rect 34250 17658 34316 17692
rect 34350 17658 34416 17692
rect 34450 17658 34516 17692
rect 34550 17658 35356 17692
rect 35390 17658 35456 17692
rect 35490 17658 35556 17692
rect 35590 17658 35656 17692
rect 35690 17658 35756 17692
rect 35790 17658 35856 17692
rect 35890 17658 36696 17692
rect 36730 17658 36796 17692
rect 36830 17658 36896 17692
rect 36930 17658 36996 17692
rect 37030 17658 37096 17692
rect 37130 17658 37196 17692
rect 37230 17658 38036 17692
rect 38070 17658 38136 17692
rect 38170 17658 38236 17692
rect 38270 17658 38336 17692
rect 38370 17658 38436 17692
rect 38470 17658 38536 17692
rect 38570 17658 38616 17692
rect 28624 17626 28724 17658
rect 28718 17620 28724 17626
rect 28776 17626 38616 17658
rect 39267 17661 39677 17673
rect 28776 17620 28782 17626
rect 26737 17579 26743 17613
rect 26777 17579 26783 17613
rect 26737 17541 26783 17579
rect 26737 17507 26743 17541
rect 26777 17507 26783 17541
rect 26737 17469 26783 17507
rect 26737 17435 26743 17469
rect 26777 17435 26783 17469
rect 26737 17397 26783 17435
rect 26737 17363 26743 17397
rect 26777 17363 26783 17397
rect 26737 17347 26783 17363
rect 23382 17280 23388 17332
rect 23440 17280 23446 17332
rect 23400 17252 23428 17280
rect 23937 17255 23995 17261
rect 23937 17252 23949 17255
rect 23400 17224 23949 17252
rect 23937 17221 23949 17224
rect 23983 17221 23995 17255
rect 23937 17215 23995 17221
rect 26510 17144 26516 17196
rect 26568 17144 26574 17196
rect 15392 17107 15824 17123
rect 26513 17119 26525 17144
rect 26559 17119 26571 17144
rect 26513 17113 26571 17119
rect 39267 17123 39275 17661
rect 39669 17123 39677 17661
rect 39267 17111 39677 17123
rect 41264 17661 41696 18071
rect 41264 17123 41282 17661
rect 41676 17123 41696 17661
rect 41264 17107 41696 17123
rect 900 17050 47736 17052
rect 900 16934 922 17050
rect 2510 17009 46126 17050
rect 2510 16975 6197 17009
rect 6231 16975 6597 17009
rect 6631 16975 6997 17009
rect 7031 16975 7397 17009
rect 7431 16975 7797 17009
rect 7831 16975 8197 17009
rect 8231 16975 8597 17009
rect 8631 16975 8997 17009
rect 9031 16975 9397 17009
rect 9431 16975 9797 17009
rect 9831 16975 10823 17009
rect 10857 16975 11023 17009
rect 11057 16975 11223 17009
rect 11257 16975 11423 17009
rect 11457 16975 11623 17009
rect 11657 16975 11823 17009
rect 11857 16975 12023 17009
rect 12057 16975 12223 17009
rect 12257 16975 12423 17009
rect 12457 16975 12623 17009
rect 12657 16975 12823 17009
rect 12857 16975 13567 17009
rect 13601 16975 13767 17009
rect 13801 16975 13967 17009
rect 14001 16975 14167 17009
rect 14201 16975 14367 17009
rect 14401 16975 14567 17009
rect 14601 16975 14767 17009
rect 14801 16975 14967 17009
rect 15001 16975 15167 17009
rect 15201 16975 15367 17009
rect 15401 16975 15567 17009
rect 15601 16975 16293 17009
rect 16327 16975 16693 17009
rect 16727 16975 17093 17009
rect 17127 16992 17493 17009
rect 17127 16975 17408 16992
rect 2510 16940 17408 16975
rect 17460 16975 17493 16992
rect 17527 16975 17893 17009
rect 17927 16975 18293 17009
rect 18327 16975 18693 17009
rect 18727 16975 19093 17009
rect 19127 16975 19493 17009
rect 19527 16975 19893 17009
rect 19927 16975 20293 17009
rect 20327 16975 20693 17009
rect 20727 16975 21093 17009
rect 21127 16975 21493 17009
rect 21527 16975 21893 17009
rect 21927 16975 22293 17009
rect 22327 16975 22693 17009
rect 22727 16975 23093 17009
rect 23127 16975 24131 17009
rect 24165 16975 24531 17009
rect 24565 16975 24931 17009
rect 24965 16975 25331 17009
rect 25365 16975 25731 17009
rect 25765 16975 26131 17009
rect 26165 16975 26531 17009
rect 26565 16975 28443 17009
rect 28477 16992 28643 17009
rect 28677 16992 28843 17009
rect 28477 16975 28632 16992
rect 28684 16975 28843 16992
rect 28877 16975 29043 17009
rect 29077 16975 29243 17009
rect 29277 16975 29443 17009
rect 29477 16975 29643 17009
rect 29677 16975 29843 17009
rect 29877 16975 30043 17009
rect 30077 16975 30243 17009
rect 30277 16975 30443 17009
rect 30477 16975 30643 17009
rect 30677 16975 30843 17009
rect 30877 16975 31043 17009
rect 31077 16975 31243 17009
rect 31277 16975 31443 17009
rect 31477 16975 31643 17009
rect 31677 16975 31843 17009
rect 31877 16975 32043 17009
rect 32077 16975 32243 17009
rect 32277 16975 32443 17009
rect 32477 16975 32643 17009
rect 32677 16975 32843 17009
rect 32877 16975 33043 17009
rect 33077 16975 33243 17009
rect 33277 16975 33443 17009
rect 33477 16975 33643 17009
rect 33677 16975 33843 17009
rect 33877 16975 34043 17009
rect 34077 16975 34243 17009
rect 34277 16975 34443 17009
rect 34477 16975 34643 17009
rect 34677 16975 34843 17009
rect 34877 16975 35043 17009
rect 35077 16975 35243 17009
rect 35277 16975 35443 17009
rect 35477 16975 35643 17009
rect 35677 16975 35843 17009
rect 35877 16975 36043 17009
rect 36077 16975 36243 17009
rect 36277 16975 36443 17009
rect 36477 16975 36643 17009
rect 36677 16975 36843 17009
rect 36877 16975 37043 17009
rect 37077 16975 37243 17009
rect 37277 16975 37443 17009
rect 37477 16975 37643 17009
rect 37677 16975 37843 17009
rect 37877 16975 38043 17009
rect 38077 16975 38243 17009
rect 38277 16975 38443 17009
rect 38477 16975 38643 17009
rect 38677 16975 38843 17009
rect 38877 16975 39439 17009
rect 39473 16975 39639 17009
rect 39673 16975 39839 17009
rect 39873 16975 40039 17009
rect 40073 16975 40239 17009
rect 40273 16975 40439 17009
rect 40473 16975 40639 17009
rect 40673 16975 40839 17009
rect 40873 16975 41039 17009
rect 41073 16975 41239 17009
rect 41273 16975 41439 17009
rect 41473 16975 46126 17009
rect 17460 16940 28632 16975
rect 28684 16940 46126 16975
rect 2510 16934 46126 16940
rect 47714 16934 47736 17050
rect 900 16932 47736 16934
rect 27614 15444 27620 15496
rect 27672 15444 27678 15496
rect 8110 15376 8116 15428
rect 8168 15416 8174 15428
rect 27632 15416 27660 15444
rect 8168 15388 27660 15416
rect 8168 15376 8174 15388
rect 3348 15170 45288 15172
rect 3348 15054 3370 15170
rect 4958 15129 43678 15170
rect 4958 15095 8079 15129
rect 8113 15095 8279 15129
rect 8313 15095 8479 15129
rect 8513 15095 8679 15129
rect 8713 15095 8879 15129
rect 8913 15095 9079 15129
rect 9113 15095 9279 15129
rect 9313 15095 9479 15129
rect 9513 15095 9679 15129
rect 9713 15095 9879 15129
rect 9913 15095 10079 15129
rect 10113 15095 10823 15129
rect 10857 15095 11023 15129
rect 11057 15095 11223 15129
rect 11257 15095 11423 15129
rect 11457 15095 11623 15129
rect 11657 15095 11823 15129
rect 11857 15095 12023 15129
rect 12057 15095 12223 15129
rect 12257 15095 12423 15129
rect 12457 15095 12623 15129
rect 12657 15095 12823 15129
rect 12857 15095 13567 15129
rect 13601 15095 13767 15129
rect 13801 15095 13967 15129
rect 14001 15095 14167 15129
rect 14201 15095 14367 15129
rect 14401 15095 14567 15129
rect 14601 15095 14767 15129
rect 14801 15095 14967 15129
rect 15001 15095 15167 15129
rect 15201 15095 15367 15129
rect 15401 15095 15567 15129
rect 15601 15095 16293 15129
rect 16327 15095 16693 15129
rect 16727 15095 17093 15129
rect 17127 15095 17493 15129
rect 17527 15095 17893 15129
rect 17927 15095 18293 15129
rect 18327 15095 18693 15129
rect 18727 15095 19093 15129
rect 19127 15095 19493 15129
rect 19527 15095 19893 15129
rect 19927 15095 20293 15129
rect 20327 15095 20693 15129
rect 20727 15095 21093 15129
rect 21127 15095 21493 15129
rect 21527 15095 21893 15129
rect 21927 15095 22293 15129
rect 22327 15095 22693 15129
rect 22727 15095 23093 15129
rect 23127 15095 23759 15129
rect 23793 15095 23959 15129
rect 23993 15095 24159 15129
rect 24193 15095 24359 15129
rect 24393 15095 24559 15129
rect 24593 15095 24759 15129
rect 24793 15095 24959 15129
rect 24993 15095 25159 15129
rect 25193 15095 25359 15129
rect 25393 15095 25559 15129
rect 25593 15095 25759 15129
rect 25793 15095 28443 15129
rect 28477 15095 28643 15129
rect 28677 15095 28843 15129
rect 28877 15095 29043 15129
rect 29077 15095 29243 15129
rect 29277 15095 29443 15129
rect 29477 15095 29643 15129
rect 29677 15095 29843 15129
rect 29877 15095 30043 15129
rect 30077 15095 30243 15129
rect 30277 15095 30443 15129
rect 30477 15095 30643 15129
rect 30677 15095 30843 15129
rect 30877 15095 31043 15129
rect 31077 15095 31243 15129
rect 31277 15095 31443 15129
rect 31477 15095 31643 15129
rect 31677 15095 31843 15129
rect 31877 15095 32043 15129
rect 32077 15095 32243 15129
rect 32277 15095 32443 15129
rect 32477 15095 32643 15129
rect 32677 15095 32843 15129
rect 32877 15095 33043 15129
rect 33077 15095 33243 15129
rect 33277 15095 33443 15129
rect 33477 15095 33643 15129
rect 33677 15095 33843 15129
rect 33877 15095 34043 15129
rect 34077 15095 34243 15129
rect 34277 15095 34443 15129
rect 34477 15095 34643 15129
rect 34677 15095 34843 15129
rect 34877 15095 35043 15129
rect 35077 15095 35243 15129
rect 35277 15095 35443 15129
rect 35477 15095 35643 15129
rect 35677 15095 35843 15129
rect 35877 15095 36043 15129
rect 36077 15095 36243 15129
rect 36277 15095 36443 15129
rect 36477 15095 36643 15129
rect 36677 15095 36843 15129
rect 36877 15095 37043 15129
rect 37077 15095 37243 15129
rect 37277 15095 37443 15129
rect 37477 15095 37643 15129
rect 37677 15095 37843 15129
rect 37877 15095 38043 15129
rect 38077 15095 38243 15129
rect 38277 15095 38443 15129
rect 38477 15095 38643 15129
rect 38677 15095 38843 15129
rect 38877 15095 39439 15129
rect 39473 15095 39639 15129
rect 39673 15095 39839 15129
rect 39873 15095 40039 15129
rect 40073 15095 40239 15129
rect 40273 15095 40439 15129
rect 40473 15095 40639 15129
rect 40673 15095 40839 15129
rect 40873 15095 41039 15129
rect 41073 15095 41239 15129
rect 41273 15095 41439 15129
rect 41473 15095 43678 15129
rect 4958 15054 43678 15095
rect 45266 15054 45288 15170
rect 3348 15052 45288 15054
rect 7907 14872 8317 14873
rect 8754 14872 8760 14884
rect 7907 14861 8760 14872
rect 7907 14323 7915 14861
rect 8309 14844 8760 14861
rect 8309 14323 8317 14844
rect 8754 14832 8760 14844
rect 8812 14832 8818 14884
rect 39298 14873 39304 14884
rect 9915 14861 10325 14873
rect 7907 14311 8317 14323
rect 9915 14323 9922 14861
rect 10316 14323 10325 14861
rect 10651 14861 11061 14873
rect 10410 14356 10416 14408
rect 10468 14396 10474 14408
rect 10651 14396 10659 14861
rect 10468 14368 10659 14396
rect 10468 14356 10474 14368
rect 9915 14311 10325 14323
rect 10651 14323 10659 14368
rect 11053 14323 11061 14861
rect 10651 14311 11061 14323
rect 12659 14861 13069 14873
rect 12659 14323 12666 14861
rect 13060 14323 13069 14861
rect 12659 14311 13069 14323
rect 13395 14861 13805 14873
rect 13395 14323 13403 14861
rect 13797 14396 13805 14861
rect 15403 14861 15813 14873
rect 14734 14396 14740 14408
rect 13797 14368 14740 14396
rect 13797 14323 13805 14368
rect 14734 14356 14740 14368
rect 14792 14356 14798 14408
rect 13395 14311 13805 14323
rect 15403 14323 15410 14861
rect 15804 14323 15813 14861
rect 23587 14861 23997 14873
rect 23587 14340 23595 14861
rect 15403 14311 15813 14323
rect 7907 13901 8317 13913
rect 7907 13363 7915 13901
rect 8309 13363 8317 13901
rect 7907 13351 7932 13363
rect 7926 13336 7932 13351
rect 7984 13351 8317 13363
rect 9904 13901 10336 14311
rect 9904 13363 9922 13901
rect 10316 13363 10336 13901
rect 7984 13336 7990 13351
rect 9904 13347 10336 13363
rect 10651 13901 11061 13913
rect 10651 13363 10659 13901
rect 11053 13363 11061 13901
rect 10651 13351 10692 13363
rect 10686 13336 10692 13351
rect 10744 13351 11061 13363
rect 12648 13901 13080 14311
rect 12648 13363 12666 13901
rect 13060 13363 13080 13901
rect 10744 13336 10750 13351
rect 12648 13347 13080 13363
rect 13395 13901 13805 13913
rect 13395 13363 13403 13901
rect 13797 13363 13805 13901
rect 13395 13351 13728 13363
rect 13722 13336 13728 13351
rect 13780 13351 13805 13363
rect 15392 13901 15824 14311
rect 23566 14288 23572 14340
rect 23989 14323 23997 14861
rect 23624 14311 23997 14323
rect 25595 14861 26005 14873
rect 25595 14323 25602 14861
rect 25996 14323 26005 14861
rect 39267 14861 39304 14873
rect 39356 14873 39362 14884
rect 39356 14861 39677 14873
rect 28286 14796 38954 14802
rect 28286 14762 28306 14796
rect 28340 14762 28396 14796
rect 28430 14762 28486 14796
rect 28520 14762 28576 14796
rect 28610 14762 28666 14796
rect 28700 14762 28756 14796
rect 28790 14762 28846 14796
rect 28880 14762 28936 14796
rect 28970 14762 29026 14796
rect 29060 14762 29116 14796
rect 29150 14762 29206 14796
rect 29240 14762 29296 14796
rect 29330 14762 29386 14796
rect 29420 14762 29476 14796
rect 29510 14762 29646 14796
rect 29680 14762 29736 14796
rect 29770 14762 29826 14796
rect 29860 14762 29916 14796
rect 29950 14762 30006 14796
rect 30040 14762 30096 14796
rect 30130 14762 30186 14796
rect 30220 14762 30276 14796
rect 30310 14762 30366 14796
rect 30400 14762 30456 14796
rect 30490 14762 30546 14796
rect 30580 14762 30636 14796
rect 30670 14762 30726 14796
rect 30760 14762 30816 14796
rect 30850 14762 30986 14796
rect 31020 14762 31076 14796
rect 31110 14762 31166 14796
rect 31200 14762 31256 14796
rect 31290 14762 31346 14796
rect 31380 14762 31436 14796
rect 31470 14762 31526 14796
rect 31560 14762 31616 14796
rect 31650 14762 31706 14796
rect 31740 14762 31796 14796
rect 31830 14762 31886 14796
rect 31920 14762 31976 14796
rect 32010 14762 32066 14796
rect 32100 14762 32156 14796
rect 32190 14762 32326 14796
rect 32360 14762 32416 14796
rect 32450 14762 32506 14796
rect 32540 14762 32596 14796
rect 32630 14762 32686 14796
rect 32720 14762 32776 14796
rect 32810 14762 32866 14796
rect 32900 14762 32956 14796
rect 32990 14762 33046 14796
rect 33080 14762 33136 14796
rect 33170 14762 33226 14796
rect 33260 14762 33316 14796
rect 33350 14762 33406 14796
rect 33440 14762 33496 14796
rect 33530 14762 33666 14796
rect 33700 14762 33756 14796
rect 33790 14762 33846 14796
rect 33880 14762 33936 14796
rect 33970 14762 34026 14796
rect 34060 14762 34116 14796
rect 34150 14762 34206 14796
rect 34240 14762 34296 14796
rect 34330 14762 34386 14796
rect 34420 14762 34476 14796
rect 34510 14762 34566 14796
rect 34600 14762 34656 14796
rect 34690 14762 34746 14796
rect 34780 14762 34836 14796
rect 34870 14762 35006 14796
rect 35040 14762 35096 14796
rect 35130 14762 35186 14796
rect 35220 14762 35276 14796
rect 35310 14762 35366 14796
rect 35400 14762 35456 14796
rect 35490 14762 35546 14796
rect 35580 14762 35636 14796
rect 35670 14762 35726 14796
rect 35760 14762 35816 14796
rect 35850 14762 35906 14796
rect 35940 14762 35996 14796
rect 36030 14762 36086 14796
rect 36120 14762 36176 14796
rect 36210 14762 36346 14796
rect 36380 14762 36436 14796
rect 36470 14762 36526 14796
rect 36560 14762 36616 14796
rect 36650 14762 36706 14796
rect 36740 14762 36796 14796
rect 36830 14762 36886 14796
rect 36920 14762 36976 14796
rect 37010 14762 37066 14796
rect 37100 14762 37156 14796
rect 37190 14762 37246 14796
rect 37280 14762 37336 14796
rect 37370 14762 37426 14796
rect 37460 14762 37516 14796
rect 37550 14762 37686 14796
rect 37720 14762 37776 14796
rect 37810 14762 37866 14796
rect 37900 14762 37956 14796
rect 37990 14762 38046 14796
rect 38080 14762 38136 14796
rect 38170 14762 38226 14796
rect 38260 14762 38316 14796
rect 38350 14762 38406 14796
rect 38440 14762 38496 14796
rect 38530 14762 38586 14796
rect 38620 14762 38676 14796
rect 38710 14762 38766 14796
rect 38800 14762 38856 14796
rect 38890 14762 38954 14796
rect 28286 14732 38954 14762
rect 28644 14652 28672 14732
rect 28450 14636 38790 14652
rect 28450 14602 28470 14636
rect 28504 14602 28560 14636
rect 28594 14612 28650 14636
rect 28594 14602 28632 14612
rect 28684 14602 28740 14636
rect 28774 14602 28830 14636
rect 28864 14602 28920 14636
rect 28954 14602 29010 14636
rect 29044 14602 29100 14636
rect 29134 14602 29190 14636
rect 29224 14602 29280 14636
rect 29314 14602 29370 14636
rect 29404 14602 29810 14636
rect 29844 14602 29900 14636
rect 29934 14602 29990 14636
rect 30024 14602 30080 14636
rect 30114 14602 30170 14636
rect 30204 14602 30260 14636
rect 30294 14602 30350 14636
rect 30384 14602 30440 14636
rect 30474 14602 30530 14636
rect 30564 14602 30620 14636
rect 30654 14602 30710 14636
rect 30744 14602 31150 14636
rect 31184 14602 31240 14636
rect 31274 14602 31330 14636
rect 31364 14602 31420 14636
rect 31454 14602 31510 14636
rect 31544 14602 31600 14636
rect 31634 14602 31690 14636
rect 31724 14602 31780 14636
rect 31814 14602 31870 14636
rect 31904 14602 31960 14636
rect 31994 14602 32050 14636
rect 32084 14602 32490 14636
rect 32524 14602 32580 14636
rect 32614 14602 32670 14636
rect 32704 14602 32760 14636
rect 32794 14602 32850 14636
rect 32884 14602 32940 14636
rect 32974 14602 33030 14636
rect 33064 14602 33120 14636
rect 33154 14602 33210 14636
rect 33244 14602 33300 14636
rect 33334 14602 33390 14636
rect 33424 14602 33830 14636
rect 33864 14602 33920 14636
rect 33954 14602 34010 14636
rect 34044 14602 34100 14636
rect 34134 14602 34190 14636
rect 34224 14602 34280 14636
rect 34314 14602 34370 14636
rect 34404 14602 34460 14636
rect 34494 14602 34550 14636
rect 34584 14602 34640 14636
rect 34674 14602 34730 14636
rect 34764 14602 35170 14636
rect 35204 14602 35260 14636
rect 35294 14602 35350 14636
rect 35384 14602 35440 14636
rect 35474 14602 35530 14636
rect 35564 14602 35620 14636
rect 35654 14602 35710 14636
rect 35744 14602 35800 14636
rect 35834 14602 35890 14636
rect 35924 14602 35980 14636
rect 36014 14602 36070 14636
rect 36104 14602 36510 14636
rect 36544 14602 36600 14636
rect 36634 14602 36690 14636
rect 36724 14602 36780 14636
rect 36814 14602 36870 14636
rect 36904 14602 36960 14636
rect 36994 14602 37050 14636
rect 37084 14602 37140 14636
rect 37174 14602 37230 14636
rect 37264 14602 37320 14636
rect 37354 14602 37410 14636
rect 37444 14602 37850 14636
rect 37884 14602 37940 14636
rect 37974 14602 38030 14636
rect 38064 14602 38120 14636
rect 38154 14602 38210 14636
rect 38244 14602 38300 14636
rect 38334 14602 38390 14636
rect 38424 14602 38480 14636
rect 38514 14602 38570 14636
rect 38604 14602 38660 14636
rect 38694 14602 38750 14636
rect 38784 14602 38790 14636
rect 28450 14582 28632 14602
rect 28626 14560 28632 14582
rect 28684 14582 38790 14602
rect 28684 14560 28690 14582
rect 25595 14311 26005 14323
rect 28624 14476 38616 14478
rect 28624 14432 28724 14476
rect 28776 14432 38616 14476
rect 28624 14398 28656 14432
rect 28690 14424 28724 14432
rect 28690 14398 28756 14424
rect 28790 14398 28856 14432
rect 28890 14398 28956 14432
rect 28990 14398 29056 14432
rect 29090 14398 29156 14432
rect 29190 14398 29996 14432
rect 30030 14398 30096 14432
rect 30130 14398 30196 14432
rect 30230 14398 30296 14432
rect 30330 14398 30396 14432
rect 30430 14398 30496 14432
rect 30530 14398 31336 14432
rect 31370 14398 31436 14432
rect 31470 14398 31536 14432
rect 31570 14398 31636 14432
rect 31670 14398 31736 14432
rect 31770 14398 31836 14432
rect 31870 14398 32676 14432
rect 32710 14398 32776 14432
rect 32810 14398 32876 14432
rect 32910 14398 32976 14432
rect 33010 14398 33076 14432
rect 33110 14398 33176 14432
rect 33210 14398 34016 14432
rect 34050 14398 34116 14432
rect 34150 14398 34216 14432
rect 34250 14398 34316 14432
rect 34350 14398 34416 14432
rect 34450 14398 34516 14432
rect 34550 14398 35356 14432
rect 35390 14398 35456 14432
rect 35490 14398 35556 14432
rect 35590 14398 35656 14432
rect 35690 14398 35756 14432
rect 35790 14398 35856 14432
rect 35890 14398 36696 14432
rect 36730 14398 36796 14432
rect 36830 14398 36896 14432
rect 36930 14398 36996 14432
rect 37030 14398 37096 14432
rect 37130 14398 37196 14432
rect 37230 14398 38036 14432
rect 38070 14398 38136 14432
rect 38170 14398 38236 14432
rect 38270 14398 38336 14432
rect 38370 14398 38436 14432
rect 38470 14398 38536 14432
rect 38570 14398 38616 14432
rect 28624 14332 38616 14398
rect 23624 14288 23630 14311
rect 15392 13363 15410 13901
rect 15804 13363 15824 13901
rect 23587 13901 23997 13913
rect 20070 13404 20076 13456
rect 20128 13444 20134 13456
rect 23587 13444 23595 13901
rect 20128 13416 23595 13444
rect 20128 13404 20134 13416
rect 13780 13336 13786 13351
rect 15392 13347 15824 13363
rect 23587 13363 23595 13416
rect 23989 13363 23997 13901
rect 23587 13351 23997 13363
rect 25584 13901 26016 14311
rect 25584 13363 25602 13901
rect 25996 13363 26016 13901
rect 28624 14298 28656 14332
rect 28690 14298 28756 14332
rect 28790 14298 28856 14332
rect 28890 14298 28956 14332
rect 28990 14298 29056 14332
rect 29090 14298 29156 14332
rect 29190 14298 29996 14332
rect 30030 14298 30096 14332
rect 30130 14298 30196 14332
rect 30230 14298 30296 14332
rect 30330 14298 30396 14332
rect 30430 14298 30496 14332
rect 30530 14298 31336 14332
rect 31370 14298 31436 14332
rect 31470 14298 31536 14332
rect 31570 14298 31636 14332
rect 31670 14298 31736 14332
rect 31770 14298 31836 14332
rect 31870 14298 32676 14332
rect 32710 14298 32776 14332
rect 32810 14298 32876 14332
rect 32910 14298 32976 14332
rect 33010 14298 33076 14332
rect 33110 14298 33176 14332
rect 33210 14298 34016 14332
rect 34050 14298 34116 14332
rect 34150 14298 34216 14332
rect 34250 14298 34316 14332
rect 34350 14298 34416 14332
rect 34450 14298 34516 14332
rect 34550 14298 35356 14332
rect 35390 14298 35456 14332
rect 35490 14298 35556 14332
rect 35590 14298 35656 14332
rect 35690 14298 35756 14332
rect 35790 14298 35856 14332
rect 35890 14298 36696 14332
rect 36730 14298 36796 14332
rect 36830 14298 36896 14332
rect 36930 14298 36996 14332
rect 37030 14298 37096 14332
rect 37130 14298 37196 14332
rect 37230 14298 38036 14332
rect 38070 14298 38136 14332
rect 38170 14298 38236 14332
rect 38270 14298 38336 14332
rect 38370 14298 38436 14332
rect 38470 14298 38536 14332
rect 38570 14298 38616 14332
rect 39267 14323 39275 14861
rect 39669 14323 39677 14861
rect 39267 14311 39677 14323
rect 41275 14861 41685 14873
rect 41275 14323 41282 14861
rect 41676 14323 41685 14861
rect 41275 14311 41685 14323
rect 28624 14232 38616 14298
rect 28624 14198 28656 14232
rect 28690 14198 28756 14232
rect 28790 14198 28856 14232
rect 28890 14198 28956 14232
rect 28990 14198 29056 14232
rect 29090 14198 29156 14232
rect 29190 14198 29996 14232
rect 30030 14198 30096 14232
rect 30130 14198 30196 14232
rect 30230 14198 30296 14232
rect 30330 14198 30396 14232
rect 30430 14198 30496 14232
rect 30530 14198 31336 14232
rect 31370 14198 31436 14232
rect 31470 14198 31536 14232
rect 31570 14198 31636 14232
rect 31670 14198 31736 14232
rect 31770 14198 31836 14232
rect 31870 14198 32676 14232
rect 32710 14198 32776 14232
rect 32810 14198 32876 14232
rect 32910 14198 32976 14232
rect 33010 14198 33076 14232
rect 33110 14198 33176 14232
rect 33210 14198 34016 14232
rect 34050 14198 34116 14232
rect 34150 14198 34216 14232
rect 34250 14198 34316 14232
rect 34350 14198 34416 14232
rect 34450 14198 34516 14232
rect 34550 14198 35356 14232
rect 35390 14198 35456 14232
rect 35490 14198 35556 14232
rect 35590 14198 35656 14232
rect 35690 14198 35756 14232
rect 35790 14198 35856 14232
rect 35890 14198 36696 14232
rect 36730 14198 36796 14232
rect 36830 14198 36896 14232
rect 36930 14198 36996 14232
rect 37030 14198 37096 14232
rect 37130 14198 37196 14232
rect 37230 14198 38036 14232
rect 38070 14198 38136 14232
rect 38170 14198 38236 14232
rect 38270 14198 38336 14232
rect 38370 14198 38436 14232
rect 38470 14198 38536 14232
rect 38570 14198 38616 14232
rect 28624 14132 38616 14198
rect 28624 14098 28656 14132
rect 28690 14098 28756 14132
rect 28790 14098 28856 14132
rect 28890 14098 28956 14132
rect 28990 14098 29056 14132
rect 29090 14098 29156 14132
rect 29190 14098 29996 14132
rect 30030 14098 30096 14132
rect 30130 14098 30196 14132
rect 30230 14098 30296 14132
rect 30330 14098 30396 14132
rect 30430 14098 30496 14132
rect 30530 14098 31336 14132
rect 31370 14098 31436 14132
rect 31470 14098 31536 14132
rect 31570 14098 31636 14132
rect 31670 14098 31736 14132
rect 31770 14098 31836 14132
rect 31870 14098 32676 14132
rect 32710 14098 32776 14132
rect 32810 14098 32876 14132
rect 32910 14098 32976 14132
rect 33010 14098 33076 14132
rect 33110 14098 33176 14132
rect 33210 14098 34016 14132
rect 34050 14098 34116 14132
rect 34150 14098 34216 14132
rect 34250 14098 34316 14132
rect 34350 14098 34416 14132
rect 34450 14098 34516 14132
rect 34550 14098 35356 14132
rect 35390 14098 35456 14132
rect 35490 14098 35556 14132
rect 35590 14098 35656 14132
rect 35690 14098 35756 14132
rect 35790 14098 35856 14132
rect 35890 14098 36696 14132
rect 36730 14098 36796 14132
rect 36830 14098 36896 14132
rect 36930 14098 36996 14132
rect 37030 14098 37096 14132
rect 37130 14098 37196 14132
rect 37230 14098 38036 14132
rect 38070 14098 38136 14132
rect 38170 14098 38236 14132
rect 38270 14098 38336 14132
rect 38370 14098 38436 14132
rect 38470 14098 38536 14132
rect 38570 14098 38616 14132
rect 28624 14032 38616 14098
rect 28624 13998 28656 14032
rect 28690 13998 28756 14032
rect 28790 13998 28856 14032
rect 28890 13998 28956 14032
rect 28990 13998 29056 14032
rect 29090 13998 29156 14032
rect 29190 13998 29996 14032
rect 30030 13998 30096 14032
rect 30130 13998 30196 14032
rect 30230 13998 30296 14032
rect 30330 13998 30396 14032
rect 30430 13998 30496 14032
rect 30530 13998 31336 14032
rect 31370 13998 31436 14032
rect 31470 13998 31536 14032
rect 31570 13998 31636 14032
rect 31670 13998 31736 14032
rect 31770 13998 31836 14032
rect 31870 13998 32676 14032
rect 32710 13998 32776 14032
rect 32810 13998 32876 14032
rect 32910 13998 32976 14032
rect 33010 13998 33076 14032
rect 33110 13998 33176 14032
rect 33210 13998 34016 14032
rect 34050 13998 34116 14032
rect 34150 13998 34216 14032
rect 34250 13998 34316 14032
rect 34350 13998 34416 14032
rect 34450 13998 34516 14032
rect 34550 13998 35356 14032
rect 35390 13998 35456 14032
rect 35490 13998 35556 14032
rect 35590 13998 35656 14032
rect 35690 13998 35756 14032
rect 35790 13998 35856 14032
rect 35890 13998 36696 14032
rect 36730 13998 36796 14032
rect 36830 13998 36896 14032
rect 36930 13998 36996 14032
rect 37030 13998 37096 14032
rect 37130 13998 37196 14032
rect 37230 13998 38036 14032
rect 38070 13998 38136 14032
rect 38170 13998 38236 14032
rect 38270 13998 38336 14032
rect 38370 13998 38436 14032
rect 38470 13998 38536 14032
rect 38570 13998 38616 14032
rect 28624 13932 38616 13998
rect 28624 13898 28656 13932
rect 28690 13898 28756 13932
rect 28790 13898 28856 13932
rect 28890 13898 28956 13932
rect 28990 13898 29056 13932
rect 29090 13898 29156 13932
rect 29190 13898 29996 13932
rect 30030 13898 30096 13932
rect 30130 13898 30196 13932
rect 30230 13898 30296 13932
rect 30330 13898 30396 13932
rect 30430 13898 30496 13932
rect 30530 13898 31336 13932
rect 31370 13898 31436 13932
rect 31470 13898 31536 13932
rect 31570 13898 31636 13932
rect 31670 13898 31736 13932
rect 31770 13898 31836 13932
rect 31870 13898 32676 13932
rect 32710 13898 32776 13932
rect 32810 13898 32876 13932
rect 32910 13898 32976 13932
rect 33010 13898 33076 13932
rect 33110 13898 33176 13932
rect 33210 13898 34016 13932
rect 34050 13898 34116 13932
rect 34150 13898 34216 13932
rect 34250 13898 34316 13932
rect 34350 13898 34416 13932
rect 34450 13898 34516 13932
rect 34550 13898 35356 13932
rect 35390 13898 35456 13932
rect 35490 13898 35556 13932
rect 35590 13898 35656 13932
rect 35690 13898 35756 13932
rect 35790 13898 35856 13932
rect 35890 13898 36696 13932
rect 36730 13898 36796 13932
rect 36830 13898 36896 13932
rect 36930 13898 36996 13932
rect 37030 13898 37096 13932
rect 37130 13898 37196 13932
rect 37230 13898 38036 13932
rect 38070 13898 38136 13932
rect 38170 13898 38236 13932
rect 38270 13898 38336 13932
rect 38370 13898 38436 13932
rect 38470 13898 38536 13932
rect 38570 13898 38616 13932
rect 28624 13866 38616 13898
rect 39267 13901 39677 13913
rect 39267 13444 39275 13901
rect 38212 13416 39275 13444
rect 38212 13388 38240 13416
rect 25584 13347 26016 13363
rect 38194 13336 38200 13388
rect 38252 13336 38258 13388
rect 39267 13363 39275 13416
rect 39669 13363 39677 13901
rect 39267 13351 39677 13363
rect 41264 13901 41696 14311
rect 41264 13363 41282 13901
rect 41676 13363 41696 13901
rect 41264 13347 41696 13363
rect 900 13290 47736 13292
rect 900 13174 922 13290
rect 2510 13252 46126 13290
rect 2510 13249 17132 13252
rect 2510 13215 8079 13249
rect 8113 13215 8279 13249
rect 8313 13215 8479 13249
rect 8513 13215 8679 13249
rect 8713 13215 8879 13249
rect 8913 13215 9079 13249
rect 9113 13215 9279 13249
rect 9313 13215 9479 13249
rect 9513 13215 9679 13249
rect 9713 13215 9879 13249
rect 9913 13215 10079 13249
rect 10113 13215 10823 13249
rect 10857 13215 11023 13249
rect 11057 13215 11223 13249
rect 11257 13215 11423 13249
rect 11457 13215 11623 13249
rect 11657 13215 11823 13249
rect 11857 13215 12023 13249
rect 12057 13215 12223 13249
rect 12257 13215 12423 13249
rect 12457 13215 12623 13249
rect 12657 13215 12823 13249
rect 12857 13215 13567 13249
rect 13601 13215 13767 13249
rect 13801 13215 13967 13249
rect 14001 13215 14167 13249
rect 14201 13215 14367 13249
rect 14401 13215 14567 13249
rect 14601 13215 14767 13249
rect 14801 13215 14967 13249
rect 15001 13215 15167 13249
rect 15201 13215 15367 13249
rect 15401 13215 15567 13249
rect 15601 13215 16293 13249
rect 16327 13215 16693 13249
rect 16727 13215 17093 13249
rect 17127 13215 17132 13249
rect 2510 13200 17132 13215
rect 17184 13249 28632 13252
rect 28684 13249 46126 13252
rect 17184 13215 17493 13249
rect 17527 13215 17893 13249
rect 17927 13215 18293 13249
rect 18327 13215 18693 13249
rect 18727 13215 19093 13249
rect 19127 13215 19493 13249
rect 19527 13215 19893 13249
rect 19927 13215 20293 13249
rect 20327 13215 20693 13249
rect 20727 13215 21093 13249
rect 21127 13215 21493 13249
rect 21527 13215 21893 13249
rect 21927 13215 22293 13249
rect 22327 13215 22693 13249
rect 22727 13215 23093 13249
rect 23127 13215 23759 13249
rect 23793 13215 23959 13249
rect 23993 13215 24159 13249
rect 24193 13215 24359 13249
rect 24393 13215 24559 13249
rect 24593 13215 24759 13249
rect 24793 13215 24959 13249
rect 24993 13215 25159 13249
rect 25193 13215 25359 13249
rect 25393 13215 25559 13249
rect 25593 13215 25759 13249
rect 25793 13215 28443 13249
rect 28477 13215 28632 13249
rect 28684 13215 28843 13249
rect 28877 13215 29043 13249
rect 29077 13215 29243 13249
rect 29277 13215 29443 13249
rect 29477 13215 29643 13249
rect 29677 13215 29843 13249
rect 29877 13215 30043 13249
rect 30077 13215 30243 13249
rect 30277 13215 30443 13249
rect 30477 13215 30643 13249
rect 30677 13215 30843 13249
rect 30877 13215 31043 13249
rect 31077 13215 31243 13249
rect 31277 13215 31443 13249
rect 31477 13215 31643 13249
rect 31677 13215 31843 13249
rect 31877 13215 32043 13249
rect 32077 13215 32243 13249
rect 32277 13215 32443 13249
rect 32477 13215 32643 13249
rect 32677 13215 32843 13249
rect 32877 13215 33043 13249
rect 33077 13215 33243 13249
rect 33277 13215 33443 13249
rect 33477 13215 33643 13249
rect 33677 13215 33843 13249
rect 33877 13215 34043 13249
rect 34077 13215 34243 13249
rect 34277 13215 34443 13249
rect 34477 13215 34643 13249
rect 34677 13215 34843 13249
rect 34877 13215 35043 13249
rect 35077 13215 35243 13249
rect 35277 13215 35443 13249
rect 35477 13215 35643 13249
rect 35677 13215 35843 13249
rect 35877 13215 36043 13249
rect 36077 13215 36243 13249
rect 36277 13215 36443 13249
rect 36477 13215 36643 13249
rect 36677 13215 36843 13249
rect 36877 13215 37043 13249
rect 37077 13215 37243 13249
rect 37277 13215 37443 13249
rect 37477 13215 37643 13249
rect 37677 13215 37843 13249
rect 37877 13215 38043 13249
rect 38077 13215 38243 13249
rect 38277 13215 38443 13249
rect 38477 13215 38643 13249
rect 38677 13215 38843 13249
rect 38877 13215 39439 13249
rect 39473 13215 39639 13249
rect 39673 13215 39839 13249
rect 39873 13215 40039 13249
rect 40073 13215 40239 13249
rect 40273 13215 40439 13249
rect 40473 13215 40639 13249
rect 40673 13215 40839 13249
rect 40873 13215 41039 13249
rect 41073 13215 41239 13249
rect 41273 13215 41439 13249
rect 41473 13215 46126 13249
rect 17184 13200 28632 13215
rect 28684 13200 46126 13215
rect 2510 13174 46126 13200
rect 47714 13174 47736 13290
rect 900 13172 47736 13174
rect 10686 12492 10692 12504
rect 8220 12464 10692 12492
rect 8220 12436 8248 12464
rect 10686 12452 10692 12464
rect 10744 12452 10750 12504
rect 8202 12384 8208 12436
rect 8260 12384 8266 12436
rect 13722 11908 13728 11960
rect 13780 11948 13786 11960
rect 19426 11948 19432 11960
rect 13780 11920 19432 11948
rect 13780 11908 13786 11920
rect 19426 11908 19432 11920
rect 19484 11908 19490 11960
rect 13906 11636 13912 11688
rect 13964 11676 13970 11688
rect 20070 11676 20076 11688
rect 13964 11648 20076 11676
rect 13964 11636 13970 11648
rect 20070 11636 20076 11648
rect 20128 11636 20134 11688
rect 34054 11500 34060 11552
rect 34112 11540 34118 11552
rect 35434 11540 35440 11552
rect 34112 11512 35440 11540
rect 34112 11500 34118 11512
rect 35434 11500 35440 11512
rect 35492 11500 35498 11552
rect 3348 11410 45288 11412
rect 3348 11294 3370 11410
rect 4958 11369 43678 11410
rect 4958 11335 8079 11369
rect 8113 11335 8279 11369
rect 8313 11335 8479 11369
rect 8513 11335 8679 11369
rect 8713 11335 8879 11369
rect 8913 11335 9079 11369
rect 9113 11335 9279 11369
rect 9313 11335 9479 11369
rect 9513 11335 9679 11369
rect 9713 11335 9879 11369
rect 9913 11335 10079 11369
rect 10113 11335 10823 11369
rect 10857 11335 11023 11369
rect 11057 11335 11223 11369
rect 11257 11335 11423 11369
rect 11457 11335 11623 11369
rect 11657 11335 11823 11369
rect 11857 11335 12023 11369
rect 12057 11335 12223 11369
rect 12257 11335 12423 11369
rect 12457 11335 12623 11369
rect 12657 11335 12823 11369
rect 12857 11335 13567 11369
rect 13601 11335 13767 11369
rect 13801 11335 13967 11369
rect 14001 11335 14167 11369
rect 14201 11335 14367 11369
rect 14401 11335 14567 11369
rect 14601 11335 14767 11369
rect 14801 11335 14967 11369
rect 15001 11335 15167 11369
rect 15201 11335 15367 11369
rect 15401 11335 15567 11369
rect 15601 11335 16293 11369
rect 16327 11335 16693 11369
rect 16727 11335 17093 11369
rect 17127 11335 17493 11369
rect 17527 11335 17893 11369
rect 17927 11335 18293 11369
rect 18327 11335 18693 11369
rect 18727 11335 19093 11369
rect 19127 11335 19493 11369
rect 19527 11335 19893 11369
rect 19927 11335 20293 11369
rect 20327 11335 20693 11369
rect 20727 11335 21093 11369
rect 21127 11335 21493 11369
rect 21527 11335 21893 11369
rect 21927 11335 22293 11369
rect 22327 11335 22693 11369
rect 22727 11335 23093 11369
rect 23127 11335 23761 11369
rect 23795 11335 23961 11369
rect 23995 11335 24161 11369
rect 24195 11335 24361 11369
rect 24395 11335 24561 11369
rect 24595 11335 24761 11369
rect 24795 11335 24961 11369
rect 24995 11335 25161 11369
rect 25195 11335 25361 11369
rect 25395 11335 25561 11369
rect 25595 11335 25761 11369
rect 25795 11335 25961 11369
rect 25995 11335 26161 11369
rect 26195 11335 26361 11369
rect 26395 11335 27091 11369
rect 27125 11335 27291 11369
rect 27325 11335 27491 11369
rect 27525 11335 27691 11369
rect 27725 11335 27891 11369
rect 27925 11335 28091 11369
rect 28125 11335 28291 11369
rect 28325 11335 28491 11369
rect 28525 11335 28691 11369
rect 28725 11335 28891 11369
rect 28925 11335 29091 11369
rect 29125 11335 29835 11369
rect 29869 11335 30035 11369
rect 30069 11335 30235 11369
rect 30269 11335 30435 11369
rect 30469 11335 30635 11369
rect 30669 11335 30835 11369
rect 30869 11335 31035 11369
rect 31069 11335 31235 11369
rect 31269 11335 31435 11369
rect 31469 11335 31635 11369
rect 31669 11335 31835 11369
rect 31869 11335 32579 11369
rect 32613 11335 32779 11369
rect 32813 11335 32979 11369
rect 33013 11335 33179 11369
rect 33213 11335 33379 11369
rect 33413 11335 33579 11369
rect 33613 11335 33779 11369
rect 33813 11335 33979 11369
rect 34013 11335 34179 11369
rect 34213 11335 34379 11369
rect 34413 11335 34579 11369
rect 34613 11335 35323 11369
rect 35357 11335 35523 11369
rect 35557 11335 35723 11369
rect 35757 11335 35923 11369
rect 35957 11335 36123 11369
rect 36157 11335 36323 11369
rect 36357 11335 36523 11369
rect 36557 11335 36723 11369
rect 36757 11335 36923 11369
rect 36957 11335 37123 11369
rect 37157 11335 37323 11369
rect 37357 11335 38067 11369
rect 38101 11335 38267 11369
rect 38301 11335 38467 11369
rect 38501 11335 38667 11369
rect 38701 11335 38867 11369
rect 38901 11335 39067 11369
rect 39101 11335 39267 11369
rect 39301 11335 39467 11369
rect 39501 11335 39667 11369
rect 39701 11335 39867 11369
rect 39901 11335 40067 11369
rect 40101 11335 43678 11369
rect 4958 11294 43678 11335
rect 45266 11294 45288 11410
rect 3348 11292 45288 11294
rect 10980 11172 20576 11200
rect 10980 11113 11008 11172
rect 20548 11144 20576 11172
rect 23658 11160 23664 11212
rect 23716 11200 23722 11212
rect 23716 11172 29408 11200
rect 23716 11160 23722 11172
rect 7907 11101 8317 11113
rect 7907 10563 7915 11101
rect 8309 10563 8317 11101
rect 7907 10551 8317 10563
rect 9915 11101 10325 11113
rect 9915 10563 9922 11101
rect 10316 10563 10325 11101
rect 9915 10551 10325 10563
rect 10651 11101 11061 11113
rect 10651 10563 10659 11101
rect 11053 10563 11061 11101
rect 10651 10551 11061 10563
rect 12659 11101 13069 11113
rect 12659 10563 12666 11101
rect 13060 10563 13069 11101
rect 12659 10551 13069 10563
rect 13395 11101 13805 11113
rect 13395 10563 13403 11101
rect 13797 11064 13805 11101
rect 15403 11101 15813 11113
rect 13906 11064 13912 11076
rect 13797 11036 13912 11064
rect 13797 10563 13805 11036
rect 13906 11024 13912 11036
rect 13964 11024 13970 11076
rect 13395 10551 13805 10563
rect 15403 10563 15410 11101
rect 15804 10563 15813 11101
rect 20530 11092 20536 11144
rect 20588 11092 20594 11144
rect 23588 11101 23998 11113
rect 19426 11024 19432 11076
rect 19484 11064 19490 11076
rect 23588 11064 23596 11101
rect 19484 11036 23596 11064
rect 19484 11024 19490 11036
rect 15403 10551 15813 10563
rect 23588 10563 23596 11036
rect 23990 10563 23998 11101
rect 23588 10551 23998 10563
rect 26170 11101 26580 11113
rect 26170 10563 26177 11101
rect 26571 10563 26580 11101
rect 26170 10551 26580 10563
rect 26919 11101 27329 11113
rect 26919 10563 26927 11101
rect 27321 10588 27329 11101
rect 28927 11101 29337 11113
rect 28810 10588 28816 10600
rect 27321 10563 28816 10588
rect 26919 10560 28816 10563
rect 26919 10551 27329 10560
rect 7907 10141 8317 10153
rect 7907 9603 7915 10141
rect 8309 9636 8317 10141
rect 9904 10141 10336 10551
rect 9766 9636 9772 9648
rect 8309 9608 9772 9636
rect 8309 9603 8317 9608
rect 7907 9591 8317 9603
rect 9766 9596 9772 9608
rect 9824 9596 9830 9648
rect 9904 9603 9922 10141
rect 10316 9603 10336 10141
rect 9904 9587 10336 9603
rect 10651 10141 11061 10153
rect 10651 9603 10659 10141
rect 11053 9636 11061 10141
rect 12648 10141 13080 10551
rect 12526 9636 12532 9648
rect 11053 9608 12532 9636
rect 11053 9603 11061 9608
rect 10651 9591 11061 9603
rect 12526 9596 12532 9608
rect 12584 9596 12590 9648
rect 12648 9603 12666 10141
rect 13060 9603 13080 10141
rect 12648 9587 13080 9603
rect 13395 10141 13805 10153
rect 13395 9603 13403 10141
rect 13797 9636 13805 10141
rect 15392 10141 15824 10551
rect 13906 9636 13912 9648
rect 13797 9608 13912 9636
rect 13797 9603 13805 9608
rect 13395 9591 13805 9603
rect 13906 9596 13912 9608
rect 13964 9596 13970 9648
rect 15392 9603 15410 10141
rect 15804 9603 15824 10141
rect 15392 9587 15824 9603
rect 23588 10141 23998 10153
rect 23588 9603 23596 10141
rect 23990 9603 23998 10141
rect 23588 9591 23998 9603
rect 26159 10141 26591 10551
rect 28810 10548 28816 10560
rect 28868 10548 28874 10600
rect 28927 10563 28934 11101
rect 29328 10563 29337 11101
rect 29380 11064 29408 11172
rect 31496 11172 37688 11200
rect 31496 11144 31524 11172
rect 29663 11101 30073 11113
rect 29663 11064 29671 11101
rect 29380 11036 29671 11064
rect 28927 10551 29337 10563
rect 29663 10563 29671 11036
rect 30065 10563 30073 11101
rect 31478 11092 31484 11144
rect 31536 11092 31542 11144
rect 31671 11101 32081 11113
rect 29663 10551 30073 10563
rect 31671 10563 31678 11101
rect 32072 10563 32081 11101
rect 31671 10551 32081 10563
rect 32407 11101 32817 11113
rect 32407 10563 32415 11101
rect 32809 11064 32817 11101
rect 34415 11101 34825 11113
rect 34054 11064 34060 11076
rect 32809 11036 34060 11064
rect 32809 10563 32817 11036
rect 34054 11024 34060 11036
rect 34112 11024 34118 11076
rect 32407 10551 32817 10563
rect 34415 10563 34422 11101
rect 34816 10563 34825 11101
rect 34415 10551 34825 10563
rect 35151 11101 35561 11113
rect 35151 10563 35159 11101
rect 35553 10588 35561 11101
rect 37159 11101 37569 11113
rect 36998 10588 37004 10600
rect 35553 10563 37004 10588
rect 35151 10560 37004 10563
rect 35151 10551 35561 10560
rect 26159 9603 26177 10141
rect 26571 9603 26591 10141
rect 23952 9532 23980 9591
rect 26159 9587 26591 9603
rect 26919 10141 27329 10153
rect 26919 9603 26927 10141
rect 27321 9636 27329 10141
rect 28916 10141 29348 10551
rect 28534 9636 28540 9648
rect 27321 9608 28540 9636
rect 27321 9603 27329 9608
rect 26919 9591 27329 9603
rect 28534 9596 28540 9608
rect 28592 9596 28598 9648
rect 28916 9603 28934 10141
rect 29328 9603 29348 10141
rect 29663 10141 30073 10153
rect 29454 10072 29460 10124
rect 29512 10112 29518 10124
rect 29663 10112 29671 10141
rect 29512 10084 29671 10112
rect 29512 10072 29518 10084
rect 28916 9587 29348 9603
rect 29663 9603 29671 10084
rect 30065 9603 30073 10141
rect 29663 9591 30073 9603
rect 31660 10141 32092 10551
rect 31660 9603 31678 10141
rect 32072 9603 32092 10141
rect 32407 10141 32817 10153
rect 31660 9587 32092 9603
rect 32122 9596 32128 9648
rect 32180 9636 32186 9648
rect 32407 9636 32415 10141
rect 32180 9608 32415 9636
rect 32180 9596 32186 9608
rect 32407 9603 32415 9608
rect 32809 9603 32817 10141
rect 32407 9591 32817 9603
rect 34404 10141 34836 10551
rect 36998 10548 37004 10560
rect 37056 10548 37062 10600
rect 37159 10563 37166 11101
rect 37560 10563 37569 11101
rect 37660 11064 37688 11172
rect 37895 11101 38305 11113
rect 37895 11064 37903 11101
rect 37660 11036 37903 11064
rect 37159 10551 37569 10563
rect 37895 10563 37903 11036
rect 38297 10563 38305 11101
rect 37895 10551 38305 10563
rect 39903 11101 40313 11113
rect 39903 10563 39910 11101
rect 40304 10563 40313 11101
rect 39903 10551 40313 10563
rect 34404 9603 34422 10141
rect 34816 9603 34836 10141
rect 35151 10141 35561 10153
rect 34404 9587 34836 9603
rect 34974 9596 34980 9648
rect 35032 9636 35038 9648
rect 35151 9636 35159 10141
rect 35032 9608 35159 9636
rect 35032 9596 35038 9608
rect 35151 9603 35159 9608
rect 35553 9603 35561 10141
rect 35151 9591 35561 9603
rect 37148 10141 37580 10551
rect 37148 9603 37166 10141
rect 37560 9603 37580 10141
rect 37895 10141 38305 10153
rect 37148 9587 37580 9603
rect 37642 9596 37648 9648
rect 37700 9636 37706 9648
rect 37895 9636 37903 10141
rect 37700 9608 37903 9636
rect 37700 9596 37706 9608
rect 37895 9603 37903 9608
rect 38297 9603 38305 10141
rect 37895 9591 38305 9603
rect 39892 10141 40324 10551
rect 39892 9603 39910 10141
rect 40304 9603 40324 10141
rect 39892 9587 40324 9603
rect 900 9530 47736 9532
rect 900 9414 922 9530
rect 2510 9512 46126 9530
rect 2510 9489 17132 9512
rect 2510 9455 8079 9489
rect 8113 9455 8279 9489
rect 8313 9455 8479 9489
rect 8513 9455 8679 9489
rect 8713 9455 8879 9489
rect 8913 9455 9079 9489
rect 9113 9455 9279 9489
rect 9313 9455 9479 9489
rect 9513 9455 9679 9489
rect 9713 9455 9879 9489
rect 9913 9455 10079 9489
rect 10113 9455 10823 9489
rect 10857 9455 11023 9489
rect 11057 9455 11223 9489
rect 11257 9455 11423 9489
rect 11457 9455 11623 9489
rect 11657 9455 11823 9489
rect 11857 9455 12023 9489
rect 12057 9455 12223 9489
rect 12257 9455 12423 9489
rect 12457 9455 12623 9489
rect 12657 9455 12823 9489
rect 12857 9455 13567 9489
rect 13601 9455 13767 9489
rect 13801 9455 13967 9489
rect 14001 9455 14167 9489
rect 14201 9455 14367 9489
rect 14401 9455 14567 9489
rect 14601 9455 14767 9489
rect 14801 9455 14967 9489
rect 15001 9455 15167 9489
rect 15201 9455 15367 9489
rect 15401 9455 15567 9489
rect 15601 9455 16293 9489
rect 16327 9455 16693 9489
rect 16727 9455 17093 9489
rect 17127 9460 17132 9489
rect 17184 9489 46126 9512
rect 17184 9460 17493 9489
rect 17127 9455 17493 9460
rect 17527 9455 17893 9489
rect 17927 9455 18293 9489
rect 18327 9455 18693 9489
rect 18727 9455 19093 9489
rect 19127 9455 19493 9489
rect 19527 9455 19893 9489
rect 19927 9455 20293 9489
rect 20327 9455 20693 9489
rect 20727 9455 21093 9489
rect 21127 9455 21493 9489
rect 21527 9455 21893 9489
rect 21927 9455 22293 9489
rect 22327 9455 22693 9489
rect 22727 9455 23093 9489
rect 23127 9455 23761 9489
rect 23795 9455 23961 9489
rect 23995 9455 24161 9489
rect 24195 9455 24361 9489
rect 24395 9455 24561 9489
rect 24595 9455 24761 9489
rect 24795 9455 24961 9489
rect 24995 9455 25161 9489
rect 25195 9455 25361 9489
rect 25395 9455 25561 9489
rect 25595 9455 25761 9489
rect 25795 9455 25961 9489
rect 25995 9455 26161 9489
rect 26195 9455 26361 9489
rect 26395 9455 27091 9489
rect 27125 9455 27291 9489
rect 27325 9455 27491 9489
rect 27525 9455 27691 9489
rect 27725 9455 27891 9489
rect 27925 9455 28091 9489
rect 28125 9455 28291 9489
rect 28325 9455 28491 9489
rect 28525 9455 28691 9489
rect 28725 9455 28891 9489
rect 28925 9455 29091 9489
rect 29125 9455 29835 9489
rect 29869 9455 30035 9489
rect 30069 9455 30235 9489
rect 30269 9455 30435 9489
rect 30469 9455 30635 9489
rect 30669 9455 30835 9489
rect 30869 9455 31035 9489
rect 31069 9455 31235 9489
rect 31269 9455 31435 9489
rect 31469 9455 31635 9489
rect 31669 9455 31835 9489
rect 31869 9455 32579 9489
rect 32613 9455 32779 9489
rect 32813 9455 32979 9489
rect 33013 9455 33179 9489
rect 33213 9455 33379 9489
rect 33413 9455 33579 9489
rect 33613 9455 33779 9489
rect 33813 9455 33979 9489
rect 34013 9455 34179 9489
rect 34213 9455 34379 9489
rect 34413 9455 34579 9489
rect 34613 9455 35323 9489
rect 35357 9455 35523 9489
rect 35557 9455 35723 9489
rect 35757 9455 35923 9489
rect 35957 9455 36123 9489
rect 36157 9455 36323 9489
rect 36357 9455 36523 9489
rect 36557 9455 36723 9489
rect 36757 9455 36923 9489
rect 36957 9455 37123 9489
rect 37157 9455 37323 9489
rect 37357 9455 38067 9489
rect 38101 9455 38267 9489
rect 38301 9455 38467 9489
rect 38501 9455 38667 9489
rect 38701 9455 38867 9489
rect 38901 9455 39067 9489
rect 39101 9455 39267 9489
rect 39301 9455 39467 9489
rect 39501 9455 39667 9489
rect 39701 9455 39867 9489
rect 39901 9455 40067 9489
rect 40101 9455 46126 9489
rect 2510 9414 46126 9455
rect 47714 9414 47736 9530
rect 900 9412 47736 9414
rect 32490 9324 32496 9376
rect 32548 9364 32554 9376
rect 34974 9364 34980 9376
rect 32548 9336 34980 9364
rect 32548 9324 32554 9336
rect 34974 9324 34980 9336
rect 35032 9324 35038 9376
rect 36998 9324 37004 9376
rect 37056 9364 37062 9376
rect 38102 9364 38108 9376
rect 37056 9336 38108 9364
rect 37056 9324 37062 9336
rect 38102 9324 38108 9336
rect 38160 9324 38166 9376
rect 14734 9188 14740 9240
rect 14792 9228 14798 9240
rect 32122 9228 32128 9240
rect 14792 9200 32128 9228
rect 14792 9188 14798 9200
rect 32122 9188 32128 9200
rect 32180 9188 32186 9240
rect 12526 8916 12532 8968
rect 12584 8956 12590 8968
rect 23198 8956 23204 8968
rect 12584 8928 23204 8956
rect 12584 8916 12590 8928
rect 23198 8916 23204 8928
rect 23256 8916 23262 8968
rect 3348 7650 45288 7652
rect 3348 7534 3370 7650
rect 4958 7609 43678 7650
rect 4958 7575 8079 7609
rect 8113 7575 8279 7609
rect 8313 7575 8479 7609
rect 8513 7575 8679 7609
rect 8713 7575 8879 7609
rect 8913 7575 9079 7609
rect 9113 7575 9279 7609
rect 9313 7575 9479 7609
rect 9513 7575 9679 7609
rect 9713 7575 9879 7609
rect 9913 7575 10079 7609
rect 10113 7575 14451 7609
rect 14485 7575 14651 7609
rect 14685 7575 14851 7609
rect 14885 7575 15051 7609
rect 15085 7575 15251 7609
rect 15285 7575 15451 7609
rect 15485 7575 15651 7609
rect 15685 7575 15851 7609
rect 15885 7575 16051 7609
rect 16085 7575 16251 7609
rect 16285 7575 16451 7609
rect 16485 7575 16651 7609
rect 16685 7575 16851 7609
rect 16885 7575 17051 7609
rect 17085 7575 17781 7609
rect 17815 7575 17981 7609
rect 18015 7575 18181 7609
rect 18215 7575 18381 7609
rect 18415 7575 18581 7609
rect 18615 7575 18781 7609
rect 18815 7575 18981 7609
rect 19015 7575 19181 7609
rect 19215 7575 19381 7609
rect 19415 7575 19581 7609
rect 19615 7575 19781 7609
rect 19815 7575 20525 7609
rect 20559 7575 20725 7609
rect 20759 7575 20925 7609
rect 20959 7575 21125 7609
rect 21159 7575 21325 7609
rect 21359 7575 21525 7609
rect 21559 7575 21725 7609
rect 21759 7575 21925 7609
rect 21959 7575 22125 7609
rect 22159 7575 22325 7609
rect 22359 7575 22525 7609
rect 22559 7575 23269 7609
rect 23303 7575 23469 7609
rect 23503 7575 23669 7609
rect 23703 7575 23869 7609
rect 23903 7575 24069 7609
rect 24103 7575 24269 7609
rect 24303 7575 24469 7609
rect 24503 7575 24669 7609
rect 24703 7575 24869 7609
rect 24903 7575 25069 7609
rect 25103 7575 25269 7609
rect 25303 7575 26013 7609
rect 26047 7575 26213 7609
rect 26247 7575 26413 7609
rect 26447 7575 26613 7609
rect 26647 7575 26813 7609
rect 26847 7575 27013 7609
rect 27047 7575 27213 7609
rect 27247 7575 27413 7609
rect 27447 7575 27613 7609
rect 27647 7575 27813 7609
rect 27847 7575 28013 7609
rect 28047 7575 28757 7609
rect 28791 7575 28957 7609
rect 28991 7575 29157 7609
rect 29191 7575 29357 7609
rect 29391 7575 29557 7609
rect 29591 7575 29757 7609
rect 29791 7575 29957 7609
rect 29991 7575 30157 7609
rect 30191 7575 30357 7609
rect 30391 7575 30557 7609
rect 30591 7575 30757 7609
rect 30791 7575 31501 7609
rect 31535 7575 31701 7609
rect 31735 7575 31901 7609
rect 31935 7575 32101 7609
rect 32135 7575 32301 7609
rect 32335 7575 32501 7609
rect 32535 7575 32701 7609
rect 32735 7575 32901 7609
rect 32935 7575 33101 7609
rect 33135 7575 33301 7609
rect 33335 7575 33501 7609
rect 33535 7575 35323 7609
rect 35357 7575 35523 7609
rect 35557 7575 35723 7609
rect 35757 7575 35923 7609
rect 35957 7575 36123 7609
rect 36157 7575 36323 7609
rect 36357 7575 36523 7609
rect 36557 7575 36723 7609
rect 36757 7575 36923 7609
rect 36957 7575 37123 7609
rect 37157 7575 37323 7609
rect 37357 7575 38067 7609
rect 38101 7575 38267 7609
rect 38301 7575 38467 7609
rect 38501 7575 38667 7609
rect 38701 7575 38867 7609
rect 38901 7575 39067 7609
rect 39101 7575 39267 7609
rect 39301 7575 39467 7609
rect 39501 7575 39667 7609
rect 39701 7575 39867 7609
rect 39901 7575 40067 7609
rect 40101 7575 43678 7609
rect 4958 7534 43678 7575
rect 45266 7534 45288 7650
rect 3348 7532 45288 7534
rect 25590 7460 25596 7472
rect 22296 7432 25596 7460
rect 8202 7353 8208 7404
rect 7907 7352 8208 7353
rect 8260 7353 8266 7404
rect 8260 7352 8317 7353
rect 7907 7341 8317 7352
rect 7907 6803 7915 7341
rect 8309 6803 8317 7341
rect 7907 6791 8317 6803
rect 9915 7341 10325 7353
rect 9915 6803 9922 7341
rect 10316 6803 10325 7341
rect 14278 7341 14688 7353
rect 13906 7284 13912 7336
rect 13964 7324 13970 7336
rect 14278 7324 14286 7341
rect 13964 7296 14286 7324
rect 13964 7284 13970 7296
rect 9915 6791 10325 6803
rect 14278 6803 14286 7296
rect 14680 6803 14688 7341
rect 14278 6791 14688 6803
rect 16860 7341 17270 7353
rect 16860 6803 16867 7341
rect 17261 6803 17270 7341
rect 16860 6791 17270 6803
rect 17609 7341 18019 7353
rect 17609 6803 17617 7341
rect 18011 6803 18019 7341
rect 17609 6791 18019 6803
rect 19617 7341 20027 7353
rect 19617 6803 19624 7341
rect 20018 6803 20027 7341
rect 19617 6791 20027 6803
rect 20353 7341 20763 7353
rect 20353 6803 20361 7341
rect 20755 7324 20763 7341
rect 22296 7324 22324 7432
rect 25590 7420 25596 7432
rect 25648 7420 25654 7472
rect 37642 7460 37648 7472
rect 37016 7432 37648 7460
rect 20755 7296 22324 7324
rect 22361 7341 22771 7353
rect 20755 6803 20763 7296
rect 20353 6791 20763 6803
rect 22361 6803 22368 7341
rect 22762 6803 22771 7341
rect 22361 6791 22771 6803
rect 23097 7341 23507 7353
rect 23097 6803 23105 7341
rect 23499 6803 23507 7341
rect 23097 6791 23507 6803
rect 25105 7341 25515 7353
rect 25105 6803 25112 7341
rect 25506 6803 25515 7341
rect 25841 7341 26251 7353
rect 25682 6808 25688 6860
rect 25740 6848 25746 6860
rect 25841 6848 25849 7341
rect 25740 6820 25849 6848
rect 25740 6808 25746 6820
rect 25105 6791 25515 6803
rect 25841 6803 25849 6820
rect 26243 6803 26251 7341
rect 25841 6791 26251 6803
rect 27849 7341 28259 7353
rect 27849 6803 27856 7341
rect 28250 6803 28259 7341
rect 28585 7341 28995 7353
rect 28585 7336 28593 7341
rect 28534 7284 28540 7336
rect 28592 7284 28593 7336
rect 27849 6791 28259 6803
rect 28585 6803 28593 7284
rect 28987 6803 28995 7341
rect 28585 6791 28995 6803
rect 30593 7341 31003 7353
rect 30593 6803 30600 7341
rect 30994 6803 31003 7341
rect 30593 6791 31003 6803
rect 31329 7341 31739 7353
rect 31329 6803 31337 7341
rect 31731 7324 31739 7341
rect 33337 7341 33747 7353
rect 32490 7324 32496 7336
rect 31731 7296 32496 7324
rect 31731 6803 31739 7296
rect 32490 7284 32496 7296
rect 32548 7284 32554 7336
rect 31329 6791 31739 6803
rect 33337 6803 33344 7341
rect 33738 6803 33747 7341
rect 33337 6791 33747 6803
rect 35151 7341 35561 7353
rect 35151 6803 35159 7341
rect 35553 7324 35561 7341
rect 37016 7324 37044 7432
rect 37642 7420 37648 7432
rect 37700 7420 37706 7472
rect 38194 7353 38200 7404
rect 35553 7296 37044 7324
rect 37159 7341 37569 7353
rect 35553 6803 35561 7296
rect 35151 6791 35561 6803
rect 37159 6803 37166 7341
rect 37560 6803 37569 7341
rect 37159 6791 37569 6803
rect 37895 7352 38200 7353
rect 38252 7353 38258 7404
rect 38252 7352 38305 7353
rect 37895 7341 38305 7352
rect 37895 6803 37903 7341
rect 38297 6803 38305 7341
rect 37895 6791 38305 6803
rect 39903 7341 40313 7353
rect 39903 6803 39910 7341
rect 40304 6803 40313 7341
rect 39903 6791 40313 6803
rect 8110 6468 8116 6520
rect 8168 6468 8174 6520
rect 8128 6393 8156 6468
rect 7907 6381 8317 6393
rect 7907 5843 7915 6381
rect 8309 5843 8317 6381
rect 7907 5831 8317 5843
rect 9904 6381 10336 6791
rect 9904 5843 9922 6381
rect 10316 5843 10336 6381
rect 9904 5827 10336 5843
rect 14278 6381 14688 6393
rect 14278 5843 14286 6381
rect 14680 5843 14688 6381
rect 14278 5831 14688 5843
rect 16849 6381 17281 6791
rect 16849 5843 16867 6381
rect 17261 5843 17281 6381
rect 14292 5772 14320 5831
rect 16849 5827 17281 5843
rect 17609 6381 18019 6393
rect 17609 5843 17617 6381
rect 18011 6372 18019 6381
rect 19524 6384 19576 6390
rect 18011 6344 19524 6372
rect 18011 5843 18019 6344
rect 19524 6326 19576 6332
rect 19606 6381 20038 6791
rect 17609 5831 18019 5843
rect 19606 5843 19624 6381
rect 20018 5843 20038 6381
rect 19606 5827 20038 5843
rect 20353 6384 20763 6393
rect 20353 6381 20536 6384
rect 20588 6381 20763 6384
rect 20353 5843 20361 6381
rect 20755 5843 20763 6381
rect 20353 5831 20763 5843
rect 22350 6381 22782 6791
rect 22350 5843 22368 6381
rect 22762 5843 22782 6381
rect 22350 5827 22782 5843
rect 23097 6381 23507 6393
rect 23097 5843 23105 6381
rect 23499 6372 23507 6381
rect 23566 6372 23572 6384
rect 23499 6344 23572 6372
rect 23499 5843 23507 6344
rect 23566 6332 23572 6344
rect 23624 6332 23630 6384
rect 25094 6381 25526 6791
rect 23097 5831 23507 5843
rect 25094 5843 25112 6381
rect 25506 5843 25526 6381
rect 25590 6332 25596 6384
rect 25648 6372 25654 6384
rect 25841 6381 26251 6393
rect 25841 6372 25849 6381
rect 25648 6344 25849 6372
rect 25648 6332 25654 6344
rect 25094 5827 25526 5843
rect 25841 5843 25849 6344
rect 26243 5843 26251 6381
rect 25841 5831 26251 5843
rect 27838 6381 28270 6791
rect 27838 5843 27856 6381
rect 28250 5843 28270 6381
rect 28585 6381 28995 6393
rect 28350 6060 28356 6112
rect 28408 6100 28414 6112
rect 28585 6100 28593 6381
rect 28408 6072 28593 6100
rect 28408 6060 28414 6072
rect 27838 5827 28270 5843
rect 28585 5843 28593 6072
rect 28987 5843 28995 6381
rect 28585 5831 28995 5843
rect 30582 6381 31014 6791
rect 30582 5843 30600 6381
rect 30994 5843 31014 6381
rect 30582 5827 31014 5843
rect 31329 6384 31739 6393
rect 31329 6381 31484 6384
rect 31536 6381 31739 6384
rect 31329 5843 31337 6381
rect 31731 5843 31739 6381
rect 31329 5831 31739 5843
rect 33326 6381 33758 6791
rect 35342 6468 35348 6520
rect 35400 6468 35406 6520
rect 35360 6393 35388 6468
rect 33326 5843 33344 6381
rect 33738 5843 33758 6381
rect 33326 5827 33758 5843
rect 35151 6381 35561 6393
rect 35151 5843 35159 6381
rect 35553 5843 35561 6381
rect 35151 5831 35561 5843
rect 37148 6381 37580 6791
rect 38102 6468 38108 6520
rect 38160 6468 38166 6520
rect 38120 6393 38148 6468
rect 37148 5843 37166 6381
rect 37560 5843 37580 6381
rect 37148 5827 37580 5843
rect 37895 6381 38305 6393
rect 37895 5843 37903 6381
rect 38297 5843 38305 6381
rect 37895 5831 38305 5843
rect 39892 6381 40324 6791
rect 39892 5843 39910 6381
rect 40304 5843 40324 6381
rect 39892 5827 40324 5843
rect 900 5770 47736 5772
rect 900 5654 922 5770
rect 2510 5729 46126 5770
rect 2510 5695 8079 5729
rect 8113 5695 8279 5729
rect 8313 5695 8479 5729
rect 8513 5695 8679 5729
rect 8713 5695 8879 5729
rect 8913 5695 9079 5729
rect 9113 5695 9279 5729
rect 9313 5695 9479 5729
rect 9513 5695 9679 5729
rect 9713 5695 9879 5729
rect 9913 5695 10079 5729
rect 10113 5695 14451 5729
rect 14485 5695 14651 5729
rect 14685 5695 14851 5729
rect 14885 5695 15051 5729
rect 15085 5695 15251 5729
rect 15285 5695 15451 5729
rect 15485 5695 15651 5729
rect 15685 5695 15851 5729
rect 15885 5695 16051 5729
rect 16085 5695 16251 5729
rect 16285 5695 16451 5729
rect 16485 5695 16651 5729
rect 16685 5695 16851 5729
rect 16885 5695 17051 5729
rect 17085 5695 17781 5729
rect 17815 5695 17981 5729
rect 18015 5695 18181 5729
rect 18215 5695 18381 5729
rect 18415 5695 18581 5729
rect 18615 5695 18781 5729
rect 18815 5695 18981 5729
rect 19015 5695 19181 5729
rect 19215 5695 19381 5729
rect 19415 5695 19581 5729
rect 19615 5695 19781 5729
rect 19815 5695 20525 5729
rect 20559 5695 20725 5729
rect 20759 5695 20925 5729
rect 20959 5695 21125 5729
rect 21159 5695 21325 5729
rect 21359 5695 21525 5729
rect 21559 5695 21725 5729
rect 21759 5695 21925 5729
rect 21959 5695 22125 5729
rect 22159 5695 22325 5729
rect 22359 5695 22525 5729
rect 22559 5695 23269 5729
rect 23303 5695 23469 5729
rect 23503 5695 23669 5729
rect 23703 5695 23869 5729
rect 23903 5695 24069 5729
rect 24103 5695 24269 5729
rect 24303 5695 24469 5729
rect 24503 5695 24669 5729
rect 24703 5695 24869 5729
rect 24903 5695 25069 5729
rect 25103 5695 25269 5729
rect 25303 5695 26013 5729
rect 26047 5695 26213 5729
rect 26247 5695 26413 5729
rect 26447 5695 26613 5729
rect 26647 5695 26813 5729
rect 26847 5695 27013 5729
rect 27047 5695 27213 5729
rect 27247 5695 27413 5729
rect 27447 5695 27613 5729
rect 27647 5695 27813 5729
rect 27847 5695 28013 5729
rect 28047 5695 28757 5729
rect 28791 5695 28957 5729
rect 28991 5695 29157 5729
rect 29191 5695 29357 5729
rect 29391 5695 29557 5729
rect 29591 5695 29757 5729
rect 29791 5695 29957 5729
rect 29991 5695 30157 5729
rect 30191 5695 30357 5729
rect 30391 5695 30557 5729
rect 30591 5695 30757 5729
rect 30791 5695 31501 5729
rect 31535 5695 31701 5729
rect 31735 5695 31901 5729
rect 31935 5695 32101 5729
rect 32135 5695 32301 5729
rect 32335 5695 32501 5729
rect 32535 5695 32701 5729
rect 32735 5695 32901 5729
rect 32935 5695 33101 5729
rect 33135 5695 33301 5729
rect 33335 5695 33501 5729
rect 33535 5695 35323 5729
rect 35357 5695 35523 5729
rect 35557 5695 35723 5729
rect 35757 5695 35923 5729
rect 35957 5695 36123 5729
rect 36157 5695 36323 5729
rect 36357 5695 36523 5729
rect 36557 5695 36723 5729
rect 36757 5695 36923 5729
rect 36957 5695 37123 5729
rect 37157 5695 37323 5729
rect 37357 5695 38067 5729
rect 38101 5695 38267 5729
rect 38301 5695 38467 5729
rect 38501 5695 38667 5729
rect 38701 5695 38867 5729
rect 38901 5695 39067 5729
rect 39101 5695 39267 5729
rect 39301 5695 39467 5729
rect 39501 5695 39667 5729
rect 39701 5695 39867 5729
rect 39901 5695 40067 5729
rect 40101 5695 46126 5729
rect 2510 5654 46126 5695
rect 47714 5654 47736 5770
rect 900 5652 47736 5654
<< via1 >>
rect 3370 41374 4958 41490
rect 12440 41420 12492 41472
rect 43678 41374 45266 41490
rect 27344 41148 27396 41200
rect 38660 39831 38712 39840
rect 38660 39797 38669 39831
rect 38669 39797 38703 39831
rect 38703 39797 38712 39831
rect 38660 39788 38712 39797
rect 9588 39652 9640 39704
rect 15016 39695 15068 39704
rect 15016 39661 15025 39695
rect 15025 39661 15059 39695
rect 15059 39661 15068 39695
rect 15016 39652 15068 39661
rect 27620 39695 27672 39704
rect 27620 39661 27629 39695
rect 27629 39661 27663 39695
rect 27663 39661 27672 39695
rect 27620 39652 27672 39661
rect 922 39494 2510 39610
rect 46126 39494 47714 39610
rect 3370 37614 4958 37730
rect 12992 37612 13044 37664
rect 16856 37612 16908 37664
rect 27896 37612 27948 37664
rect 43678 37614 45266 37730
rect 30196 37162 30234 37188
rect 30234 37162 30248 37188
rect 30196 37136 30248 37162
rect 39948 36728 40000 36780
rect 31668 36456 31720 36508
rect 26240 36116 26292 36168
rect 9588 36048 9640 36100
rect 922 35734 2510 35850
rect 30196 35809 30248 35828
rect 30196 35776 30207 35809
rect 30207 35776 30241 35809
rect 30241 35776 30248 35809
rect 46126 35734 47714 35850
rect 3370 33854 4958 33970
rect 9956 33895 9987 33924
rect 9987 33895 10008 33924
rect 9956 33872 10008 33895
rect 43678 33854 45266 33970
rect 40040 32376 40092 32428
rect 26884 32283 26936 32292
rect 26884 32249 26893 32283
rect 26893 32249 26927 32283
rect 26927 32249 26936 32283
rect 26884 32240 26936 32249
rect 14188 32181 14240 32224
rect 14188 32172 14197 32181
rect 14197 32172 14231 32181
rect 14231 32172 14240 32181
rect 922 31974 2510 32090
rect 46126 31974 47714 32090
rect 3370 30094 4958 30210
rect 43678 30094 45266 30210
rect 18880 28677 18932 28688
rect 18880 28643 18885 28677
rect 18885 28643 18919 28677
rect 18919 28643 18932 28677
rect 18880 28636 18932 28643
rect 26516 28500 26568 28552
rect 40040 29860 40092 29912
rect 12532 28407 12584 28416
rect 12532 28373 12541 28407
rect 12541 28373 12575 28407
rect 12575 28373 12584 28407
rect 12532 28364 12584 28373
rect 14188 28407 14240 28416
rect 14188 28373 14197 28407
rect 14197 28373 14231 28407
rect 14231 28373 14240 28407
rect 14188 28364 14240 28373
rect 23388 28407 23440 28416
rect 23388 28373 23397 28407
rect 23397 28373 23431 28407
rect 23431 28373 23440 28407
rect 23388 28364 23440 28373
rect 39304 28908 39356 28960
rect 40040 28432 40092 28484
rect 922 28214 2510 28330
rect 46126 28214 47714 28330
rect 3370 26334 4958 26450
rect 43678 26334 45266 26450
rect 7104 25603 7133 25628
rect 7133 25603 7156 25628
rect 7104 25576 7156 25603
rect 9588 26141 9640 26172
rect 9588 26120 9589 26141
rect 9589 26120 9623 26141
rect 9623 26120 9640 26141
rect 26240 26188 26292 26240
rect 7196 24624 7248 24676
rect 31668 25712 31720 25764
rect 28632 25212 28684 25220
rect 28632 25178 28656 25212
rect 28656 25178 28684 25212
rect 28632 25168 28684 25178
rect 39396 25644 39448 25696
rect 23388 25007 23440 25016
rect 23388 24973 23397 25007
rect 23397 24973 23431 25007
rect 23431 24973 23440 25007
rect 23388 24964 23440 24973
rect 39396 24896 39448 24948
rect 23296 24871 23348 24880
rect 23296 24837 23305 24871
rect 23305 24837 23339 24871
rect 23339 24837 23348 24871
rect 23296 24828 23348 24837
rect 27620 24828 27672 24880
rect 9680 24667 9732 24676
rect 9680 24633 9689 24667
rect 9689 24633 9723 24667
rect 9723 24633 9732 24667
rect 9680 24624 9732 24633
rect 12532 24667 12584 24676
rect 12532 24633 12541 24667
rect 12541 24633 12575 24667
rect 12575 24633 12584 24667
rect 12532 24624 12584 24633
rect 922 24454 2510 24570
rect 15476 24488 15528 24540
rect 46126 24454 47714 24570
rect 7196 24216 7248 24268
rect 13360 24216 13412 24268
rect 7104 23468 7156 23520
rect 30104 23468 30156 23520
rect 3370 22574 4958 22690
rect 43678 22574 45266 22690
rect 8300 22491 8352 22500
rect 8300 22457 8309 22491
rect 8309 22457 8343 22491
rect 8343 22457 8352 22491
rect 8300 22448 8352 22457
rect 26424 22491 26476 22500
rect 26424 22457 26433 22491
rect 26433 22457 26467 22491
rect 26467 22457 26476 22491
rect 26424 22448 26476 22457
rect 38660 22380 38712 22432
rect 23296 22176 23348 22228
rect 20904 21564 20956 21616
rect 30564 22108 30616 22160
rect 28632 21972 28684 22024
rect 28724 21360 28776 21412
rect 26516 21267 26568 21276
rect 26516 21233 26525 21267
rect 26525 21233 26559 21267
rect 26559 21233 26568 21267
rect 26516 21224 26568 21233
rect 30104 21156 30156 21208
rect 26884 21131 26936 21140
rect 13268 20995 13320 21004
rect 13268 20961 13277 20995
rect 13277 20961 13311 20995
rect 13311 20961 13320 20995
rect 13268 20952 13320 20961
rect 8300 20927 8352 20936
rect 8300 20893 8309 20927
rect 8309 20893 8343 20927
rect 8343 20893 8352 20927
rect 8300 20884 8352 20893
rect 26884 21097 26893 21131
rect 26893 21097 26927 21131
rect 26927 21097 26936 21131
rect 26884 21088 26936 21097
rect 922 20694 2510 20810
rect 14096 20769 14148 20800
rect 14096 20748 14145 20769
rect 14145 20748 14148 20769
rect 30564 20748 30616 20800
rect 46126 20694 47714 20810
rect 3370 18814 4958 18930
rect 43678 18814 45266 18930
rect 9680 18335 9690 18352
rect 9690 18335 9724 18352
rect 9724 18335 9732 18352
rect 9680 18300 9732 18335
rect 12532 18096 12584 18148
rect 13360 18621 13412 18624
rect 13360 18572 13403 18621
rect 13403 18572 13412 18621
rect 8760 17144 8812 17196
rect 13176 17620 13228 17672
rect 39488 18621 39540 18624
rect 28632 18396 28684 18420
rect 28632 18368 28650 18396
rect 28650 18368 28684 18396
rect 28724 18192 28776 18216
rect 28724 18164 28756 18192
rect 28756 18164 28776 18192
rect 39488 18572 39540 18621
rect 28724 17658 28756 17672
rect 28756 17658 28776 17672
rect 28724 17620 28776 17658
rect 23388 17280 23440 17332
rect 26516 17153 26568 17196
rect 26516 17144 26525 17153
rect 26525 17144 26559 17153
rect 26559 17144 26568 17153
rect 39304 17144 39356 17196
rect 922 16934 2510 17050
rect 17408 16940 17460 16992
rect 28632 16975 28643 16992
rect 28643 16975 28677 16992
rect 28677 16975 28684 16992
rect 28632 16940 28684 16975
rect 46126 16934 47714 17050
rect 27620 15444 27672 15496
rect 8116 15376 8168 15428
rect 3370 15054 4958 15170
rect 43678 15054 45266 15170
rect 8760 14832 8812 14884
rect 10416 14356 10468 14408
rect 14740 14356 14792 14408
rect 7932 13363 7984 13388
rect 7932 13336 7984 13363
rect 10692 13363 10744 13388
rect 10692 13336 10744 13363
rect 13728 13363 13780 13388
rect 13728 13336 13780 13363
rect 23572 14323 23595 14340
rect 23595 14323 23624 14340
rect 23572 14288 23624 14323
rect 39304 14861 39356 14884
rect 28632 14602 28650 14612
rect 28650 14602 28684 14612
rect 28632 14560 28684 14602
rect 28724 14432 28776 14476
rect 28724 14424 28756 14432
rect 28756 14424 28776 14432
rect 20076 13404 20128 13456
rect 39304 14832 39356 14861
rect 38200 13336 38252 13388
rect 922 13174 2510 13290
rect 17132 13200 17184 13252
rect 28632 13249 28684 13252
rect 28632 13215 28643 13249
rect 28643 13215 28677 13249
rect 28677 13215 28684 13249
rect 28632 13200 28684 13215
rect 46126 13174 47714 13290
rect 10692 12452 10744 12504
rect 8208 12384 8260 12436
rect 13728 11908 13780 11960
rect 19432 11908 19484 11960
rect 13912 11636 13964 11688
rect 20076 11636 20128 11688
rect 34060 11500 34112 11552
rect 35440 11500 35492 11552
rect 3370 11294 4958 11410
rect 43678 11294 45266 11410
rect 23664 11160 23716 11212
rect 7932 11024 7984 11076
rect 13912 11024 13964 11076
rect 20536 11092 20588 11144
rect 19432 11024 19484 11076
rect 9772 9596 9824 9648
rect 12532 9596 12584 9648
rect 13912 9596 13964 9648
rect 28816 10548 28868 10600
rect 31484 11092 31536 11144
rect 34060 11024 34112 11076
rect 28540 9596 28592 9648
rect 29460 10072 29512 10124
rect 32128 9596 32180 9648
rect 37004 10548 37056 10600
rect 34980 9596 35032 9648
rect 37648 9596 37700 9648
rect 922 9414 2510 9530
rect 17132 9460 17184 9512
rect 46126 9414 47714 9530
rect 32496 9324 32548 9376
rect 34980 9324 35032 9376
rect 37004 9324 37056 9376
rect 38108 9324 38160 9376
rect 14740 9188 14792 9240
rect 32128 9188 32180 9240
rect 12532 8916 12584 8968
rect 23204 8916 23256 8968
rect 3370 7534 4958 7650
rect 43678 7534 45266 7650
rect 8208 7352 8260 7404
rect 13912 7284 13964 7336
rect 17776 6808 17828 6860
rect 25596 7420 25648 7472
rect 23204 7284 23256 7336
rect 25688 6808 25740 6860
rect 28540 7284 28592 7336
rect 32496 7284 32548 7336
rect 37648 7420 37700 7472
rect 38200 7352 38252 7404
rect 8116 6468 8168 6520
rect 19524 6332 19576 6384
rect 20536 6381 20588 6384
rect 20536 6332 20588 6381
rect 23572 6332 23624 6384
rect 25596 6332 25648 6384
rect 28356 6060 28408 6112
rect 31484 6381 31536 6384
rect 31484 6332 31536 6381
rect 35348 6468 35400 6520
rect 38108 6468 38160 6520
rect 922 5654 2510 5770
rect 46126 5654 47714 5770
<< metal2 >>
rect 3348 41490 4980 41492
rect 3348 41374 3370 41490
rect 4958 41374 4980 41490
rect 3348 41372 4980 41374
rect 12438 41472 12494 41478
rect 12438 41420 12440 41472
rect 12492 41420 12494 41472
rect 12438 41398 12494 41420
rect 27448 41392 27476 47192
rect 12438 41333 12494 41342
rect 27356 41364 27476 41392
rect 43656 41490 45288 41492
rect 43656 41374 43678 41490
rect 45266 41374 45288 41490
rect 43656 41372 45288 41374
rect 27356 41206 27384 41364
rect 6798 41190 6998 41202
rect 6798 41134 6830 41190
rect 6886 41134 6910 41190
rect 6966 41134 6998 41190
rect 27344 41200 27396 41206
rect 27344 41142 27396 41148
rect 6798 41122 6998 41134
rect 38660 39840 38712 39846
rect 6820 39770 6980 39792
rect 38660 39782 38712 39788
rect 6820 39714 6872 39770
rect 6928 39714 6980 39770
rect 6820 39692 6980 39714
rect 9588 39704 9640 39710
rect 15016 39704 15068 39710
rect 9588 39646 9640 39652
rect 15014 39690 15016 39699
rect 27620 39704 27672 39710
rect 15068 39690 15070 39699
rect 900 39610 2532 39612
rect 900 39494 922 39610
rect 2510 39494 2532 39610
rect 900 39492 2532 39494
rect 3348 37730 4980 37732
rect 3348 37614 3370 37730
rect 4958 37614 4980 37730
rect 3348 37612 4980 37614
rect 5916 37430 6116 37442
rect 5916 37374 5948 37430
rect 6004 37374 6028 37430
rect 6084 37374 6116 37430
rect 5916 37362 6116 37374
rect 9600 36106 9628 39646
rect 15014 39625 15070 39634
rect 27618 39690 27620 39699
rect 27672 39690 27674 39699
rect 27618 39625 27674 39634
rect 15028 39613 15056 39625
rect 27632 39613 27660 39625
rect 12992 37664 13044 37670
rect 12990 37616 12992 37625
rect 16856 37664 16908 37670
rect 13044 37616 13046 37625
rect 12990 37551 13046 37560
rect 16854 37616 16856 37625
rect 27896 37664 27948 37670
rect 16908 37616 16910 37625
rect 16854 37551 16910 37560
rect 27894 37616 27896 37625
rect 27948 37616 27950 37625
rect 27894 37551 27950 37560
rect 13364 37430 13564 37442
rect 13364 37374 13396 37430
rect 13452 37374 13476 37430
rect 13532 37374 13564 37430
rect 13364 37362 13564 37374
rect 20812 37430 21012 37442
rect 20812 37374 20844 37430
rect 20900 37374 20924 37430
rect 20980 37374 21012 37430
rect 20812 37362 21012 37374
rect 30196 37188 30248 37194
rect 30196 37130 30248 37136
rect 26240 36168 26292 36174
rect 26240 36110 26292 36116
rect 9588 36100 9640 36106
rect 9588 36042 9640 36048
rect 5938 36010 6098 36032
rect 5938 35954 5990 36010
rect 6046 35954 6098 36010
rect 5938 35932 6098 35954
rect 900 35850 2532 35852
rect 900 35734 922 35850
rect 2510 35734 2532 35850
rect 900 35732 2532 35734
rect 3348 33970 4980 33972
rect 3348 33854 3370 33970
rect 4958 33854 4980 33970
rect 3348 33852 4980 33854
rect 6602 33670 6802 33682
rect 6602 33614 6634 33670
rect 6690 33614 6714 33670
rect 6770 33614 6802 33670
rect 6602 33602 6802 33614
rect 6624 32250 6784 32272
rect 6624 32194 6676 32250
rect 6732 32194 6784 32250
rect 6624 32172 6784 32194
rect 900 32090 2532 32092
rect 900 31974 922 32090
rect 2510 31974 2532 32090
rect 900 31972 2532 31974
rect 3348 30210 4980 30212
rect 3348 30094 3370 30210
rect 4958 30094 4980 30210
rect 3348 30092 4980 30094
rect 900 28330 2532 28332
rect 900 28214 922 28330
rect 2510 28214 2532 28330
rect 900 28212 2532 28214
rect 3348 26450 4980 26452
rect 3348 26334 3370 26450
rect 4958 26334 4980 26450
rect 3348 26332 4980 26334
rect 9600 26178 9628 36042
rect 13386 36010 13546 36032
rect 13386 35954 13438 36010
rect 13494 35954 13546 36010
rect 13386 35932 13546 35954
rect 20834 36010 20994 36032
rect 20834 35954 20886 36010
rect 20942 35954 20994 36010
rect 20834 35932 20994 35954
rect 9954 33924 10010 33930
rect 9954 33872 9956 33924
rect 10008 33872 10010 33924
rect 9954 33834 10010 33872
rect 9954 33769 10010 33778
rect 14186 32248 14242 32257
rect 14186 32183 14188 32192
rect 14240 32183 14242 32192
rect 14188 32166 14240 32172
rect 14200 28422 14228 32166
rect 18880 28688 18932 28694
rect 18880 28630 18932 28636
rect 18892 28597 18920 28630
rect 18878 28588 18934 28597
rect 18878 28523 18934 28532
rect 12532 28416 12584 28422
rect 12532 28358 12584 28364
rect 14188 28416 14240 28422
rect 14188 28358 14240 28364
rect 23388 28416 23440 28422
rect 23388 28358 23440 28364
rect 9588 26172 9640 26178
rect 9588 26114 9640 26120
rect 7104 25628 7156 25634
rect 7104 25570 7156 25576
rect 900 24570 2532 24572
rect 900 24454 922 24570
rect 2510 24454 2532 24570
rect 900 24452 2532 24454
rect 7116 23526 7144 25570
rect 12544 24682 12572 28358
rect 15422 26150 15622 26162
rect 15422 26094 15454 26150
rect 15510 26094 15534 26150
rect 15590 26094 15622 26150
rect 15422 26082 15622 26094
rect 23294 25050 23350 25059
rect 23400 25022 23428 28358
rect 26252 26246 26280 36110
rect 30208 35834 30236 37130
rect 31668 36508 31720 36514
rect 31668 36450 31720 36456
rect 30196 35828 30248 35834
rect 30196 35770 30248 35776
rect 26884 32292 26936 32298
rect 26884 32234 26936 32240
rect 26516 28552 26568 28558
rect 26516 28494 26568 28500
rect 26240 26240 26292 26246
rect 26240 26182 26292 26188
rect 23294 24985 23350 24994
rect 23388 25016 23440 25022
rect 23308 24886 23336 24985
rect 23388 24958 23440 24964
rect 23296 24880 23348 24886
rect 23296 24822 23348 24828
rect 15444 24730 15604 24752
rect 7196 24676 7248 24682
rect 7196 24618 7248 24624
rect 9680 24676 9732 24682
rect 9680 24618 9732 24624
rect 12532 24676 12584 24682
rect 15444 24674 15496 24730
rect 15552 24674 15604 24730
rect 15444 24652 15604 24674
rect 12532 24618 12584 24624
rect 7208 24274 7236 24618
rect 7196 24268 7248 24274
rect 7196 24210 7248 24216
rect 7104 23520 7156 23526
rect 7104 23462 7156 23468
rect 3348 22690 4980 22692
rect 3348 22574 3370 22690
rect 4958 22574 4980 22690
rect 3348 22572 4980 22574
rect 8300 22500 8352 22506
rect 8300 22442 8352 22448
rect 8312 20942 8340 22442
rect 8300 20936 8352 20942
rect 8300 20878 8352 20884
rect 900 20810 2532 20812
rect 900 20694 922 20810
rect 2510 20694 2532 20810
rect 900 20692 2532 20694
rect 3348 18930 4980 18932
rect 3348 18814 3370 18930
rect 4958 18814 4980 18930
rect 3348 18812 4980 18814
rect 9692 18358 9720 24618
rect 15474 24562 15530 24571
rect 15474 24497 15476 24506
rect 15528 24497 15530 24506
rect 15476 24482 15528 24488
rect 15488 24474 15516 24482
rect 13360 24268 13412 24274
rect 13360 24210 13412 24216
rect 13266 22610 13322 22619
rect 13266 22545 13322 22554
rect 13280 21010 13308 22545
rect 13268 21004 13320 21010
rect 13268 20946 13320 20952
rect 13372 18630 13400 24210
rect 13560 22390 13760 22402
rect 13560 22334 13592 22390
rect 13648 22334 13672 22390
rect 13728 22334 13760 22390
rect 13560 22322 13760 22334
rect 23308 22234 23336 24822
rect 23296 22228 23348 22234
rect 23296 22170 23348 22176
rect 20902 21634 20958 21643
rect 20902 21569 20904 21578
rect 20956 21569 20958 21578
rect 20904 21558 20956 21564
rect 20916 21546 20944 21558
rect 13582 20970 13742 20992
rect 13582 20914 13634 20970
rect 13690 20914 13742 20970
rect 13582 20892 13742 20914
rect 14094 20902 14150 20911
rect 14094 20837 14150 20846
rect 14108 20806 14136 20837
rect 14096 20800 14148 20806
rect 14096 20742 14148 20748
rect 20718 18950 20774 18959
rect 20718 18885 20774 18894
rect 16108 18630 16308 18642
rect 13360 18624 13412 18630
rect 13360 18566 13412 18572
rect 16108 18574 16140 18630
rect 16196 18574 16220 18630
rect 16276 18574 16308 18630
rect 16108 18562 16308 18574
rect 9680 18352 9732 18358
rect 9680 18294 9732 18300
rect 12532 18148 12584 18154
rect 12584 18108 13216 18136
rect 12532 18090 12584 18096
rect 13188 17678 13216 18108
rect 13176 17672 13228 17678
rect 13176 17614 13228 17620
rect 16130 17210 16290 17232
rect 8760 17196 8812 17202
rect 8760 17138 8812 17144
rect 16130 17154 16182 17210
rect 16238 17154 16290 17210
rect 900 17050 2532 17052
rect 900 16934 922 17050
rect 2510 16934 2532 17050
rect 900 16932 2532 16934
rect 8116 15428 8168 15434
rect 8116 15370 8168 15376
rect 3348 15170 4980 15172
rect 3348 15054 3370 15170
rect 4958 15054 4980 15170
rect 3348 15052 4980 15054
rect 7932 13388 7984 13394
rect 7932 13330 7984 13336
rect 900 13290 2532 13292
rect 900 13174 922 13290
rect 2510 13174 2532 13290
rect 900 13172 2532 13174
rect 3348 11410 4980 11412
rect 3348 11294 3370 11410
rect 4958 11294 4980 11410
rect 3348 11292 4980 11294
rect 7944 11082 7972 13330
rect 7932 11076 7984 11082
rect 7932 11018 7984 11024
rect 900 9530 2532 9532
rect 900 9414 922 9530
rect 2510 9414 2532 9530
rect 900 9412 2532 9414
rect 3348 7650 4980 7652
rect 3348 7534 3370 7650
rect 4958 7534 4980 7650
rect 3348 7532 4980 7534
rect 8128 6526 8156 15370
rect 8772 14890 8800 17138
rect 16130 17132 16290 17154
rect 17406 16998 17462 17007
rect 17406 16940 17408 16942
rect 17460 16940 17462 16942
rect 17406 16933 17462 16940
rect 17420 16910 17448 16933
rect 20732 16397 20760 18885
rect 23400 17338 23428 24958
rect 26252 22624 26280 26182
rect 26252 22596 26464 22624
rect 26436 22506 26464 22596
rect 26424 22500 26476 22506
rect 26424 22442 26476 22448
rect 26528 21282 26556 28494
rect 26516 21276 26568 21282
rect 26516 21218 26568 21224
rect 23388 17332 23440 17338
rect 23388 17274 23440 17280
rect 26528 17202 26556 21218
rect 26896 21146 26924 32234
rect 31680 25770 31708 36450
rect 31668 25764 31720 25770
rect 31668 25706 31720 25712
rect 28632 25220 28684 25226
rect 28632 25162 28684 25168
rect 27620 24880 27672 24886
rect 27620 24822 27672 24828
rect 26884 21140 26936 21146
rect 26884 21082 26936 21088
rect 26516 17196 26568 17202
rect 26516 17138 26568 17144
rect 20718 16388 20774 16397
rect 20718 16323 20774 16332
rect 27632 15502 27660 24822
rect 28644 22030 28672 25162
rect 30104 23520 30156 23526
rect 30104 23462 30156 23468
rect 28632 22024 28684 22030
rect 28632 21966 28684 21972
rect 28724 21412 28776 21418
rect 28724 21354 28776 21360
rect 28632 18420 28684 18426
rect 28632 18362 28684 18368
rect 28644 16998 28672 18362
rect 28736 18222 28764 21354
rect 30116 21214 30144 23462
rect 38672 22438 38700 39782
rect 46104 39610 47736 39612
rect 46104 39494 46126 39610
rect 47714 39494 47736 39610
rect 46104 39492 47736 39494
rect 43656 37730 45288 37732
rect 43656 37614 43678 37730
rect 45266 37614 45288 37730
rect 43656 37612 45288 37614
rect 39948 36780 40000 36786
rect 39948 36722 40000 36728
rect 39960 29152 39988 36722
rect 46104 35850 47736 35852
rect 46104 35734 46126 35850
rect 47714 35734 47736 35850
rect 46104 35732 47736 35734
rect 43656 33970 45288 33972
rect 43656 33854 43678 33970
rect 45266 33854 45288 33970
rect 43656 33852 45288 33854
rect 40040 32428 40092 32434
rect 40040 32370 40092 32376
rect 40052 29918 40080 32370
rect 46104 32090 47736 32092
rect 46104 31974 46126 32090
rect 47714 31974 47736 32090
rect 46104 31972 47736 31974
rect 43656 30210 45288 30212
rect 43656 30094 43678 30210
rect 45266 30094 45288 30210
rect 43656 30092 45288 30094
rect 40040 29912 40092 29918
rect 40040 29854 40092 29860
rect 39316 29124 39988 29152
rect 39316 28966 39344 29124
rect 39304 28960 39356 28966
rect 39304 28902 39356 28908
rect 40040 28484 40092 28490
rect 40040 28426 40092 28432
rect 39396 25696 39448 25702
rect 39396 25638 39448 25644
rect 39408 24954 39436 25638
rect 39396 24948 39448 24954
rect 40052 24936 40080 28426
rect 46104 28330 47736 28332
rect 46104 28214 46126 28330
rect 47714 28214 47736 28330
rect 46104 28212 47736 28214
rect 43656 26450 45288 26452
rect 43656 26334 43678 26450
rect 45266 26334 45288 26450
rect 43656 26332 45288 26334
rect 39396 24890 39448 24896
rect 39500 24908 40080 24936
rect 38660 22432 38712 22438
rect 38660 22374 38712 22380
rect 30564 22160 30616 22166
rect 30564 22102 30616 22108
rect 30104 21208 30156 21214
rect 30104 21150 30156 21156
rect 30576 20806 30604 22102
rect 30564 20800 30616 20806
rect 30564 20742 30616 20748
rect 39500 18630 39528 24908
rect 46104 24570 47736 24572
rect 46104 24454 46126 24570
rect 47714 24454 47736 24570
rect 46104 24452 47736 24454
rect 43656 22690 45288 22692
rect 43656 22574 43678 22690
rect 45266 22574 45288 22690
rect 43656 22572 45288 22574
rect 46104 20810 47736 20812
rect 46104 20694 46126 20810
rect 47714 20694 47736 20810
rect 46104 20692 47736 20694
rect 43656 18930 45288 18932
rect 43656 18814 43678 18930
rect 45266 18814 45288 18930
rect 43656 18812 45288 18814
rect 39488 18624 39540 18630
rect 39488 18566 39540 18572
rect 28724 18216 28776 18222
rect 28724 18158 28776 18164
rect 28724 17672 28776 17678
rect 28724 17614 28776 17620
rect 28632 16992 28684 16998
rect 28632 16934 28684 16940
rect 27620 15496 27672 15502
rect 27620 15438 27672 15444
rect 8760 14884 8812 14890
rect 8760 14826 8812 14832
rect 16108 14870 16308 14882
rect 16108 14814 16140 14870
rect 16196 14814 16220 14870
rect 16276 14814 16308 14870
rect 16108 14802 16308 14814
rect 28632 14612 28684 14618
rect 28632 14554 28684 14560
rect 10416 14408 10468 14414
rect 10416 14350 10468 14356
rect 14740 14408 14792 14414
rect 14740 14350 14792 14356
rect 10428 14192 10456 14350
rect 9784 14164 10456 14192
rect 8208 12436 8260 12442
rect 8208 12378 8260 12384
rect 8220 7410 8248 12378
rect 9784 9654 9812 14164
rect 10692 13388 10744 13394
rect 10692 13330 10744 13336
rect 13728 13388 13780 13394
rect 13728 13330 13780 13336
rect 10704 12510 10732 13330
rect 10692 12504 10744 12510
rect 10692 12446 10744 12452
rect 13740 11966 13768 13330
rect 13728 11960 13780 11966
rect 13728 11902 13780 11908
rect 13912 11688 13964 11694
rect 13912 11630 13964 11636
rect 13924 11082 13952 11630
rect 13912 11076 13964 11082
rect 13912 11018 13964 11024
rect 9772 9648 9824 9654
rect 9772 9590 9824 9596
rect 12532 9648 12584 9654
rect 12532 9590 12584 9596
rect 13912 9648 13964 9654
rect 13912 9590 13964 9596
rect 12544 8974 12572 9590
rect 12532 8968 12584 8974
rect 12532 8910 12584 8916
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 13924 7342 13952 9590
rect 14752 9246 14780 14350
rect 23572 14340 23624 14346
rect 23572 14282 23624 14288
rect 16130 13450 16290 13472
rect 16130 13394 16182 13450
rect 16238 13394 16290 13450
rect 17130 13460 17186 13469
rect 17130 13395 17186 13404
rect 20076 13456 20128 13462
rect 20076 13398 20128 13404
rect 16130 13372 16290 13394
rect 17144 13258 17172 13395
rect 17132 13252 17184 13258
rect 17132 13194 17184 13200
rect 19432 11960 19484 11966
rect 19432 11902 19484 11908
rect 16108 11110 16308 11122
rect 16108 11054 16140 11110
rect 16196 11054 16220 11110
rect 16276 11054 16308 11110
rect 19444 11082 19472 11902
rect 20088 11694 20116 13398
rect 20076 11688 20128 11694
rect 20076 11630 20128 11636
rect 20536 11144 20588 11150
rect 20536 11086 20588 11092
rect 16108 11042 16308 11054
rect 19432 11076 19484 11082
rect 19432 11018 19484 11024
rect 16130 9690 16290 9712
rect 16130 9634 16182 9690
rect 16238 9634 16290 9690
rect 16130 9612 16290 9634
rect 17130 9678 17186 9687
rect 17130 9613 17186 9622
rect 17144 9518 17172 9613
rect 17132 9512 17184 9518
rect 17132 9454 17184 9460
rect 14740 9240 14792 9246
rect 14740 9182 14792 9188
rect 13912 7336 13964 7342
rect 13912 7278 13964 7284
rect 17776 6860 17828 6866
rect 17776 6802 17828 6808
rect 8116 6520 8168 6526
rect 8116 6462 8168 6468
rect 17788 6149 17816 6802
rect 19522 6506 19578 6515
rect 19522 6441 19578 6450
rect 19536 6390 19564 6441
rect 20548 6390 20576 11086
rect 23204 8968 23256 8974
rect 23204 8910 23256 8916
rect 23216 7342 23244 8910
rect 23204 7336 23256 7342
rect 23204 7278 23256 7284
rect 23584 6390 23612 14282
rect 28644 13258 28672 14554
rect 28736 14482 28764 17614
rect 39304 17196 39356 17202
rect 39304 17138 39356 17144
rect 39316 14890 39344 17138
rect 46104 17050 47736 17052
rect 46104 16934 46126 17050
rect 47714 16934 47736 17050
rect 46104 16932 47736 16934
rect 43656 15170 45288 15172
rect 43656 15054 43678 15170
rect 45266 15054 45288 15170
rect 43656 15052 45288 15054
rect 39304 14884 39356 14890
rect 39304 14826 39356 14832
rect 28724 14476 28776 14482
rect 28724 14418 28776 14424
rect 38200 13388 38252 13394
rect 38200 13330 38252 13336
rect 28632 13252 28684 13258
rect 28632 13194 28684 13200
rect 34060 11552 34112 11558
rect 34060 11494 34112 11500
rect 35440 11552 35492 11558
rect 35440 11494 35492 11500
rect 23662 11212 23718 11218
rect 23662 11160 23664 11212
rect 23716 11160 23718 11212
rect 23662 11142 23718 11160
rect 31484 11144 31536 11150
rect 31484 11086 31536 11092
rect 23662 11077 23718 11086
rect 28816 10600 28868 10606
rect 28816 10542 28868 10548
rect 28828 10112 28856 10542
rect 29460 10124 29512 10130
rect 28828 10084 29460 10112
rect 29460 10066 29512 10072
rect 28540 9648 28592 9654
rect 28540 9590 28592 9596
rect 25596 7472 25648 7478
rect 25596 7414 25648 7420
rect 25608 6390 25636 7414
rect 28552 7342 28580 9590
rect 28540 7336 28592 7342
rect 28540 7278 28592 7284
rect 25688 6860 25740 6866
rect 25688 6802 25740 6808
rect 25700 6515 25728 6802
rect 25686 6506 25742 6515
rect 25686 6441 25742 6450
rect 31496 6390 31524 11086
rect 34072 11082 34100 11494
rect 35452 11336 35480 11494
rect 35360 11308 35480 11336
rect 34060 11076 34112 11082
rect 34060 11018 34112 11024
rect 32128 9648 32180 9654
rect 32128 9590 32180 9596
rect 34980 9648 35032 9654
rect 34980 9590 35032 9596
rect 32140 9246 32168 9590
rect 34992 9382 35020 9590
rect 32496 9376 32548 9382
rect 32496 9318 32548 9324
rect 34980 9376 35032 9382
rect 34980 9318 35032 9324
rect 32128 9240 32180 9246
rect 32128 9182 32180 9188
rect 32508 7342 32536 9318
rect 32496 7336 32548 7342
rect 32496 7278 32548 7284
rect 35360 6526 35388 11308
rect 37004 10600 37056 10606
rect 37004 10542 37056 10548
rect 37016 9382 37044 10542
rect 37648 9648 37700 9654
rect 37648 9590 37700 9596
rect 37004 9376 37056 9382
rect 37004 9318 37056 9324
rect 37660 7478 37688 9590
rect 38108 9376 38160 9382
rect 38108 9318 38160 9324
rect 37648 7472 37700 7478
rect 37648 7414 37700 7420
rect 38120 6526 38148 9318
rect 38212 7410 38240 13330
rect 46104 13290 47736 13292
rect 46104 13174 46126 13290
rect 47714 13174 47736 13290
rect 46104 13172 47736 13174
rect 43656 11410 45288 11412
rect 43656 11294 43678 11410
rect 45266 11294 45288 11410
rect 43656 11292 45288 11294
rect 46104 9530 47736 9532
rect 46104 9414 46126 9530
rect 47714 9414 47736 9530
rect 46104 9412 47736 9414
rect 43656 7650 45288 7652
rect 43656 7534 43678 7650
rect 45266 7534 45288 7650
rect 43656 7532 45288 7534
rect 38200 7404 38252 7410
rect 38200 7346 38252 7352
rect 35348 6520 35400 6526
rect 35348 6462 35400 6468
rect 38108 6520 38160 6526
rect 38108 6462 38160 6468
rect 19524 6384 19576 6390
rect 19524 6326 19576 6332
rect 20536 6384 20588 6390
rect 20536 6326 20588 6332
rect 23572 6384 23624 6390
rect 23572 6326 23624 6332
rect 25596 6384 25648 6390
rect 25596 6326 25648 6332
rect 31484 6384 31536 6390
rect 31484 6326 31536 6332
rect 17774 6140 17830 6149
rect 17774 6075 17830 6084
rect 28354 6140 28410 6149
rect 28354 6075 28356 6084
rect 28408 6075 28410 6084
rect 28356 6054 28408 6060
rect 28368 6052 28396 6054
rect 900 5770 2532 5772
rect 900 5654 922 5770
rect 2510 5654 2532 5770
rect 900 5652 2532 5654
rect 46104 5770 47736 5772
rect 46104 5654 46126 5770
rect 47714 5654 47736 5770
rect 46104 5652 47736 5654
<< via2 >>
rect 3376 41404 3432 41460
rect 3456 41404 3512 41460
rect 3536 41404 3592 41460
rect 3616 41404 3672 41460
rect 3696 41404 3752 41460
rect 3776 41404 3832 41460
rect 3856 41404 3912 41460
rect 3936 41404 3992 41460
rect 4016 41404 4072 41460
rect 4096 41404 4152 41460
rect 4176 41404 4232 41460
rect 4256 41404 4312 41460
rect 4336 41404 4392 41460
rect 4416 41404 4472 41460
rect 4496 41404 4552 41460
rect 4576 41404 4632 41460
rect 4656 41404 4712 41460
rect 4736 41404 4792 41460
rect 4816 41404 4872 41460
rect 4896 41404 4952 41460
rect 12438 41342 12494 41398
rect 43684 41404 43740 41460
rect 43764 41404 43820 41460
rect 43844 41404 43900 41460
rect 43924 41404 43980 41460
rect 44004 41404 44060 41460
rect 44084 41404 44140 41460
rect 44164 41404 44220 41460
rect 44244 41404 44300 41460
rect 44324 41404 44380 41460
rect 44404 41404 44460 41460
rect 44484 41404 44540 41460
rect 44564 41404 44620 41460
rect 44644 41404 44700 41460
rect 44724 41404 44780 41460
rect 44804 41404 44860 41460
rect 44884 41404 44940 41460
rect 44964 41404 45020 41460
rect 45044 41404 45100 41460
rect 45124 41404 45180 41460
rect 45204 41404 45260 41460
rect 6830 41134 6886 41190
rect 6910 41134 6966 41190
rect 6872 39714 6928 39770
rect 15014 39652 15016 39690
rect 15016 39652 15068 39690
rect 15068 39652 15070 39690
rect 928 39524 984 39580
rect 1008 39524 1064 39580
rect 1088 39524 1144 39580
rect 1168 39524 1224 39580
rect 1248 39524 1304 39580
rect 1328 39524 1384 39580
rect 1408 39524 1464 39580
rect 1488 39524 1544 39580
rect 1568 39524 1624 39580
rect 1648 39524 1704 39580
rect 1728 39524 1784 39580
rect 1808 39524 1864 39580
rect 1888 39524 1944 39580
rect 1968 39524 2024 39580
rect 2048 39524 2104 39580
rect 2128 39524 2184 39580
rect 2208 39524 2264 39580
rect 2288 39524 2344 39580
rect 2368 39524 2424 39580
rect 2448 39524 2504 39580
rect 3376 37644 3432 37700
rect 3456 37644 3512 37700
rect 3536 37644 3592 37700
rect 3616 37644 3672 37700
rect 3696 37644 3752 37700
rect 3776 37644 3832 37700
rect 3856 37644 3912 37700
rect 3936 37644 3992 37700
rect 4016 37644 4072 37700
rect 4096 37644 4152 37700
rect 4176 37644 4232 37700
rect 4256 37644 4312 37700
rect 4336 37644 4392 37700
rect 4416 37644 4472 37700
rect 4496 37644 4552 37700
rect 4576 37644 4632 37700
rect 4656 37644 4712 37700
rect 4736 37644 4792 37700
rect 4816 37644 4872 37700
rect 4896 37644 4952 37700
rect 5948 37374 6004 37430
rect 6028 37374 6084 37430
rect 15014 39634 15070 39652
rect 27618 39652 27620 39690
rect 27620 39652 27672 39690
rect 27672 39652 27674 39690
rect 27618 39634 27674 39652
rect 12990 37612 12992 37616
rect 12992 37612 13044 37616
rect 13044 37612 13046 37616
rect 12990 37560 13046 37612
rect 16854 37612 16856 37616
rect 16856 37612 16908 37616
rect 16908 37612 16910 37616
rect 16854 37560 16910 37612
rect 27894 37612 27896 37616
rect 27896 37612 27948 37616
rect 27948 37612 27950 37616
rect 27894 37560 27950 37612
rect 13396 37374 13452 37430
rect 13476 37374 13532 37430
rect 20844 37374 20900 37430
rect 20924 37374 20980 37430
rect 5990 35954 6046 36010
rect 928 35764 984 35820
rect 1008 35764 1064 35820
rect 1088 35764 1144 35820
rect 1168 35764 1224 35820
rect 1248 35764 1304 35820
rect 1328 35764 1384 35820
rect 1408 35764 1464 35820
rect 1488 35764 1544 35820
rect 1568 35764 1624 35820
rect 1648 35764 1704 35820
rect 1728 35764 1784 35820
rect 1808 35764 1864 35820
rect 1888 35764 1944 35820
rect 1968 35764 2024 35820
rect 2048 35764 2104 35820
rect 2128 35764 2184 35820
rect 2208 35764 2264 35820
rect 2288 35764 2344 35820
rect 2368 35764 2424 35820
rect 2448 35764 2504 35820
rect 3376 33884 3432 33940
rect 3456 33884 3512 33940
rect 3536 33884 3592 33940
rect 3616 33884 3672 33940
rect 3696 33884 3752 33940
rect 3776 33884 3832 33940
rect 3856 33884 3912 33940
rect 3936 33884 3992 33940
rect 4016 33884 4072 33940
rect 4096 33884 4152 33940
rect 4176 33884 4232 33940
rect 4256 33884 4312 33940
rect 4336 33884 4392 33940
rect 4416 33884 4472 33940
rect 4496 33884 4552 33940
rect 4576 33884 4632 33940
rect 4656 33884 4712 33940
rect 4736 33884 4792 33940
rect 4816 33884 4872 33940
rect 4896 33884 4952 33940
rect 6634 33614 6690 33670
rect 6714 33614 6770 33670
rect 6676 32194 6732 32250
rect 928 32004 984 32060
rect 1008 32004 1064 32060
rect 1088 32004 1144 32060
rect 1168 32004 1224 32060
rect 1248 32004 1304 32060
rect 1328 32004 1384 32060
rect 1408 32004 1464 32060
rect 1488 32004 1544 32060
rect 1568 32004 1624 32060
rect 1648 32004 1704 32060
rect 1728 32004 1784 32060
rect 1808 32004 1864 32060
rect 1888 32004 1944 32060
rect 1968 32004 2024 32060
rect 2048 32004 2104 32060
rect 2128 32004 2184 32060
rect 2208 32004 2264 32060
rect 2288 32004 2344 32060
rect 2368 32004 2424 32060
rect 2448 32004 2504 32060
rect 3376 30124 3432 30180
rect 3456 30124 3512 30180
rect 3536 30124 3592 30180
rect 3616 30124 3672 30180
rect 3696 30124 3752 30180
rect 3776 30124 3832 30180
rect 3856 30124 3912 30180
rect 3936 30124 3992 30180
rect 4016 30124 4072 30180
rect 4096 30124 4152 30180
rect 4176 30124 4232 30180
rect 4256 30124 4312 30180
rect 4336 30124 4392 30180
rect 4416 30124 4472 30180
rect 4496 30124 4552 30180
rect 4576 30124 4632 30180
rect 4656 30124 4712 30180
rect 4736 30124 4792 30180
rect 4816 30124 4872 30180
rect 4896 30124 4952 30180
rect 928 28244 984 28300
rect 1008 28244 1064 28300
rect 1088 28244 1144 28300
rect 1168 28244 1224 28300
rect 1248 28244 1304 28300
rect 1328 28244 1384 28300
rect 1408 28244 1464 28300
rect 1488 28244 1544 28300
rect 1568 28244 1624 28300
rect 1648 28244 1704 28300
rect 1728 28244 1784 28300
rect 1808 28244 1864 28300
rect 1888 28244 1944 28300
rect 1968 28244 2024 28300
rect 2048 28244 2104 28300
rect 2128 28244 2184 28300
rect 2208 28244 2264 28300
rect 2288 28244 2344 28300
rect 2368 28244 2424 28300
rect 2448 28244 2504 28300
rect 3376 26364 3432 26420
rect 3456 26364 3512 26420
rect 3536 26364 3592 26420
rect 3616 26364 3672 26420
rect 3696 26364 3752 26420
rect 3776 26364 3832 26420
rect 3856 26364 3912 26420
rect 3936 26364 3992 26420
rect 4016 26364 4072 26420
rect 4096 26364 4152 26420
rect 4176 26364 4232 26420
rect 4256 26364 4312 26420
rect 4336 26364 4392 26420
rect 4416 26364 4472 26420
rect 4496 26364 4552 26420
rect 4576 26364 4632 26420
rect 4656 26364 4712 26420
rect 4736 26364 4792 26420
rect 4816 26364 4872 26420
rect 4896 26364 4952 26420
rect 13438 35954 13494 36010
rect 20886 35954 20942 36010
rect 9954 33778 10010 33834
rect 14186 32224 14242 32248
rect 14186 32192 14188 32224
rect 14188 32192 14240 32224
rect 14240 32192 14242 32224
rect 18878 28532 18934 28588
rect 928 24484 984 24540
rect 1008 24484 1064 24540
rect 1088 24484 1144 24540
rect 1168 24484 1224 24540
rect 1248 24484 1304 24540
rect 1328 24484 1384 24540
rect 1408 24484 1464 24540
rect 1488 24484 1544 24540
rect 1568 24484 1624 24540
rect 1648 24484 1704 24540
rect 1728 24484 1784 24540
rect 1808 24484 1864 24540
rect 1888 24484 1944 24540
rect 1968 24484 2024 24540
rect 2048 24484 2104 24540
rect 2128 24484 2184 24540
rect 2208 24484 2264 24540
rect 2288 24484 2344 24540
rect 2368 24484 2424 24540
rect 2448 24484 2504 24540
rect 15454 26094 15510 26150
rect 15534 26094 15590 26150
rect 23294 24994 23350 25050
rect 15496 24674 15552 24730
rect 3376 22604 3432 22660
rect 3456 22604 3512 22660
rect 3536 22604 3592 22660
rect 3616 22604 3672 22660
rect 3696 22604 3752 22660
rect 3776 22604 3832 22660
rect 3856 22604 3912 22660
rect 3936 22604 3992 22660
rect 4016 22604 4072 22660
rect 4096 22604 4152 22660
rect 4176 22604 4232 22660
rect 4256 22604 4312 22660
rect 4336 22604 4392 22660
rect 4416 22604 4472 22660
rect 4496 22604 4552 22660
rect 4576 22604 4632 22660
rect 4656 22604 4712 22660
rect 4736 22604 4792 22660
rect 4816 22604 4872 22660
rect 4896 22604 4952 22660
rect 928 20724 984 20780
rect 1008 20724 1064 20780
rect 1088 20724 1144 20780
rect 1168 20724 1224 20780
rect 1248 20724 1304 20780
rect 1328 20724 1384 20780
rect 1408 20724 1464 20780
rect 1488 20724 1544 20780
rect 1568 20724 1624 20780
rect 1648 20724 1704 20780
rect 1728 20724 1784 20780
rect 1808 20724 1864 20780
rect 1888 20724 1944 20780
rect 1968 20724 2024 20780
rect 2048 20724 2104 20780
rect 2128 20724 2184 20780
rect 2208 20724 2264 20780
rect 2288 20724 2344 20780
rect 2368 20724 2424 20780
rect 2448 20724 2504 20780
rect 3376 18844 3432 18900
rect 3456 18844 3512 18900
rect 3536 18844 3592 18900
rect 3616 18844 3672 18900
rect 3696 18844 3752 18900
rect 3776 18844 3832 18900
rect 3856 18844 3912 18900
rect 3936 18844 3992 18900
rect 4016 18844 4072 18900
rect 4096 18844 4152 18900
rect 4176 18844 4232 18900
rect 4256 18844 4312 18900
rect 4336 18844 4392 18900
rect 4416 18844 4472 18900
rect 4496 18844 4552 18900
rect 4576 18844 4632 18900
rect 4656 18844 4712 18900
rect 4736 18844 4792 18900
rect 4816 18844 4872 18900
rect 4896 18844 4952 18900
rect 15474 24540 15530 24562
rect 15474 24506 15476 24540
rect 15476 24506 15528 24540
rect 15528 24506 15530 24540
rect 13266 22554 13322 22610
rect 13592 22334 13648 22390
rect 13672 22334 13728 22390
rect 20902 21616 20958 21634
rect 20902 21578 20904 21616
rect 20904 21578 20956 21616
rect 20956 21578 20958 21616
rect 13634 20914 13690 20970
rect 14094 20846 14150 20902
rect 20718 18894 20774 18950
rect 16140 18574 16196 18630
rect 16220 18574 16276 18630
rect 16182 17154 16238 17210
rect 928 16964 984 17020
rect 1008 16964 1064 17020
rect 1088 16964 1144 17020
rect 1168 16964 1224 17020
rect 1248 16964 1304 17020
rect 1328 16964 1384 17020
rect 1408 16964 1464 17020
rect 1488 16964 1544 17020
rect 1568 16964 1624 17020
rect 1648 16964 1704 17020
rect 1728 16964 1784 17020
rect 1808 16964 1864 17020
rect 1888 16964 1944 17020
rect 1968 16964 2024 17020
rect 2048 16964 2104 17020
rect 2128 16964 2184 17020
rect 2208 16964 2264 17020
rect 2288 16964 2344 17020
rect 2368 16964 2424 17020
rect 2448 16964 2504 17020
rect 3376 15084 3432 15140
rect 3456 15084 3512 15140
rect 3536 15084 3592 15140
rect 3616 15084 3672 15140
rect 3696 15084 3752 15140
rect 3776 15084 3832 15140
rect 3856 15084 3912 15140
rect 3936 15084 3992 15140
rect 4016 15084 4072 15140
rect 4096 15084 4152 15140
rect 4176 15084 4232 15140
rect 4256 15084 4312 15140
rect 4336 15084 4392 15140
rect 4416 15084 4472 15140
rect 4496 15084 4552 15140
rect 4576 15084 4632 15140
rect 4656 15084 4712 15140
rect 4736 15084 4792 15140
rect 4816 15084 4872 15140
rect 4896 15084 4952 15140
rect 928 13204 984 13260
rect 1008 13204 1064 13260
rect 1088 13204 1144 13260
rect 1168 13204 1224 13260
rect 1248 13204 1304 13260
rect 1328 13204 1384 13260
rect 1408 13204 1464 13260
rect 1488 13204 1544 13260
rect 1568 13204 1624 13260
rect 1648 13204 1704 13260
rect 1728 13204 1784 13260
rect 1808 13204 1864 13260
rect 1888 13204 1944 13260
rect 1968 13204 2024 13260
rect 2048 13204 2104 13260
rect 2128 13204 2184 13260
rect 2208 13204 2264 13260
rect 2288 13204 2344 13260
rect 2368 13204 2424 13260
rect 2448 13204 2504 13260
rect 3376 11324 3432 11380
rect 3456 11324 3512 11380
rect 3536 11324 3592 11380
rect 3616 11324 3672 11380
rect 3696 11324 3752 11380
rect 3776 11324 3832 11380
rect 3856 11324 3912 11380
rect 3936 11324 3992 11380
rect 4016 11324 4072 11380
rect 4096 11324 4152 11380
rect 4176 11324 4232 11380
rect 4256 11324 4312 11380
rect 4336 11324 4392 11380
rect 4416 11324 4472 11380
rect 4496 11324 4552 11380
rect 4576 11324 4632 11380
rect 4656 11324 4712 11380
rect 4736 11324 4792 11380
rect 4816 11324 4872 11380
rect 4896 11324 4952 11380
rect 928 9444 984 9500
rect 1008 9444 1064 9500
rect 1088 9444 1144 9500
rect 1168 9444 1224 9500
rect 1248 9444 1304 9500
rect 1328 9444 1384 9500
rect 1408 9444 1464 9500
rect 1488 9444 1544 9500
rect 1568 9444 1624 9500
rect 1648 9444 1704 9500
rect 1728 9444 1784 9500
rect 1808 9444 1864 9500
rect 1888 9444 1944 9500
rect 1968 9444 2024 9500
rect 2048 9444 2104 9500
rect 2128 9444 2184 9500
rect 2208 9444 2264 9500
rect 2288 9444 2344 9500
rect 2368 9444 2424 9500
rect 2448 9444 2504 9500
rect 3376 7564 3432 7620
rect 3456 7564 3512 7620
rect 3536 7564 3592 7620
rect 3616 7564 3672 7620
rect 3696 7564 3752 7620
rect 3776 7564 3832 7620
rect 3856 7564 3912 7620
rect 3936 7564 3992 7620
rect 4016 7564 4072 7620
rect 4096 7564 4152 7620
rect 4176 7564 4232 7620
rect 4256 7564 4312 7620
rect 4336 7564 4392 7620
rect 4416 7564 4472 7620
rect 4496 7564 4552 7620
rect 4576 7564 4632 7620
rect 4656 7564 4712 7620
rect 4736 7564 4792 7620
rect 4816 7564 4872 7620
rect 4896 7564 4952 7620
rect 17406 16992 17462 16998
rect 17406 16942 17408 16992
rect 17408 16942 17460 16992
rect 17460 16942 17462 16992
rect 20718 16332 20774 16388
rect 46132 39524 46188 39580
rect 46212 39524 46268 39580
rect 46292 39524 46348 39580
rect 46372 39524 46428 39580
rect 46452 39524 46508 39580
rect 46532 39524 46588 39580
rect 46612 39524 46668 39580
rect 46692 39524 46748 39580
rect 46772 39524 46828 39580
rect 46852 39524 46908 39580
rect 46932 39524 46988 39580
rect 47012 39524 47068 39580
rect 47092 39524 47148 39580
rect 47172 39524 47228 39580
rect 47252 39524 47308 39580
rect 47332 39524 47388 39580
rect 47412 39524 47468 39580
rect 47492 39524 47548 39580
rect 47572 39524 47628 39580
rect 47652 39524 47708 39580
rect 43684 37644 43740 37700
rect 43764 37644 43820 37700
rect 43844 37644 43900 37700
rect 43924 37644 43980 37700
rect 44004 37644 44060 37700
rect 44084 37644 44140 37700
rect 44164 37644 44220 37700
rect 44244 37644 44300 37700
rect 44324 37644 44380 37700
rect 44404 37644 44460 37700
rect 44484 37644 44540 37700
rect 44564 37644 44620 37700
rect 44644 37644 44700 37700
rect 44724 37644 44780 37700
rect 44804 37644 44860 37700
rect 44884 37644 44940 37700
rect 44964 37644 45020 37700
rect 45044 37644 45100 37700
rect 45124 37644 45180 37700
rect 45204 37644 45260 37700
rect 46132 35764 46188 35820
rect 46212 35764 46268 35820
rect 46292 35764 46348 35820
rect 46372 35764 46428 35820
rect 46452 35764 46508 35820
rect 46532 35764 46588 35820
rect 46612 35764 46668 35820
rect 46692 35764 46748 35820
rect 46772 35764 46828 35820
rect 46852 35764 46908 35820
rect 46932 35764 46988 35820
rect 47012 35764 47068 35820
rect 47092 35764 47148 35820
rect 47172 35764 47228 35820
rect 47252 35764 47308 35820
rect 47332 35764 47388 35820
rect 47412 35764 47468 35820
rect 47492 35764 47548 35820
rect 47572 35764 47628 35820
rect 47652 35764 47708 35820
rect 43684 33884 43740 33940
rect 43764 33884 43820 33940
rect 43844 33884 43900 33940
rect 43924 33884 43980 33940
rect 44004 33884 44060 33940
rect 44084 33884 44140 33940
rect 44164 33884 44220 33940
rect 44244 33884 44300 33940
rect 44324 33884 44380 33940
rect 44404 33884 44460 33940
rect 44484 33884 44540 33940
rect 44564 33884 44620 33940
rect 44644 33884 44700 33940
rect 44724 33884 44780 33940
rect 44804 33884 44860 33940
rect 44884 33884 44940 33940
rect 44964 33884 45020 33940
rect 45044 33884 45100 33940
rect 45124 33884 45180 33940
rect 45204 33884 45260 33940
rect 46132 32004 46188 32060
rect 46212 32004 46268 32060
rect 46292 32004 46348 32060
rect 46372 32004 46428 32060
rect 46452 32004 46508 32060
rect 46532 32004 46588 32060
rect 46612 32004 46668 32060
rect 46692 32004 46748 32060
rect 46772 32004 46828 32060
rect 46852 32004 46908 32060
rect 46932 32004 46988 32060
rect 47012 32004 47068 32060
rect 47092 32004 47148 32060
rect 47172 32004 47228 32060
rect 47252 32004 47308 32060
rect 47332 32004 47388 32060
rect 47412 32004 47468 32060
rect 47492 32004 47548 32060
rect 47572 32004 47628 32060
rect 47652 32004 47708 32060
rect 43684 30124 43740 30180
rect 43764 30124 43820 30180
rect 43844 30124 43900 30180
rect 43924 30124 43980 30180
rect 44004 30124 44060 30180
rect 44084 30124 44140 30180
rect 44164 30124 44220 30180
rect 44244 30124 44300 30180
rect 44324 30124 44380 30180
rect 44404 30124 44460 30180
rect 44484 30124 44540 30180
rect 44564 30124 44620 30180
rect 44644 30124 44700 30180
rect 44724 30124 44780 30180
rect 44804 30124 44860 30180
rect 44884 30124 44940 30180
rect 44964 30124 45020 30180
rect 45044 30124 45100 30180
rect 45124 30124 45180 30180
rect 45204 30124 45260 30180
rect 46132 28244 46188 28300
rect 46212 28244 46268 28300
rect 46292 28244 46348 28300
rect 46372 28244 46428 28300
rect 46452 28244 46508 28300
rect 46532 28244 46588 28300
rect 46612 28244 46668 28300
rect 46692 28244 46748 28300
rect 46772 28244 46828 28300
rect 46852 28244 46908 28300
rect 46932 28244 46988 28300
rect 47012 28244 47068 28300
rect 47092 28244 47148 28300
rect 47172 28244 47228 28300
rect 47252 28244 47308 28300
rect 47332 28244 47388 28300
rect 47412 28244 47468 28300
rect 47492 28244 47548 28300
rect 47572 28244 47628 28300
rect 47652 28244 47708 28300
rect 43684 26364 43740 26420
rect 43764 26364 43820 26420
rect 43844 26364 43900 26420
rect 43924 26364 43980 26420
rect 44004 26364 44060 26420
rect 44084 26364 44140 26420
rect 44164 26364 44220 26420
rect 44244 26364 44300 26420
rect 44324 26364 44380 26420
rect 44404 26364 44460 26420
rect 44484 26364 44540 26420
rect 44564 26364 44620 26420
rect 44644 26364 44700 26420
rect 44724 26364 44780 26420
rect 44804 26364 44860 26420
rect 44884 26364 44940 26420
rect 44964 26364 45020 26420
rect 45044 26364 45100 26420
rect 45124 26364 45180 26420
rect 45204 26364 45260 26420
rect 46132 24484 46188 24540
rect 46212 24484 46268 24540
rect 46292 24484 46348 24540
rect 46372 24484 46428 24540
rect 46452 24484 46508 24540
rect 46532 24484 46588 24540
rect 46612 24484 46668 24540
rect 46692 24484 46748 24540
rect 46772 24484 46828 24540
rect 46852 24484 46908 24540
rect 46932 24484 46988 24540
rect 47012 24484 47068 24540
rect 47092 24484 47148 24540
rect 47172 24484 47228 24540
rect 47252 24484 47308 24540
rect 47332 24484 47388 24540
rect 47412 24484 47468 24540
rect 47492 24484 47548 24540
rect 47572 24484 47628 24540
rect 47652 24484 47708 24540
rect 43684 22604 43740 22660
rect 43764 22604 43820 22660
rect 43844 22604 43900 22660
rect 43924 22604 43980 22660
rect 44004 22604 44060 22660
rect 44084 22604 44140 22660
rect 44164 22604 44220 22660
rect 44244 22604 44300 22660
rect 44324 22604 44380 22660
rect 44404 22604 44460 22660
rect 44484 22604 44540 22660
rect 44564 22604 44620 22660
rect 44644 22604 44700 22660
rect 44724 22604 44780 22660
rect 44804 22604 44860 22660
rect 44884 22604 44940 22660
rect 44964 22604 45020 22660
rect 45044 22604 45100 22660
rect 45124 22604 45180 22660
rect 45204 22604 45260 22660
rect 46132 20724 46188 20780
rect 46212 20724 46268 20780
rect 46292 20724 46348 20780
rect 46372 20724 46428 20780
rect 46452 20724 46508 20780
rect 46532 20724 46588 20780
rect 46612 20724 46668 20780
rect 46692 20724 46748 20780
rect 46772 20724 46828 20780
rect 46852 20724 46908 20780
rect 46932 20724 46988 20780
rect 47012 20724 47068 20780
rect 47092 20724 47148 20780
rect 47172 20724 47228 20780
rect 47252 20724 47308 20780
rect 47332 20724 47388 20780
rect 47412 20724 47468 20780
rect 47492 20724 47548 20780
rect 47572 20724 47628 20780
rect 47652 20724 47708 20780
rect 43684 18844 43740 18900
rect 43764 18844 43820 18900
rect 43844 18844 43900 18900
rect 43924 18844 43980 18900
rect 44004 18844 44060 18900
rect 44084 18844 44140 18900
rect 44164 18844 44220 18900
rect 44244 18844 44300 18900
rect 44324 18844 44380 18900
rect 44404 18844 44460 18900
rect 44484 18844 44540 18900
rect 44564 18844 44620 18900
rect 44644 18844 44700 18900
rect 44724 18844 44780 18900
rect 44804 18844 44860 18900
rect 44884 18844 44940 18900
rect 44964 18844 45020 18900
rect 45044 18844 45100 18900
rect 45124 18844 45180 18900
rect 45204 18844 45260 18900
rect 16140 14814 16196 14870
rect 16220 14814 16276 14870
rect 16182 13394 16238 13450
rect 17130 13404 17186 13460
rect 16140 11054 16196 11110
rect 16220 11054 16276 11110
rect 16182 9634 16238 9690
rect 17130 9622 17186 9678
rect 19522 6450 19578 6506
rect 46132 16964 46188 17020
rect 46212 16964 46268 17020
rect 46292 16964 46348 17020
rect 46372 16964 46428 17020
rect 46452 16964 46508 17020
rect 46532 16964 46588 17020
rect 46612 16964 46668 17020
rect 46692 16964 46748 17020
rect 46772 16964 46828 17020
rect 46852 16964 46908 17020
rect 46932 16964 46988 17020
rect 47012 16964 47068 17020
rect 47092 16964 47148 17020
rect 47172 16964 47228 17020
rect 47252 16964 47308 17020
rect 47332 16964 47388 17020
rect 47412 16964 47468 17020
rect 47492 16964 47548 17020
rect 47572 16964 47628 17020
rect 47652 16964 47708 17020
rect 43684 15084 43740 15140
rect 43764 15084 43820 15140
rect 43844 15084 43900 15140
rect 43924 15084 43980 15140
rect 44004 15084 44060 15140
rect 44084 15084 44140 15140
rect 44164 15084 44220 15140
rect 44244 15084 44300 15140
rect 44324 15084 44380 15140
rect 44404 15084 44460 15140
rect 44484 15084 44540 15140
rect 44564 15084 44620 15140
rect 44644 15084 44700 15140
rect 44724 15084 44780 15140
rect 44804 15084 44860 15140
rect 44884 15084 44940 15140
rect 44964 15084 45020 15140
rect 45044 15084 45100 15140
rect 45124 15084 45180 15140
rect 45204 15084 45260 15140
rect 23662 11086 23718 11142
rect 25686 6450 25742 6506
rect 46132 13204 46188 13260
rect 46212 13204 46268 13260
rect 46292 13204 46348 13260
rect 46372 13204 46428 13260
rect 46452 13204 46508 13260
rect 46532 13204 46588 13260
rect 46612 13204 46668 13260
rect 46692 13204 46748 13260
rect 46772 13204 46828 13260
rect 46852 13204 46908 13260
rect 46932 13204 46988 13260
rect 47012 13204 47068 13260
rect 47092 13204 47148 13260
rect 47172 13204 47228 13260
rect 47252 13204 47308 13260
rect 47332 13204 47388 13260
rect 47412 13204 47468 13260
rect 47492 13204 47548 13260
rect 47572 13204 47628 13260
rect 47652 13204 47708 13260
rect 43684 11324 43740 11380
rect 43764 11324 43820 11380
rect 43844 11324 43900 11380
rect 43924 11324 43980 11380
rect 44004 11324 44060 11380
rect 44084 11324 44140 11380
rect 44164 11324 44220 11380
rect 44244 11324 44300 11380
rect 44324 11324 44380 11380
rect 44404 11324 44460 11380
rect 44484 11324 44540 11380
rect 44564 11324 44620 11380
rect 44644 11324 44700 11380
rect 44724 11324 44780 11380
rect 44804 11324 44860 11380
rect 44884 11324 44940 11380
rect 44964 11324 45020 11380
rect 45044 11324 45100 11380
rect 45124 11324 45180 11380
rect 45204 11324 45260 11380
rect 46132 9444 46188 9500
rect 46212 9444 46268 9500
rect 46292 9444 46348 9500
rect 46372 9444 46428 9500
rect 46452 9444 46508 9500
rect 46532 9444 46588 9500
rect 46612 9444 46668 9500
rect 46692 9444 46748 9500
rect 46772 9444 46828 9500
rect 46852 9444 46908 9500
rect 46932 9444 46988 9500
rect 47012 9444 47068 9500
rect 47092 9444 47148 9500
rect 47172 9444 47228 9500
rect 47252 9444 47308 9500
rect 47332 9444 47388 9500
rect 47412 9444 47468 9500
rect 47492 9444 47548 9500
rect 47572 9444 47628 9500
rect 47652 9444 47708 9500
rect 43684 7564 43740 7620
rect 43764 7564 43820 7620
rect 43844 7564 43900 7620
rect 43924 7564 43980 7620
rect 44004 7564 44060 7620
rect 44084 7564 44140 7620
rect 44164 7564 44220 7620
rect 44244 7564 44300 7620
rect 44324 7564 44380 7620
rect 44404 7564 44460 7620
rect 44484 7564 44540 7620
rect 44564 7564 44620 7620
rect 44644 7564 44700 7620
rect 44724 7564 44780 7620
rect 44804 7564 44860 7620
rect 44884 7564 44940 7620
rect 44964 7564 45020 7620
rect 45044 7564 45100 7620
rect 45124 7564 45180 7620
rect 45204 7564 45260 7620
rect 17774 6084 17830 6140
rect 28354 6112 28410 6140
rect 28354 6084 28356 6112
rect 28356 6084 28408 6112
rect 28408 6084 28410 6112
rect 928 5684 984 5740
rect 1008 5684 1064 5740
rect 1088 5684 1144 5740
rect 1168 5684 1224 5740
rect 1248 5684 1304 5740
rect 1328 5684 1384 5740
rect 1408 5684 1464 5740
rect 1488 5684 1544 5740
rect 1568 5684 1624 5740
rect 1648 5684 1704 5740
rect 1728 5684 1784 5740
rect 1808 5684 1864 5740
rect 1888 5684 1944 5740
rect 1968 5684 2024 5740
rect 2048 5684 2104 5740
rect 2128 5684 2184 5740
rect 2208 5684 2264 5740
rect 2288 5684 2344 5740
rect 2368 5684 2424 5740
rect 2448 5684 2504 5740
rect 46132 5684 46188 5740
rect 46212 5684 46268 5740
rect 46292 5684 46348 5740
rect 46372 5684 46428 5740
rect 46452 5684 46508 5740
rect 46532 5684 46588 5740
rect 46612 5684 46668 5740
rect 46692 5684 46748 5740
rect 46772 5684 46828 5740
rect 46852 5684 46908 5740
rect 46932 5684 46988 5740
rect 47012 5684 47068 5740
rect 47092 5684 47148 5740
rect 47172 5684 47228 5740
rect 47252 5684 47308 5740
rect 47332 5684 47388 5740
rect 47412 5684 47468 5740
rect 47492 5684 47548 5740
rect 47572 5684 47628 5740
rect 47652 5684 47708 5740
<< metal3 >>
rect 3348 41464 4980 41492
rect 3348 41400 3372 41464
rect 3436 41400 3452 41464
rect 3516 41400 3532 41464
rect 3596 41400 3612 41464
rect 3676 41400 3692 41464
rect 3756 41400 3772 41464
rect 3836 41400 3852 41464
rect 3916 41400 3932 41464
rect 3996 41400 4012 41464
rect 4076 41400 4092 41464
rect 4156 41400 4172 41464
rect 4236 41400 4252 41464
rect 4316 41400 4332 41464
rect 4396 41400 4412 41464
rect 4476 41400 4492 41464
rect 4556 41400 4572 41464
rect 4636 41400 4652 41464
rect 4716 41400 4732 41464
rect 4796 41400 4812 41464
rect 4876 41400 4892 41464
rect 4956 41400 4980 41464
rect 43656 41464 45288 41492
rect 12433 41402 12499 41403
rect 12428 41400 12434 41402
rect 3348 41372 4980 41400
rect 12344 41340 12434 41400
rect 12428 41338 12434 41340
rect 12498 41338 12504 41402
rect 43656 41400 43680 41464
rect 43744 41400 43760 41464
rect 43824 41400 43840 41464
rect 43904 41400 43920 41464
rect 43984 41400 44000 41464
rect 44064 41400 44080 41464
rect 44144 41400 44160 41464
rect 44224 41400 44240 41464
rect 44304 41400 44320 41464
rect 44384 41400 44400 41464
rect 44464 41400 44480 41464
rect 44544 41400 44560 41464
rect 44624 41400 44640 41464
rect 44704 41400 44720 41464
rect 44784 41400 44800 41464
rect 44864 41400 44880 41464
rect 44944 41400 44960 41464
rect 45024 41400 45040 41464
rect 45104 41400 45120 41464
rect 45184 41400 45200 41464
rect 45264 41400 45288 41464
rect 43656 41372 45288 41400
rect 12433 41337 12499 41338
rect 6798 41190 13970 41202
rect 6798 41134 6830 41190
rect 6886 41134 6910 41190
rect 6966 41174 13970 41190
rect 6966 41134 7414 41174
rect 6798 41110 7414 41134
rect 7478 41110 8133 41174
rect 8197 41110 8852 41174
rect 8916 41110 9571 41174
rect 9635 41110 10290 41174
rect 10354 41110 11009 41174
rect 11073 41110 11728 41174
rect 11792 41110 12447 41174
rect 12511 41110 13166 41174
rect 13230 41110 13885 41174
rect 13949 41110 13970 41174
rect 6798 41094 13970 41110
rect 6798 41030 7414 41094
rect 7478 41030 8133 41094
rect 8197 41030 8852 41094
rect 8916 41030 9571 41094
rect 9635 41030 10290 41094
rect 10354 41030 11009 41094
rect 11073 41030 11728 41094
rect 11792 41030 12447 41094
rect 12511 41030 13166 41094
rect 13230 41030 13885 41094
rect 13949 41030 13970 41094
rect 6798 41014 13970 41030
rect 6798 40950 7414 41014
rect 7478 40950 8133 41014
rect 8197 40950 8852 41014
rect 8916 40950 9571 41014
rect 9635 40950 10290 41014
rect 10354 40950 11009 41014
rect 11073 40950 11728 41014
rect 11792 40950 12447 41014
rect 12511 40950 13166 41014
rect 13230 40950 13885 41014
rect 13949 40950 13970 41014
rect 6798 40934 13970 40950
rect 6798 40870 7414 40934
rect 7478 40870 8133 40934
rect 8197 40870 8852 40934
rect 8916 40870 9571 40934
rect 9635 40870 10290 40934
rect 10354 40870 11009 40934
rect 11073 40870 11728 40934
rect 11792 40870 12447 40934
rect 12511 40870 13166 40934
rect 13230 40870 13885 40934
rect 13949 40870 13970 40934
rect 6798 40854 13970 40870
rect 6798 40790 7414 40854
rect 7478 40790 8133 40854
rect 8197 40790 8852 40854
rect 8916 40790 9571 40854
rect 9635 40790 10290 40854
rect 10354 40790 11009 40854
rect 11073 40790 11728 40854
rect 11792 40790 12447 40854
rect 12511 40790 13166 40854
rect 13230 40790 13885 40854
rect 13949 40790 13970 40854
rect 6798 40774 13970 40790
rect 6798 40710 7414 40774
rect 7478 40710 8133 40774
rect 8197 40710 8852 40774
rect 8916 40710 9571 40774
rect 9635 40710 10290 40774
rect 10354 40710 11009 40774
rect 11073 40710 11728 40774
rect 11792 40710 12447 40774
rect 12511 40710 13166 40774
rect 13230 40710 13885 40774
rect 13949 40710 13970 40774
rect 6798 40694 13970 40710
rect 6798 40630 7414 40694
rect 7478 40630 8133 40694
rect 8197 40630 8852 40694
rect 8916 40630 9571 40694
rect 9635 40630 10290 40694
rect 10354 40630 11009 40694
rect 11073 40630 11728 40694
rect 11792 40630 12447 40694
rect 12511 40630 13166 40694
rect 13230 40630 13885 40694
rect 13949 40630 13970 40694
rect 6798 40474 13970 40630
rect 6798 40410 7414 40474
rect 7478 40410 8133 40474
rect 8197 40410 8852 40474
rect 8916 40410 9571 40474
rect 9635 40410 10290 40474
rect 10354 40410 11009 40474
rect 11073 40410 11728 40474
rect 11792 40410 12447 40474
rect 12511 40410 13166 40474
rect 13230 40410 13885 40474
rect 13949 40410 13970 40474
rect 6798 40394 13970 40410
rect 6798 40330 7414 40394
rect 7478 40330 8133 40394
rect 8197 40330 8852 40394
rect 8916 40330 9571 40394
rect 9635 40330 10290 40394
rect 10354 40330 11009 40394
rect 11073 40330 11728 40394
rect 11792 40330 12447 40394
rect 12511 40330 13166 40394
rect 13230 40330 13885 40394
rect 13949 40330 13970 40394
rect 6798 40314 13970 40330
rect 6798 40250 7414 40314
rect 7478 40250 8133 40314
rect 8197 40250 8852 40314
rect 8916 40250 9571 40314
rect 9635 40250 10290 40314
rect 10354 40250 11009 40314
rect 11073 40250 11728 40314
rect 11792 40250 12447 40314
rect 12511 40250 13166 40314
rect 13230 40250 13885 40314
rect 13949 40250 13970 40314
rect 6798 40234 13970 40250
rect 6798 40170 7414 40234
rect 7478 40170 8133 40234
rect 8197 40170 8852 40234
rect 8916 40170 9571 40234
rect 9635 40170 10290 40234
rect 10354 40170 11009 40234
rect 11073 40170 11728 40234
rect 11792 40170 12447 40234
rect 12511 40170 13166 40234
rect 13230 40170 13885 40234
rect 13949 40170 13970 40234
rect 6798 40154 13970 40170
rect 6798 40090 7414 40154
rect 7478 40090 8133 40154
rect 8197 40090 8852 40154
rect 8916 40090 9571 40154
rect 9635 40090 10290 40154
rect 10354 40090 11009 40154
rect 11073 40090 11728 40154
rect 11792 40090 12447 40154
rect 12511 40090 13166 40154
rect 13230 40090 13885 40154
rect 13949 40090 13970 40154
rect 6798 40074 13970 40090
rect 6798 40010 7414 40074
rect 7478 40010 8133 40074
rect 8197 40010 8852 40074
rect 8916 40010 9571 40074
rect 9635 40010 10290 40074
rect 10354 40010 11009 40074
rect 11073 40010 11728 40074
rect 11792 40010 12447 40074
rect 12511 40010 13166 40074
rect 13230 40010 13885 40074
rect 13949 40010 13970 40074
rect 6798 39994 13970 40010
rect 6798 39930 7414 39994
rect 7478 39930 8133 39994
rect 8197 39930 8852 39994
rect 8916 39930 9571 39994
rect 9635 39930 10290 39994
rect 10354 39930 11009 39994
rect 11073 39930 11728 39994
rect 11792 39930 12447 39994
rect 12511 39930 13166 39994
rect 13230 39930 13885 39994
rect 13949 39930 13970 39994
rect 6798 39902 13970 39930
rect 6800 39774 7000 39802
rect 6800 39710 6828 39774
rect 6892 39770 6908 39774
rect 6892 39710 6908 39714
rect 6972 39710 7000 39774
rect 6800 39682 7000 39710
rect 13670 39630 13676 39694
rect 13740 39692 13746 39694
rect 15009 39692 15075 39695
rect 27613 39694 27679 39695
rect 27608 39692 27614 39694
rect 13740 39690 15075 39692
rect 13740 39634 15014 39690
rect 15070 39634 15075 39690
rect 13740 39632 15075 39634
rect 27524 39632 27614 39692
rect 13740 39630 13746 39632
rect 15009 39629 15075 39632
rect 27608 39630 27614 39632
rect 27678 39630 27684 39694
rect 27613 39629 27679 39630
rect 900 39584 2532 39612
rect 900 39520 924 39584
rect 988 39520 1004 39584
rect 1068 39520 1084 39584
rect 1148 39520 1164 39584
rect 1228 39520 1244 39584
rect 1308 39520 1324 39584
rect 1388 39520 1404 39584
rect 1468 39520 1484 39584
rect 1548 39520 1564 39584
rect 1628 39520 1644 39584
rect 1708 39520 1724 39584
rect 1788 39520 1804 39584
rect 1868 39520 1884 39584
rect 1948 39520 1964 39584
rect 2028 39520 2044 39584
rect 2108 39520 2124 39584
rect 2188 39520 2204 39584
rect 2268 39520 2284 39584
rect 2348 39520 2364 39584
rect 2428 39520 2444 39584
rect 2508 39520 2532 39584
rect 900 39492 2532 39520
rect 46104 39584 47736 39612
rect 46104 39520 46128 39584
rect 46192 39520 46208 39584
rect 46272 39520 46288 39584
rect 46352 39520 46368 39584
rect 46432 39520 46448 39584
rect 46512 39520 46528 39584
rect 46592 39520 46608 39584
rect 46672 39520 46688 39584
rect 46752 39520 46768 39584
rect 46832 39520 46848 39584
rect 46912 39520 46928 39584
rect 46992 39520 47008 39584
rect 47072 39520 47088 39584
rect 47152 39520 47168 39584
rect 47232 39520 47248 39584
rect 47312 39520 47328 39584
rect 47392 39520 47408 39584
rect 47472 39520 47488 39584
rect 47552 39520 47568 39584
rect 47632 39520 47648 39584
rect 47712 39520 47736 39584
rect 46104 39492 47736 39520
rect 3348 37704 4980 37732
rect 3348 37640 3372 37704
rect 3436 37640 3452 37704
rect 3516 37640 3532 37704
rect 3596 37640 3612 37704
rect 3676 37640 3692 37704
rect 3756 37640 3772 37704
rect 3836 37640 3852 37704
rect 3916 37640 3932 37704
rect 3996 37640 4012 37704
rect 4076 37640 4092 37704
rect 4156 37640 4172 37704
rect 4236 37640 4252 37704
rect 4316 37640 4332 37704
rect 4396 37640 4412 37704
rect 4476 37640 4492 37704
rect 4556 37640 4572 37704
rect 4636 37640 4652 37704
rect 4716 37640 4732 37704
rect 4796 37640 4812 37704
rect 4876 37640 4892 37704
rect 4956 37640 4980 37704
rect 3348 37612 4980 37640
rect 43656 37704 45288 37732
rect 43656 37640 43680 37704
rect 43744 37640 43760 37704
rect 43824 37640 43840 37704
rect 43904 37640 43920 37704
rect 43984 37640 44000 37704
rect 44064 37640 44080 37704
rect 44144 37640 44160 37704
rect 44224 37640 44240 37704
rect 44304 37640 44320 37704
rect 44384 37640 44400 37704
rect 44464 37640 44480 37704
rect 44544 37640 44560 37704
rect 44624 37640 44640 37704
rect 44704 37640 44720 37704
rect 44784 37640 44800 37704
rect 44864 37640 44880 37704
rect 44944 37640 44960 37704
rect 45024 37640 45040 37704
rect 45104 37640 45120 37704
rect 45184 37640 45200 37704
rect 45264 37640 45288 37704
rect 12985 37620 13051 37621
rect 16849 37620 16915 37621
rect 27889 37620 27955 37621
rect 12980 37618 12986 37620
rect 12896 37558 12986 37618
rect 12980 37556 12986 37558
rect 13050 37556 13056 37620
rect 16844 37618 16850 37620
rect 16760 37558 16850 37618
rect 16844 37556 16850 37558
rect 16914 37556 16920 37620
rect 27884 37618 27890 37620
rect 27800 37558 27890 37618
rect 27884 37556 27890 37558
rect 27954 37556 27960 37620
rect 43656 37612 45288 37640
rect 12985 37555 13051 37556
rect 16849 37555 16915 37556
rect 27889 37555 27955 37556
rect 5916 37430 13088 37442
rect 5916 37374 5948 37430
rect 6004 37374 6028 37430
rect 6084 37414 13088 37430
rect 6084 37374 6532 37414
rect 5916 37350 6532 37374
rect 6596 37350 7251 37414
rect 7315 37350 7970 37414
rect 8034 37350 8689 37414
rect 8753 37350 9408 37414
rect 9472 37350 10127 37414
rect 10191 37350 10846 37414
rect 10910 37350 11565 37414
rect 11629 37350 12284 37414
rect 12348 37350 13003 37414
rect 13067 37350 13088 37414
rect 5916 37334 13088 37350
rect 5916 37270 6532 37334
rect 6596 37270 7251 37334
rect 7315 37270 7970 37334
rect 8034 37270 8689 37334
rect 8753 37270 9408 37334
rect 9472 37270 10127 37334
rect 10191 37270 10846 37334
rect 10910 37270 11565 37334
rect 11629 37270 12284 37334
rect 12348 37270 13003 37334
rect 13067 37270 13088 37334
rect 5916 37254 13088 37270
rect 5916 37190 6532 37254
rect 6596 37190 7251 37254
rect 7315 37190 7970 37254
rect 8034 37190 8689 37254
rect 8753 37190 9408 37254
rect 9472 37190 10127 37254
rect 10191 37190 10846 37254
rect 10910 37190 11565 37254
rect 11629 37190 12284 37254
rect 12348 37190 13003 37254
rect 13067 37190 13088 37254
rect 5916 37174 13088 37190
rect 5916 37110 6532 37174
rect 6596 37110 7251 37174
rect 7315 37110 7970 37174
rect 8034 37110 8689 37174
rect 8753 37110 9408 37174
rect 9472 37110 10127 37174
rect 10191 37110 10846 37174
rect 10910 37110 11565 37174
rect 11629 37110 12284 37174
rect 12348 37110 13003 37174
rect 13067 37110 13088 37174
rect 5916 37094 13088 37110
rect 5916 37030 6532 37094
rect 6596 37030 7251 37094
rect 7315 37030 7970 37094
rect 8034 37030 8689 37094
rect 8753 37030 9408 37094
rect 9472 37030 10127 37094
rect 10191 37030 10846 37094
rect 10910 37030 11565 37094
rect 11629 37030 12284 37094
rect 12348 37030 13003 37094
rect 13067 37030 13088 37094
rect 5916 37014 13088 37030
rect 5916 36950 6532 37014
rect 6596 36950 7251 37014
rect 7315 36950 7970 37014
rect 8034 36950 8689 37014
rect 8753 36950 9408 37014
rect 9472 36950 10127 37014
rect 10191 36950 10846 37014
rect 10910 36950 11565 37014
rect 11629 36950 12284 37014
rect 12348 36950 13003 37014
rect 13067 36950 13088 37014
rect 5916 36934 13088 36950
rect 5916 36870 6532 36934
rect 6596 36870 7251 36934
rect 7315 36870 7970 36934
rect 8034 36870 8689 36934
rect 8753 36870 9408 36934
rect 9472 36870 10127 36934
rect 10191 36870 10846 36934
rect 10910 36870 11565 36934
rect 11629 36870 12284 36934
rect 12348 36870 13003 36934
rect 13067 36870 13088 36934
rect 5916 36714 13088 36870
rect 5916 36650 6532 36714
rect 6596 36650 7251 36714
rect 7315 36650 7970 36714
rect 8034 36650 8689 36714
rect 8753 36650 9408 36714
rect 9472 36650 10127 36714
rect 10191 36650 10846 36714
rect 10910 36650 11565 36714
rect 11629 36650 12284 36714
rect 12348 36650 13003 36714
rect 13067 36650 13088 36714
rect 5916 36634 13088 36650
rect 5916 36570 6532 36634
rect 6596 36570 7251 36634
rect 7315 36570 7970 36634
rect 8034 36570 8689 36634
rect 8753 36570 9408 36634
rect 9472 36570 10127 36634
rect 10191 36570 10846 36634
rect 10910 36570 11565 36634
rect 11629 36570 12284 36634
rect 12348 36570 13003 36634
rect 13067 36570 13088 36634
rect 5916 36554 13088 36570
rect 5916 36490 6532 36554
rect 6596 36490 7251 36554
rect 7315 36490 7970 36554
rect 8034 36490 8689 36554
rect 8753 36490 9408 36554
rect 9472 36490 10127 36554
rect 10191 36490 10846 36554
rect 10910 36490 11565 36554
rect 11629 36490 12284 36554
rect 12348 36490 13003 36554
rect 13067 36490 13088 36554
rect 5916 36474 13088 36490
rect 5916 36410 6532 36474
rect 6596 36410 7251 36474
rect 7315 36410 7970 36474
rect 8034 36410 8689 36474
rect 8753 36410 9408 36474
rect 9472 36410 10127 36474
rect 10191 36410 10846 36474
rect 10910 36410 11565 36474
rect 11629 36410 12284 36474
rect 12348 36410 13003 36474
rect 13067 36410 13088 36474
rect 5916 36394 13088 36410
rect 5916 36330 6532 36394
rect 6596 36330 7251 36394
rect 7315 36330 7970 36394
rect 8034 36330 8689 36394
rect 8753 36330 9408 36394
rect 9472 36330 10127 36394
rect 10191 36330 10846 36394
rect 10910 36330 11565 36394
rect 11629 36330 12284 36394
rect 12348 36330 13003 36394
rect 13067 36330 13088 36394
rect 5916 36314 13088 36330
rect 5916 36250 6532 36314
rect 6596 36250 7251 36314
rect 7315 36250 7970 36314
rect 8034 36250 8689 36314
rect 8753 36250 9408 36314
rect 9472 36250 10127 36314
rect 10191 36250 10846 36314
rect 10910 36250 11565 36314
rect 11629 36250 12284 36314
rect 12348 36250 13003 36314
rect 13067 36250 13088 36314
rect 5916 36234 13088 36250
rect 5916 36170 6532 36234
rect 6596 36170 7251 36234
rect 7315 36170 7970 36234
rect 8034 36170 8689 36234
rect 8753 36170 9408 36234
rect 9472 36170 10127 36234
rect 10191 36170 10846 36234
rect 10910 36170 11565 36234
rect 11629 36170 12284 36234
rect 12348 36170 13003 36234
rect 13067 36170 13088 36234
rect 5916 36142 13088 36170
rect 13364 37430 20536 37442
rect 13364 37374 13396 37430
rect 13452 37374 13476 37430
rect 13532 37414 20536 37430
rect 13532 37374 13980 37414
rect 13364 37350 13980 37374
rect 14044 37350 14699 37414
rect 14763 37350 15418 37414
rect 15482 37350 16137 37414
rect 16201 37350 16856 37414
rect 16920 37350 17575 37414
rect 17639 37350 18294 37414
rect 18358 37350 19013 37414
rect 19077 37350 19732 37414
rect 19796 37350 20451 37414
rect 20515 37350 20536 37414
rect 13364 37334 20536 37350
rect 13364 37270 13980 37334
rect 14044 37270 14699 37334
rect 14763 37270 15418 37334
rect 15482 37270 16137 37334
rect 16201 37270 16856 37334
rect 16920 37270 17575 37334
rect 17639 37270 18294 37334
rect 18358 37270 19013 37334
rect 19077 37270 19732 37334
rect 19796 37270 20451 37334
rect 20515 37270 20536 37334
rect 13364 37254 20536 37270
rect 13364 37190 13980 37254
rect 14044 37190 14699 37254
rect 14763 37190 15418 37254
rect 15482 37190 16137 37254
rect 16201 37190 16856 37254
rect 16920 37190 17575 37254
rect 17639 37190 18294 37254
rect 18358 37190 19013 37254
rect 19077 37190 19732 37254
rect 19796 37190 20451 37254
rect 20515 37190 20536 37254
rect 13364 37174 20536 37190
rect 13364 37110 13980 37174
rect 14044 37110 14699 37174
rect 14763 37110 15418 37174
rect 15482 37110 16137 37174
rect 16201 37110 16856 37174
rect 16920 37110 17575 37174
rect 17639 37110 18294 37174
rect 18358 37110 19013 37174
rect 19077 37110 19732 37174
rect 19796 37110 20451 37174
rect 20515 37110 20536 37174
rect 13364 37094 20536 37110
rect 13364 37030 13980 37094
rect 14044 37030 14699 37094
rect 14763 37030 15418 37094
rect 15482 37030 16137 37094
rect 16201 37030 16856 37094
rect 16920 37030 17575 37094
rect 17639 37030 18294 37094
rect 18358 37030 19013 37094
rect 19077 37030 19732 37094
rect 19796 37030 20451 37094
rect 20515 37030 20536 37094
rect 13364 37014 20536 37030
rect 13364 36950 13980 37014
rect 14044 36950 14699 37014
rect 14763 36950 15418 37014
rect 15482 36950 16137 37014
rect 16201 36950 16856 37014
rect 16920 36950 17575 37014
rect 17639 36950 18294 37014
rect 18358 36950 19013 37014
rect 19077 36950 19732 37014
rect 19796 36950 20451 37014
rect 20515 36950 20536 37014
rect 13364 36934 20536 36950
rect 13364 36870 13980 36934
rect 14044 36870 14699 36934
rect 14763 36870 15418 36934
rect 15482 36870 16137 36934
rect 16201 36870 16856 36934
rect 16920 36870 17575 36934
rect 17639 36870 18294 36934
rect 18358 36870 19013 36934
rect 19077 36870 19732 36934
rect 19796 36870 20451 36934
rect 20515 36870 20536 36934
rect 13364 36714 20536 36870
rect 13364 36650 13980 36714
rect 14044 36650 14699 36714
rect 14763 36650 15418 36714
rect 15482 36650 16137 36714
rect 16201 36650 16856 36714
rect 16920 36650 17575 36714
rect 17639 36650 18294 36714
rect 18358 36650 19013 36714
rect 19077 36650 19732 36714
rect 19796 36650 20451 36714
rect 20515 36650 20536 36714
rect 13364 36634 20536 36650
rect 13364 36570 13980 36634
rect 14044 36570 14699 36634
rect 14763 36570 15418 36634
rect 15482 36570 16137 36634
rect 16201 36570 16856 36634
rect 16920 36570 17575 36634
rect 17639 36570 18294 36634
rect 18358 36570 19013 36634
rect 19077 36570 19732 36634
rect 19796 36570 20451 36634
rect 20515 36570 20536 36634
rect 13364 36554 20536 36570
rect 13364 36490 13980 36554
rect 14044 36490 14699 36554
rect 14763 36490 15418 36554
rect 15482 36490 16137 36554
rect 16201 36490 16856 36554
rect 16920 36490 17575 36554
rect 17639 36490 18294 36554
rect 18358 36490 19013 36554
rect 19077 36490 19732 36554
rect 19796 36490 20451 36554
rect 20515 36490 20536 36554
rect 13364 36474 20536 36490
rect 13364 36410 13980 36474
rect 14044 36410 14699 36474
rect 14763 36410 15418 36474
rect 15482 36410 16137 36474
rect 16201 36410 16856 36474
rect 16920 36410 17575 36474
rect 17639 36410 18294 36474
rect 18358 36410 19013 36474
rect 19077 36410 19732 36474
rect 19796 36410 20451 36474
rect 20515 36410 20536 36474
rect 13364 36394 20536 36410
rect 13364 36330 13980 36394
rect 14044 36330 14699 36394
rect 14763 36330 15418 36394
rect 15482 36330 16137 36394
rect 16201 36330 16856 36394
rect 16920 36330 17575 36394
rect 17639 36330 18294 36394
rect 18358 36330 19013 36394
rect 19077 36330 19732 36394
rect 19796 36330 20451 36394
rect 20515 36330 20536 36394
rect 13364 36314 20536 36330
rect 13364 36250 13980 36314
rect 14044 36250 14699 36314
rect 14763 36250 15418 36314
rect 15482 36250 16137 36314
rect 16201 36250 16856 36314
rect 16920 36250 17575 36314
rect 17639 36250 18294 36314
rect 18358 36250 19013 36314
rect 19077 36250 19732 36314
rect 19796 36250 20451 36314
rect 20515 36250 20536 36314
rect 13364 36234 20536 36250
rect 13364 36170 13980 36234
rect 14044 36170 14699 36234
rect 14763 36170 15418 36234
rect 15482 36170 16137 36234
rect 16201 36170 16856 36234
rect 16920 36170 17575 36234
rect 17639 36170 18294 36234
rect 18358 36170 19013 36234
rect 19077 36170 19732 36234
rect 19796 36170 20451 36234
rect 20515 36170 20536 36234
rect 13364 36142 20536 36170
rect 20812 37430 27984 37442
rect 20812 37374 20844 37430
rect 20900 37374 20924 37430
rect 20980 37414 27984 37430
rect 20980 37374 21428 37414
rect 20812 37350 21428 37374
rect 21492 37350 22147 37414
rect 22211 37350 22866 37414
rect 22930 37350 23585 37414
rect 23649 37350 24304 37414
rect 24368 37350 25023 37414
rect 25087 37350 25742 37414
rect 25806 37350 26461 37414
rect 26525 37350 27180 37414
rect 27244 37350 27899 37414
rect 27963 37350 27984 37414
rect 20812 37334 27984 37350
rect 20812 37270 21428 37334
rect 21492 37270 22147 37334
rect 22211 37270 22866 37334
rect 22930 37270 23585 37334
rect 23649 37270 24304 37334
rect 24368 37270 25023 37334
rect 25087 37270 25742 37334
rect 25806 37270 26461 37334
rect 26525 37270 27180 37334
rect 27244 37270 27899 37334
rect 27963 37270 27984 37334
rect 20812 37254 27984 37270
rect 20812 37190 21428 37254
rect 21492 37190 22147 37254
rect 22211 37190 22866 37254
rect 22930 37190 23585 37254
rect 23649 37190 24304 37254
rect 24368 37190 25023 37254
rect 25087 37190 25742 37254
rect 25806 37190 26461 37254
rect 26525 37190 27180 37254
rect 27244 37190 27899 37254
rect 27963 37190 27984 37254
rect 20812 37174 27984 37190
rect 20812 37110 21428 37174
rect 21492 37110 22147 37174
rect 22211 37110 22866 37174
rect 22930 37110 23585 37174
rect 23649 37110 24304 37174
rect 24368 37110 25023 37174
rect 25087 37110 25742 37174
rect 25806 37110 26461 37174
rect 26525 37110 27180 37174
rect 27244 37110 27899 37174
rect 27963 37110 27984 37174
rect 20812 37094 27984 37110
rect 20812 37030 21428 37094
rect 21492 37030 22147 37094
rect 22211 37030 22866 37094
rect 22930 37030 23585 37094
rect 23649 37030 24304 37094
rect 24368 37030 25023 37094
rect 25087 37030 25742 37094
rect 25806 37030 26461 37094
rect 26525 37030 27180 37094
rect 27244 37030 27899 37094
rect 27963 37030 27984 37094
rect 20812 37014 27984 37030
rect 20812 36950 21428 37014
rect 21492 36950 22147 37014
rect 22211 36950 22866 37014
rect 22930 36950 23585 37014
rect 23649 36950 24304 37014
rect 24368 36950 25023 37014
rect 25087 36950 25742 37014
rect 25806 36950 26461 37014
rect 26525 36950 27180 37014
rect 27244 36950 27899 37014
rect 27963 36950 27984 37014
rect 20812 36934 27984 36950
rect 20812 36870 21428 36934
rect 21492 36870 22147 36934
rect 22211 36870 22866 36934
rect 22930 36870 23585 36934
rect 23649 36870 24304 36934
rect 24368 36870 25023 36934
rect 25087 36870 25742 36934
rect 25806 36870 26461 36934
rect 26525 36870 27180 36934
rect 27244 36870 27899 36934
rect 27963 36870 27984 36934
rect 20812 36714 27984 36870
rect 20812 36650 21428 36714
rect 21492 36650 22147 36714
rect 22211 36650 22866 36714
rect 22930 36650 23585 36714
rect 23649 36650 24304 36714
rect 24368 36650 25023 36714
rect 25087 36650 25742 36714
rect 25806 36650 26461 36714
rect 26525 36650 27180 36714
rect 27244 36650 27899 36714
rect 27963 36650 27984 36714
rect 20812 36634 27984 36650
rect 20812 36570 21428 36634
rect 21492 36570 22147 36634
rect 22211 36570 22866 36634
rect 22930 36570 23585 36634
rect 23649 36570 24304 36634
rect 24368 36570 25023 36634
rect 25087 36570 25742 36634
rect 25806 36570 26461 36634
rect 26525 36570 27180 36634
rect 27244 36570 27899 36634
rect 27963 36570 27984 36634
rect 20812 36554 27984 36570
rect 20812 36490 21428 36554
rect 21492 36490 22147 36554
rect 22211 36490 22866 36554
rect 22930 36490 23585 36554
rect 23649 36490 24304 36554
rect 24368 36490 25023 36554
rect 25087 36490 25742 36554
rect 25806 36490 26461 36554
rect 26525 36490 27180 36554
rect 27244 36490 27899 36554
rect 27963 36490 27984 36554
rect 20812 36474 27984 36490
rect 20812 36410 21428 36474
rect 21492 36410 22147 36474
rect 22211 36410 22866 36474
rect 22930 36410 23585 36474
rect 23649 36410 24304 36474
rect 24368 36410 25023 36474
rect 25087 36410 25742 36474
rect 25806 36410 26461 36474
rect 26525 36410 27180 36474
rect 27244 36410 27899 36474
rect 27963 36410 27984 36474
rect 20812 36394 27984 36410
rect 20812 36330 21428 36394
rect 21492 36330 22147 36394
rect 22211 36330 22866 36394
rect 22930 36330 23585 36394
rect 23649 36330 24304 36394
rect 24368 36330 25023 36394
rect 25087 36330 25742 36394
rect 25806 36330 26461 36394
rect 26525 36330 27180 36394
rect 27244 36330 27899 36394
rect 27963 36330 27984 36394
rect 20812 36314 27984 36330
rect 20812 36250 21428 36314
rect 21492 36250 22147 36314
rect 22211 36250 22866 36314
rect 22930 36250 23585 36314
rect 23649 36250 24304 36314
rect 24368 36250 25023 36314
rect 25087 36250 25742 36314
rect 25806 36250 26461 36314
rect 26525 36250 27180 36314
rect 27244 36250 27899 36314
rect 27963 36250 27984 36314
rect 20812 36234 27984 36250
rect 20812 36170 21428 36234
rect 21492 36170 22147 36234
rect 22211 36170 22866 36234
rect 22930 36170 23585 36234
rect 23649 36170 24304 36234
rect 24368 36170 25023 36234
rect 25087 36170 25742 36234
rect 25806 36170 26461 36234
rect 26525 36170 27180 36234
rect 27244 36170 27899 36234
rect 27963 36170 27984 36234
rect 20812 36142 27984 36170
rect 5918 36014 6118 36042
rect 5918 35950 5946 36014
rect 6010 36010 6026 36014
rect 6010 35950 6026 35954
rect 6090 35950 6118 36014
rect 5918 35922 6118 35950
rect 13366 36014 13566 36042
rect 13366 35950 13394 36014
rect 13458 36010 13474 36014
rect 13458 35950 13474 35954
rect 13538 35950 13566 36014
rect 13366 35922 13566 35950
rect 20814 36014 21014 36042
rect 20814 35950 20842 36014
rect 20906 36010 20922 36014
rect 20906 35950 20922 35954
rect 20986 35950 21014 36014
rect 20814 35922 21014 35950
rect 900 35824 2532 35852
rect 900 35760 924 35824
rect 988 35760 1004 35824
rect 1068 35760 1084 35824
rect 1148 35760 1164 35824
rect 1228 35760 1244 35824
rect 1308 35760 1324 35824
rect 1388 35760 1404 35824
rect 1468 35760 1484 35824
rect 1548 35760 1564 35824
rect 1628 35760 1644 35824
rect 1708 35760 1724 35824
rect 1788 35760 1804 35824
rect 1868 35760 1884 35824
rect 1948 35760 1964 35824
rect 2028 35760 2044 35824
rect 2108 35760 2124 35824
rect 2188 35760 2204 35824
rect 2268 35760 2284 35824
rect 2348 35760 2364 35824
rect 2428 35760 2444 35824
rect 2508 35760 2532 35824
rect 900 35732 2532 35760
rect 46104 35824 47736 35852
rect 46104 35760 46128 35824
rect 46192 35760 46208 35824
rect 46272 35760 46288 35824
rect 46352 35760 46368 35824
rect 46432 35760 46448 35824
rect 46512 35760 46528 35824
rect 46592 35760 46608 35824
rect 46672 35760 46688 35824
rect 46752 35760 46768 35824
rect 46832 35760 46848 35824
rect 46912 35760 46928 35824
rect 46992 35760 47008 35824
rect 47072 35760 47088 35824
rect 47152 35760 47168 35824
rect 47232 35760 47248 35824
rect 47312 35760 47328 35824
rect 47392 35760 47408 35824
rect 47472 35760 47488 35824
rect 47552 35760 47568 35824
rect 47632 35760 47648 35824
rect 47712 35760 47736 35824
rect 46104 35732 47736 35760
rect 3348 33944 4980 33972
rect 3348 33880 3372 33944
rect 3436 33880 3452 33944
rect 3516 33880 3532 33944
rect 3596 33880 3612 33944
rect 3676 33880 3692 33944
rect 3756 33880 3772 33944
rect 3836 33880 3852 33944
rect 3916 33880 3932 33944
rect 3996 33880 4012 33944
rect 4076 33880 4092 33944
rect 4156 33880 4172 33944
rect 4236 33880 4252 33944
rect 4316 33880 4332 33944
rect 4396 33880 4412 33944
rect 4476 33880 4492 33944
rect 4556 33880 4572 33944
rect 4636 33880 4652 33944
rect 4716 33880 4732 33944
rect 4796 33880 4812 33944
rect 4876 33880 4892 33944
rect 4956 33880 4980 33944
rect 3348 33852 4980 33880
rect 43656 33944 45288 33972
rect 43656 33880 43680 33944
rect 43744 33880 43760 33944
rect 43824 33880 43840 33944
rect 43904 33880 43920 33944
rect 43984 33880 44000 33944
rect 44064 33880 44080 33944
rect 44144 33880 44160 33944
rect 44224 33880 44240 33944
rect 44304 33880 44320 33944
rect 44384 33880 44400 33944
rect 44464 33880 44480 33944
rect 44544 33880 44560 33944
rect 44624 33880 44640 33944
rect 44704 33880 44720 33944
rect 44784 33880 44800 33944
rect 44864 33880 44880 33944
rect 44944 33880 44960 33944
rect 45024 33880 45040 33944
rect 45104 33880 45120 33944
rect 45184 33880 45200 33944
rect 45264 33880 45288 33944
rect 43656 33852 45288 33880
rect 9949 33836 10015 33839
rect 10082 33836 10088 33838
rect 9949 33834 10088 33836
rect 9949 33778 9954 33834
rect 10010 33778 10088 33834
rect 9949 33776 10088 33778
rect 9949 33773 10015 33776
rect 10082 33774 10088 33776
rect 10152 33774 10158 33838
rect 6602 33670 13774 33682
rect 6602 33614 6634 33670
rect 6690 33614 6714 33670
rect 6770 33654 13774 33670
rect 6770 33614 7218 33654
rect 6602 33590 7218 33614
rect 7282 33590 7937 33654
rect 8001 33590 8656 33654
rect 8720 33590 9375 33654
rect 9439 33590 10094 33654
rect 10158 33590 10813 33654
rect 10877 33590 11532 33654
rect 11596 33590 12251 33654
rect 12315 33590 12970 33654
rect 13034 33590 13689 33654
rect 13753 33590 13774 33654
rect 6602 33574 13774 33590
rect 6602 33510 7218 33574
rect 7282 33510 7937 33574
rect 8001 33510 8656 33574
rect 8720 33510 9375 33574
rect 9439 33510 10094 33574
rect 10158 33510 10813 33574
rect 10877 33510 11532 33574
rect 11596 33510 12251 33574
rect 12315 33510 12970 33574
rect 13034 33510 13689 33574
rect 13753 33510 13774 33574
rect 6602 33494 13774 33510
rect 6602 33430 7218 33494
rect 7282 33430 7937 33494
rect 8001 33430 8656 33494
rect 8720 33430 9375 33494
rect 9439 33430 10094 33494
rect 10158 33430 10813 33494
rect 10877 33430 11532 33494
rect 11596 33430 12251 33494
rect 12315 33430 12970 33494
rect 13034 33430 13689 33494
rect 13753 33430 13774 33494
rect 6602 33414 13774 33430
rect 6602 33350 7218 33414
rect 7282 33350 7937 33414
rect 8001 33350 8656 33414
rect 8720 33350 9375 33414
rect 9439 33350 10094 33414
rect 10158 33350 10813 33414
rect 10877 33350 11532 33414
rect 11596 33350 12251 33414
rect 12315 33350 12970 33414
rect 13034 33350 13689 33414
rect 13753 33350 13774 33414
rect 6602 33334 13774 33350
rect 6602 33270 7218 33334
rect 7282 33270 7937 33334
rect 8001 33270 8656 33334
rect 8720 33270 9375 33334
rect 9439 33270 10094 33334
rect 10158 33270 10813 33334
rect 10877 33270 11532 33334
rect 11596 33270 12251 33334
rect 12315 33270 12970 33334
rect 13034 33270 13689 33334
rect 13753 33270 13774 33334
rect 6602 33254 13774 33270
rect 6602 33190 7218 33254
rect 7282 33190 7937 33254
rect 8001 33190 8656 33254
rect 8720 33190 9375 33254
rect 9439 33190 10094 33254
rect 10158 33190 10813 33254
rect 10877 33190 11532 33254
rect 11596 33190 12251 33254
rect 12315 33190 12970 33254
rect 13034 33190 13689 33254
rect 13753 33190 13774 33254
rect 6602 33174 13774 33190
rect 6602 33110 7218 33174
rect 7282 33110 7937 33174
rect 8001 33110 8656 33174
rect 8720 33110 9375 33174
rect 9439 33110 10094 33174
rect 10158 33110 10813 33174
rect 10877 33110 11532 33174
rect 11596 33110 12251 33174
rect 12315 33110 12970 33174
rect 13034 33110 13689 33174
rect 13753 33110 13774 33174
rect 6602 32954 13774 33110
rect 6602 32890 7218 32954
rect 7282 32890 7937 32954
rect 8001 32890 8656 32954
rect 8720 32890 9375 32954
rect 9439 32890 10094 32954
rect 10158 32890 10813 32954
rect 10877 32890 11532 32954
rect 11596 32890 12251 32954
rect 12315 32890 12970 32954
rect 13034 32890 13689 32954
rect 13753 32890 13774 32954
rect 6602 32874 13774 32890
rect 6602 32810 7218 32874
rect 7282 32810 7937 32874
rect 8001 32810 8656 32874
rect 8720 32810 9375 32874
rect 9439 32810 10094 32874
rect 10158 32810 10813 32874
rect 10877 32810 11532 32874
rect 11596 32810 12251 32874
rect 12315 32810 12970 32874
rect 13034 32810 13689 32874
rect 13753 32810 13774 32874
rect 6602 32794 13774 32810
rect 6602 32730 7218 32794
rect 7282 32730 7937 32794
rect 8001 32730 8656 32794
rect 8720 32730 9375 32794
rect 9439 32730 10094 32794
rect 10158 32730 10813 32794
rect 10877 32730 11532 32794
rect 11596 32730 12251 32794
rect 12315 32730 12970 32794
rect 13034 32730 13689 32794
rect 13753 32730 13774 32794
rect 6602 32714 13774 32730
rect 6602 32650 7218 32714
rect 7282 32650 7937 32714
rect 8001 32650 8656 32714
rect 8720 32650 9375 32714
rect 9439 32650 10094 32714
rect 10158 32650 10813 32714
rect 10877 32650 11532 32714
rect 11596 32650 12251 32714
rect 12315 32650 12970 32714
rect 13034 32650 13689 32714
rect 13753 32650 13774 32714
rect 6602 32634 13774 32650
rect 6602 32570 7218 32634
rect 7282 32570 7937 32634
rect 8001 32570 8656 32634
rect 8720 32570 9375 32634
rect 9439 32570 10094 32634
rect 10158 32570 10813 32634
rect 10877 32570 11532 32634
rect 11596 32570 12251 32634
rect 12315 32570 12970 32634
rect 13034 32570 13689 32634
rect 13753 32570 13774 32634
rect 6602 32554 13774 32570
rect 6602 32490 7218 32554
rect 7282 32490 7937 32554
rect 8001 32490 8656 32554
rect 8720 32490 9375 32554
rect 9439 32490 10094 32554
rect 10158 32490 10813 32554
rect 10877 32490 11532 32554
rect 11596 32490 12251 32554
rect 12315 32490 12970 32554
rect 13034 32490 13689 32554
rect 13753 32490 13774 32554
rect 6602 32474 13774 32490
rect 6602 32410 7218 32474
rect 7282 32410 7937 32474
rect 8001 32410 8656 32474
rect 8720 32410 9375 32474
rect 9439 32410 10094 32474
rect 10158 32410 10813 32474
rect 10877 32410 11532 32474
rect 11596 32410 12251 32474
rect 12315 32410 12970 32474
rect 13034 32410 13689 32474
rect 13753 32410 13774 32474
rect 6602 32382 13774 32410
rect 6604 32254 6804 32282
rect 6604 32190 6632 32254
rect 6696 32250 6712 32254
rect 6696 32190 6712 32194
rect 6776 32190 6804 32254
rect 6604 32162 6804 32190
rect 13532 32188 13538 32252
rect 13602 32250 13608 32252
rect 14181 32250 14247 32253
rect 13602 32248 14247 32250
rect 13602 32192 14186 32248
rect 14242 32192 14247 32248
rect 13602 32190 14247 32192
rect 13602 32188 13608 32190
rect 14181 32187 14247 32190
rect 900 32064 2532 32092
rect 900 32000 924 32064
rect 988 32000 1004 32064
rect 1068 32000 1084 32064
rect 1148 32000 1164 32064
rect 1228 32000 1244 32064
rect 1308 32000 1324 32064
rect 1388 32000 1404 32064
rect 1468 32000 1484 32064
rect 1548 32000 1564 32064
rect 1628 32000 1644 32064
rect 1708 32000 1724 32064
rect 1788 32000 1804 32064
rect 1868 32000 1884 32064
rect 1948 32000 1964 32064
rect 2028 32000 2044 32064
rect 2108 32000 2124 32064
rect 2188 32000 2204 32064
rect 2268 32000 2284 32064
rect 2348 32000 2364 32064
rect 2428 32000 2444 32064
rect 2508 32000 2532 32064
rect 900 31972 2532 32000
rect 46104 32064 47736 32092
rect 46104 32000 46128 32064
rect 46192 32000 46208 32064
rect 46272 32000 46288 32064
rect 46352 32000 46368 32064
rect 46432 32000 46448 32064
rect 46512 32000 46528 32064
rect 46592 32000 46608 32064
rect 46672 32000 46688 32064
rect 46752 32000 46768 32064
rect 46832 32000 46848 32064
rect 46912 32000 46928 32064
rect 46992 32000 47008 32064
rect 47072 32000 47088 32064
rect 47152 32000 47168 32064
rect 47232 32000 47248 32064
rect 47312 32000 47328 32064
rect 47392 32000 47408 32064
rect 47472 32000 47488 32064
rect 47552 32000 47568 32064
rect 47632 32000 47648 32064
rect 47712 32000 47736 32064
rect 46104 31972 47736 32000
rect 3348 30184 4980 30212
rect 3348 30120 3372 30184
rect 3436 30120 3452 30184
rect 3516 30120 3532 30184
rect 3596 30120 3612 30184
rect 3676 30120 3692 30184
rect 3756 30120 3772 30184
rect 3836 30120 3852 30184
rect 3916 30120 3932 30184
rect 3996 30120 4012 30184
rect 4076 30120 4092 30184
rect 4156 30120 4172 30184
rect 4236 30120 4252 30184
rect 4316 30120 4332 30184
rect 4396 30120 4412 30184
rect 4476 30120 4492 30184
rect 4556 30120 4572 30184
rect 4636 30120 4652 30184
rect 4716 30120 4732 30184
rect 4796 30120 4812 30184
rect 4876 30120 4892 30184
rect 4956 30120 4980 30184
rect 3348 30092 4980 30120
rect 43656 30184 45288 30212
rect 43656 30120 43680 30184
rect 43744 30120 43760 30184
rect 43824 30120 43840 30184
rect 43904 30120 43920 30184
rect 43984 30120 44000 30184
rect 44064 30120 44080 30184
rect 44144 30120 44160 30184
rect 44224 30120 44240 30184
rect 44304 30120 44320 30184
rect 44384 30120 44400 30184
rect 44464 30120 44480 30184
rect 44544 30120 44560 30184
rect 44624 30120 44640 30184
rect 44704 30120 44720 30184
rect 44784 30120 44800 30184
rect 44864 30120 44880 30184
rect 44944 30120 44960 30184
rect 45024 30120 45040 30184
rect 45104 30120 45120 30184
rect 45184 30120 45200 30184
rect 45264 30120 45288 30184
rect 43656 30092 45288 30120
rect 18873 28592 18939 28593
rect 18873 28590 18920 28592
rect 18830 28588 18920 28590
rect 18830 28532 18878 28588
rect 18830 28530 18920 28532
rect 18873 28528 18920 28530
rect 18984 28528 18990 28592
rect 18873 28527 18939 28528
rect 900 28304 2532 28332
rect 900 28240 924 28304
rect 988 28240 1004 28304
rect 1068 28240 1084 28304
rect 1148 28240 1164 28304
rect 1228 28240 1244 28304
rect 1308 28240 1324 28304
rect 1388 28240 1404 28304
rect 1468 28240 1484 28304
rect 1548 28240 1564 28304
rect 1628 28240 1644 28304
rect 1708 28240 1724 28304
rect 1788 28240 1804 28304
rect 1868 28240 1884 28304
rect 1948 28240 1964 28304
rect 2028 28240 2044 28304
rect 2108 28240 2124 28304
rect 2188 28240 2204 28304
rect 2268 28240 2284 28304
rect 2348 28240 2364 28304
rect 2428 28240 2444 28304
rect 2508 28240 2532 28304
rect 900 28212 2532 28240
rect 46104 28304 47736 28332
rect 46104 28240 46128 28304
rect 46192 28240 46208 28304
rect 46272 28240 46288 28304
rect 46352 28240 46368 28304
rect 46432 28240 46448 28304
rect 46512 28240 46528 28304
rect 46592 28240 46608 28304
rect 46672 28240 46688 28304
rect 46752 28240 46768 28304
rect 46832 28240 46848 28304
rect 46912 28240 46928 28304
rect 46992 28240 47008 28304
rect 47072 28240 47088 28304
rect 47152 28240 47168 28304
rect 47232 28240 47248 28304
rect 47312 28240 47328 28304
rect 47392 28240 47408 28304
rect 47472 28240 47488 28304
rect 47552 28240 47568 28304
rect 47632 28240 47648 28304
rect 47712 28240 47736 28304
rect 46104 28212 47736 28240
rect 3348 26424 4980 26452
rect 3348 26360 3372 26424
rect 3436 26360 3452 26424
rect 3516 26360 3532 26424
rect 3596 26360 3612 26424
rect 3676 26360 3692 26424
rect 3756 26360 3772 26424
rect 3836 26360 3852 26424
rect 3916 26360 3932 26424
rect 3996 26360 4012 26424
rect 4076 26360 4092 26424
rect 4156 26360 4172 26424
rect 4236 26360 4252 26424
rect 4316 26360 4332 26424
rect 4396 26360 4412 26424
rect 4476 26360 4492 26424
rect 4556 26360 4572 26424
rect 4636 26360 4652 26424
rect 4716 26360 4732 26424
rect 4796 26360 4812 26424
rect 4876 26360 4892 26424
rect 4956 26360 4980 26424
rect 3348 26332 4980 26360
rect 43656 26424 45288 26452
rect 43656 26360 43680 26424
rect 43744 26360 43760 26424
rect 43824 26360 43840 26424
rect 43904 26360 43920 26424
rect 43984 26360 44000 26424
rect 44064 26360 44080 26424
rect 44144 26360 44160 26424
rect 44224 26360 44240 26424
rect 44304 26360 44320 26424
rect 44384 26360 44400 26424
rect 44464 26360 44480 26424
rect 44544 26360 44560 26424
rect 44624 26360 44640 26424
rect 44704 26360 44720 26424
rect 44784 26360 44800 26424
rect 44864 26360 44880 26424
rect 44944 26360 44960 26424
rect 45024 26360 45040 26424
rect 45104 26360 45120 26424
rect 45184 26360 45200 26424
rect 45264 26360 45288 26424
rect 43656 26332 45288 26360
rect 15422 26150 22594 26162
rect 15422 26094 15454 26150
rect 15510 26094 15534 26150
rect 15590 26134 22594 26150
rect 15590 26094 16038 26134
rect 15422 26070 16038 26094
rect 16102 26070 16757 26134
rect 16821 26070 17476 26134
rect 17540 26070 18195 26134
rect 18259 26070 18914 26134
rect 18978 26070 19633 26134
rect 19697 26070 20352 26134
rect 20416 26070 21071 26134
rect 21135 26070 21790 26134
rect 21854 26070 22509 26134
rect 22573 26070 22594 26134
rect 15422 26054 22594 26070
rect 15422 25990 16038 26054
rect 16102 25990 16757 26054
rect 16821 25990 17476 26054
rect 17540 25990 18195 26054
rect 18259 25990 18914 26054
rect 18978 25990 19633 26054
rect 19697 25990 20352 26054
rect 20416 25990 21071 26054
rect 21135 25990 21790 26054
rect 21854 25990 22509 26054
rect 22573 25990 22594 26054
rect 15422 25974 22594 25990
rect 15422 25910 16038 25974
rect 16102 25910 16757 25974
rect 16821 25910 17476 25974
rect 17540 25910 18195 25974
rect 18259 25910 18914 25974
rect 18978 25910 19633 25974
rect 19697 25910 20352 25974
rect 20416 25910 21071 25974
rect 21135 25910 21790 25974
rect 21854 25910 22509 25974
rect 22573 25910 22594 25974
rect 15422 25894 22594 25910
rect 15422 25830 16038 25894
rect 16102 25830 16757 25894
rect 16821 25830 17476 25894
rect 17540 25830 18195 25894
rect 18259 25830 18914 25894
rect 18978 25830 19633 25894
rect 19697 25830 20352 25894
rect 20416 25830 21071 25894
rect 21135 25830 21790 25894
rect 21854 25830 22509 25894
rect 22573 25830 22594 25894
rect 15422 25814 22594 25830
rect 15422 25750 16038 25814
rect 16102 25750 16757 25814
rect 16821 25750 17476 25814
rect 17540 25750 18195 25814
rect 18259 25750 18914 25814
rect 18978 25750 19633 25814
rect 19697 25750 20352 25814
rect 20416 25750 21071 25814
rect 21135 25750 21790 25814
rect 21854 25750 22509 25814
rect 22573 25750 22594 25814
rect 15422 25734 22594 25750
rect 15422 25670 16038 25734
rect 16102 25670 16757 25734
rect 16821 25670 17476 25734
rect 17540 25670 18195 25734
rect 18259 25670 18914 25734
rect 18978 25670 19633 25734
rect 19697 25670 20352 25734
rect 20416 25670 21071 25734
rect 21135 25670 21790 25734
rect 21854 25670 22509 25734
rect 22573 25670 22594 25734
rect 15422 25654 22594 25670
rect 15422 25590 16038 25654
rect 16102 25590 16757 25654
rect 16821 25590 17476 25654
rect 17540 25590 18195 25654
rect 18259 25590 18914 25654
rect 18978 25590 19633 25654
rect 19697 25590 20352 25654
rect 20416 25590 21071 25654
rect 21135 25590 21790 25654
rect 21854 25590 22509 25654
rect 22573 25590 22594 25654
rect 15422 25434 22594 25590
rect 15422 25370 16038 25434
rect 16102 25370 16757 25434
rect 16821 25370 17476 25434
rect 17540 25370 18195 25434
rect 18259 25370 18914 25434
rect 18978 25370 19633 25434
rect 19697 25370 20352 25434
rect 20416 25370 21071 25434
rect 21135 25370 21790 25434
rect 21854 25370 22509 25434
rect 22573 25370 22594 25434
rect 15422 25354 22594 25370
rect 15422 25290 16038 25354
rect 16102 25290 16757 25354
rect 16821 25290 17476 25354
rect 17540 25290 18195 25354
rect 18259 25290 18914 25354
rect 18978 25290 19633 25354
rect 19697 25290 20352 25354
rect 20416 25290 21071 25354
rect 21135 25290 21790 25354
rect 21854 25290 22509 25354
rect 22573 25290 22594 25354
rect 15422 25274 22594 25290
rect 15422 25210 16038 25274
rect 16102 25210 16757 25274
rect 16821 25210 17476 25274
rect 17540 25210 18195 25274
rect 18259 25210 18914 25274
rect 18978 25210 19633 25274
rect 19697 25210 20352 25274
rect 20416 25210 21071 25274
rect 21135 25210 21790 25274
rect 21854 25210 22509 25274
rect 22573 25210 22594 25274
rect 15422 25194 22594 25210
rect 15422 25130 16038 25194
rect 16102 25130 16757 25194
rect 16821 25130 17476 25194
rect 17540 25130 18195 25194
rect 18259 25130 18914 25194
rect 18978 25130 19633 25194
rect 19697 25130 20352 25194
rect 20416 25130 21071 25194
rect 21135 25130 21790 25194
rect 21854 25130 22509 25194
rect 22573 25130 22594 25194
rect 15422 25114 22594 25130
rect 15422 25050 16038 25114
rect 16102 25050 16757 25114
rect 16821 25050 17476 25114
rect 17540 25050 18195 25114
rect 18259 25050 18914 25114
rect 18978 25050 19633 25114
rect 19697 25050 20352 25114
rect 20416 25050 21071 25114
rect 21135 25050 21790 25114
rect 21854 25050 22509 25114
rect 22573 25050 22594 25114
rect 15422 25034 22594 25050
rect 15422 24970 16038 25034
rect 16102 24970 16757 25034
rect 16821 24970 17476 25034
rect 17540 24970 18195 25034
rect 18259 24970 18914 25034
rect 18978 24970 19633 25034
rect 19697 24970 20352 25034
rect 20416 24970 21071 25034
rect 21135 24970 21790 25034
rect 21854 24970 22509 25034
rect 22573 24970 22594 25034
rect 22778 24990 22784 25054
rect 22848 25052 22854 25054
rect 23289 25052 23355 25055
rect 22848 25050 23355 25052
rect 22848 24994 23294 25050
rect 23350 24994 23355 25050
rect 22848 24992 23355 24994
rect 22848 24990 22854 24992
rect 23289 24989 23355 24992
rect 15422 24954 22594 24970
rect 15422 24890 16038 24954
rect 16102 24890 16757 24954
rect 16821 24890 17476 24954
rect 17540 24890 18195 24954
rect 18259 24890 18914 24954
rect 18978 24890 19633 24954
rect 19697 24890 20352 24954
rect 20416 24890 21071 24954
rect 21135 24890 21790 24954
rect 21854 24890 22509 24954
rect 22573 24890 22594 24954
rect 15422 24862 22594 24890
rect 15424 24734 15624 24762
rect 15424 24670 15452 24734
rect 15516 24730 15532 24734
rect 15516 24670 15532 24674
rect 15596 24670 15624 24734
rect 15424 24642 15624 24670
rect 900 24544 2532 24572
rect 15469 24566 15535 24567
rect 15464 24564 15470 24566
rect 900 24480 924 24544
rect 988 24480 1004 24544
rect 1068 24480 1084 24544
rect 1148 24480 1164 24544
rect 1228 24480 1244 24544
rect 1308 24480 1324 24544
rect 1388 24480 1404 24544
rect 1468 24480 1484 24544
rect 1548 24480 1564 24544
rect 1628 24480 1644 24544
rect 1708 24480 1724 24544
rect 1788 24480 1804 24544
rect 1868 24480 1884 24544
rect 1948 24480 1964 24544
rect 2028 24480 2044 24544
rect 2108 24480 2124 24544
rect 2188 24480 2204 24544
rect 2268 24480 2284 24544
rect 2348 24480 2364 24544
rect 2428 24480 2444 24544
rect 2508 24480 2532 24544
rect 15380 24504 15470 24564
rect 15464 24502 15470 24504
rect 15534 24502 15540 24566
rect 46104 24544 47736 24572
rect 15469 24501 15535 24502
rect 900 24452 2532 24480
rect 46104 24480 46128 24544
rect 46192 24480 46208 24544
rect 46272 24480 46288 24544
rect 46352 24480 46368 24544
rect 46432 24480 46448 24544
rect 46512 24480 46528 24544
rect 46592 24480 46608 24544
rect 46672 24480 46688 24544
rect 46752 24480 46768 24544
rect 46832 24480 46848 24544
rect 46912 24480 46928 24544
rect 46992 24480 47008 24544
rect 47072 24480 47088 24544
rect 47152 24480 47168 24544
rect 47232 24480 47248 24544
rect 47312 24480 47328 24544
rect 47392 24480 47408 24544
rect 47472 24480 47488 24544
rect 47552 24480 47568 24544
rect 47632 24480 47648 24544
rect 47712 24480 47736 24544
rect 46104 24452 47736 24480
rect 3348 22664 4980 22692
rect 3348 22600 3372 22664
rect 3436 22600 3452 22664
rect 3516 22600 3532 22664
rect 3596 22600 3612 22664
rect 3676 22600 3692 22664
rect 3756 22600 3772 22664
rect 3836 22600 3852 22664
rect 3916 22600 3932 22664
rect 3996 22600 4012 22664
rect 4076 22600 4092 22664
rect 4156 22600 4172 22664
rect 4236 22600 4252 22664
rect 4316 22600 4332 22664
rect 4396 22600 4412 22664
rect 4476 22600 4492 22664
rect 4556 22600 4572 22664
rect 4636 22600 4652 22664
rect 4716 22600 4732 22664
rect 4796 22600 4812 22664
rect 4876 22600 4892 22664
rect 4956 22600 4980 22664
rect 43656 22664 45288 22692
rect 3348 22572 4980 22600
rect 13261 22612 13327 22615
rect 14222 22612 14228 22614
rect 13261 22610 14228 22612
rect 13261 22554 13266 22610
rect 13322 22554 14228 22610
rect 13261 22552 14228 22554
rect 13261 22549 13327 22552
rect 14222 22550 14228 22552
rect 14292 22550 14298 22614
rect 43656 22600 43680 22664
rect 43744 22600 43760 22664
rect 43824 22600 43840 22664
rect 43904 22600 43920 22664
rect 43984 22600 44000 22664
rect 44064 22600 44080 22664
rect 44144 22600 44160 22664
rect 44224 22600 44240 22664
rect 44304 22600 44320 22664
rect 44384 22600 44400 22664
rect 44464 22600 44480 22664
rect 44544 22600 44560 22664
rect 44624 22600 44640 22664
rect 44704 22600 44720 22664
rect 44784 22600 44800 22664
rect 44864 22600 44880 22664
rect 44944 22600 44960 22664
rect 45024 22600 45040 22664
rect 45104 22600 45120 22664
rect 45184 22600 45200 22664
rect 45264 22600 45288 22664
rect 43656 22572 45288 22600
rect 13560 22390 20732 22402
rect 13560 22334 13592 22390
rect 13648 22334 13672 22390
rect 13728 22374 20732 22390
rect 13728 22334 14176 22374
rect 13560 22310 14176 22334
rect 14240 22310 14895 22374
rect 14959 22310 15614 22374
rect 15678 22310 16333 22374
rect 16397 22310 17052 22374
rect 17116 22310 17771 22374
rect 17835 22310 18490 22374
rect 18554 22310 19209 22374
rect 19273 22310 19928 22374
rect 19992 22310 20647 22374
rect 20711 22310 20732 22374
rect 13560 22294 20732 22310
rect 13560 22230 14176 22294
rect 14240 22230 14895 22294
rect 14959 22230 15614 22294
rect 15678 22230 16333 22294
rect 16397 22230 17052 22294
rect 17116 22230 17771 22294
rect 17835 22230 18490 22294
rect 18554 22230 19209 22294
rect 19273 22230 19928 22294
rect 19992 22230 20647 22294
rect 20711 22230 20732 22294
rect 13560 22214 20732 22230
rect 13560 22150 14176 22214
rect 14240 22150 14895 22214
rect 14959 22150 15614 22214
rect 15678 22150 16333 22214
rect 16397 22150 17052 22214
rect 17116 22150 17771 22214
rect 17835 22150 18490 22214
rect 18554 22150 19209 22214
rect 19273 22150 19928 22214
rect 19992 22150 20647 22214
rect 20711 22150 20732 22214
rect 13560 22134 20732 22150
rect 13560 22070 14176 22134
rect 14240 22070 14895 22134
rect 14959 22070 15614 22134
rect 15678 22070 16333 22134
rect 16397 22070 17052 22134
rect 17116 22070 17771 22134
rect 17835 22070 18490 22134
rect 18554 22070 19209 22134
rect 19273 22070 19928 22134
rect 19992 22070 20647 22134
rect 20711 22070 20732 22134
rect 13560 22054 20732 22070
rect 13560 21990 14176 22054
rect 14240 21990 14895 22054
rect 14959 21990 15614 22054
rect 15678 21990 16333 22054
rect 16397 21990 17052 22054
rect 17116 21990 17771 22054
rect 17835 21990 18490 22054
rect 18554 21990 19209 22054
rect 19273 21990 19928 22054
rect 19992 21990 20647 22054
rect 20711 21990 20732 22054
rect 13560 21974 20732 21990
rect 13560 21910 14176 21974
rect 14240 21910 14895 21974
rect 14959 21910 15614 21974
rect 15678 21910 16333 21974
rect 16397 21910 17052 21974
rect 17116 21910 17771 21974
rect 17835 21910 18490 21974
rect 18554 21910 19209 21974
rect 19273 21910 19928 21974
rect 19992 21910 20647 21974
rect 20711 21910 20732 21974
rect 13560 21894 20732 21910
rect 13560 21830 14176 21894
rect 14240 21830 14895 21894
rect 14959 21830 15614 21894
rect 15678 21830 16333 21894
rect 16397 21830 17052 21894
rect 17116 21830 17771 21894
rect 17835 21830 18490 21894
rect 18554 21830 19209 21894
rect 19273 21830 19928 21894
rect 19992 21830 20647 21894
rect 20711 21830 20732 21894
rect 13560 21674 20732 21830
rect 13560 21610 14176 21674
rect 14240 21610 14895 21674
rect 14959 21610 15614 21674
rect 15678 21610 16333 21674
rect 16397 21610 17052 21674
rect 17116 21610 17771 21674
rect 17835 21610 18490 21674
rect 18554 21610 19209 21674
rect 19273 21610 19928 21674
rect 19992 21610 20647 21674
rect 20711 21610 20732 21674
rect 20897 21638 20963 21639
rect 13560 21594 20732 21610
rect 13560 21530 14176 21594
rect 14240 21530 14895 21594
rect 14959 21530 15614 21594
rect 15678 21530 16333 21594
rect 16397 21530 17052 21594
rect 17116 21530 17771 21594
rect 17835 21530 18490 21594
rect 18554 21530 19209 21594
rect 19273 21530 19928 21594
rect 19992 21530 20647 21594
rect 20711 21530 20732 21594
rect 20846 21574 20852 21638
rect 20916 21636 20963 21638
rect 20916 21634 21006 21636
rect 20958 21578 21006 21634
rect 20916 21576 21006 21578
rect 20916 21574 20963 21576
rect 20897 21573 20963 21574
rect 13560 21514 20732 21530
rect 13560 21450 14176 21514
rect 14240 21450 14895 21514
rect 14959 21450 15614 21514
rect 15678 21450 16333 21514
rect 16397 21450 17052 21514
rect 17116 21450 17771 21514
rect 17835 21450 18490 21514
rect 18554 21450 19209 21514
rect 19273 21450 19928 21514
rect 19992 21450 20647 21514
rect 20711 21450 20732 21514
rect 13560 21434 20732 21450
rect 13560 21370 14176 21434
rect 14240 21370 14895 21434
rect 14959 21370 15614 21434
rect 15678 21370 16333 21434
rect 16397 21370 17052 21434
rect 17116 21370 17771 21434
rect 17835 21370 18490 21434
rect 18554 21370 19209 21434
rect 19273 21370 19928 21434
rect 19992 21370 20647 21434
rect 20711 21370 20732 21434
rect 13560 21354 20732 21370
rect 13560 21290 14176 21354
rect 14240 21290 14895 21354
rect 14959 21290 15614 21354
rect 15678 21290 16333 21354
rect 16397 21290 17052 21354
rect 17116 21290 17771 21354
rect 17835 21290 18490 21354
rect 18554 21290 19209 21354
rect 19273 21290 19928 21354
rect 19992 21290 20647 21354
rect 20711 21290 20732 21354
rect 13560 21274 20732 21290
rect 13560 21210 14176 21274
rect 14240 21210 14895 21274
rect 14959 21210 15614 21274
rect 15678 21210 16333 21274
rect 16397 21210 17052 21274
rect 17116 21210 17771 21274
rect 17835 21210 18490 21274
rect 18554 21210 19209 21274
rect 19273 21210 19928 21274
rect 19992 21210 20647 21274
rect 20711 21210 20732 21274
rect 13560 21194 20732 21210
rect 13560 21130 14176 21194
rect 14240 21130 14895 21194
rect 14959 21130 15614 21194
rect 15678 21130 16333 21194
rect 16397 21130 17052 21194
rect 17116 21130 17771 21194
rect 17835 21130 18490 21194
rect 18554 21130 19209 21194
rect 19273 21130 19928 21194
rect 19992 21130 20647 21194
rect 20711 21130 20732 21194
rect 13560 21102 20732 21130
rect 13562 20974 13762 21002
rect 13562 20910 13590 20974
rect 13654 20970 13670 20974
rect 13654 20910 13670 20914
rect 13734 20910 13762 20974
rect 13562 20882 13762 20910
rect 14089 20906 14155 20907
rect 14084 20904 14090 20906
rect 14000 20844 14090 20904
rect 14084 20842 14090 20844
rect 14154 20842 14160 20906
rect 14089 20841 14155 20842
rect 900 20784 2532 20812
rect 900 20720 924 20784
rect 988 20720 1004 20784
rect 1068 20720 1084 20784
rect 1148 20720 1164 20784
rect 1228 20720 1244 20784
rect 1308 20720 1324 20784
rect 1388 20720 1404 20784
rect 1468 20720 1484 20784
rect 1548 20720 1564 20784
rect 1628 20720 1644 20784
rect 1708 20720 1724 20784
rect 1788 20720 1804 20784
rect 1868 20720 1884 20784
rect 1948 20720 1964 20784
rect 2028 20720 2044 20784
rect 2108 20720 2124 20784
rect 2188 20720 2204 20784
rect 2268 20720 2284 20784
rect 2348 20720 2364 20784
rect 2428 20720 2444 20784
rect 2508 20720 2532 20784
rect 900 20692 2532 20720
rect 46104 20784 47736 20812
rect 46104 20720 46128 20784
rect 46192 20720 46208 20784
rect 46272 20720 46288 20784
rect 46352 20720 46368 20784
rect 46432 20720 46448 20784
rect 46512 20720 46528 20784
rect 46592 20720 46608 20784
rect 46672 20720 46688 20784
rect 46752 20720 46768 20784
rect 46832 20720 46848 20784
rect 46912 20720 46928 20784
rect 46992 20720 47008 20784
rect 47072 20720 47088 20784
rect 47152 20720 47168 20784
rect 47232 20720 47248 20784
rect 47312 20720 47328 20784
rect 47392 20720 47408 20784
rect 47472 20720 47488 20784
rect 47552 20720 47568 20784
rect 47632 20720 47648 20784
rect 47712 20720 47736 20784
rect 46104 20692 47736 20720
rect 20713 18952 20779 18955
rect 20984 18952 20990 18954
rect 20713 18950 20990 18952
rect 3348 18904 4980 18932
rect 3348 18840 3372 18904
rect 3436 18840 3452 18904
rect 3516 18840 3532 18904
rect 3596 18840 3612 18904
rect 3676 18840 3692 18904
rect 3756 18840 3772 18904
rect 3836 18840 3852 18904
rect 3916 18840 3932 18904
rect 3996 18840 4012 18904
rect 4076 18840 4092 18904
rect 4156 18840 4172 18904
rect 4236 18840 4252 18904
rect 4316 18840 4332 18904
rect 4396 18840 4412 18904
rect 4476 18840 4492 18904
rect 4556 18840 4572 18904
rect 4636 18840 4652 18904
rect 4716 18840 4732 18904
rect 4796 18840 4812 18904
rect 4876 18840 4892 18904
rect 4956 18840 4980 18904
rect 20713 18894 20718 18950
rect 20774 18894 20990 18950
rect 20713 18892 20990 18894
rect 20713 18889 20779 18892
rect 20984 18890 20990 18892
rect 21054 18890 21060 18954
rect 43656 18904 45288 18932
rect 3348 18812 4980 18840
rect 43656 18840 43680 18904
rect 43744 18840 43760 18904
rect 43824 18840 43840 18904
rect 43904 18840 43920 18904
rect 43984 18840 44000 18904
rect 44064 18840 44080 18904
rect 44144 18840 44160 18904
rect 44224 18840 44240 18904
rect 44304 18840 44320 18904
rect 44384 18840 44400 18904
rect 44464 18840 44480 18904
rect 44544 18840 44560 18904
rect 44624 18840 44640 18904
rect 44704 18840 44720 18904
rect 44784 18840 44800 18904
rect 44864 18840 44880 18904
rect 44944 18840 44960 18904
rect 45024 18840 45040 18904
rect 45104 18840 45120 18904
rect 45184 18840 45200 18904
rect 45264 18840 45288 18904
rect 43656 18812 45288 18840
rect 16108 18630 23280 18642
rect 16108 18574 16140 18630
rect 16196 18574 16220 18630
rect 16276 18614 23280 18630
rect 16276 18574 16724 18614
rect 16108 18550 16724 18574
rect 16788 18550 17443 18614
rect 17507 18550 18162 18614
rect 18226 18550 18881 18614
rect 18945 18550 19600 18614
rect 19664 18550 20319 18614
rect 20383 18550 21038 18614
rect 21102 18550 21757 18614
rect 21821 18550 22476 18614
rect 22540 18550 23195 18614
rect 23259 18550 23280 18614
rect 16108 18534 23280 18550
rect 16108 18470 16724 18534
rect 16788 18470 17443 18534
rect 17507 18470 18162 18534
rect 18226 18470 18881 18534
rect 18945 18470 19600 18534
rect 19664 18470 20319 18534
rect 20383 18470 21038 18534
rect 21102 18470 21757 18534
rect 21821 18470 22476 18534
rect 22540 18470 23195 18534
rect 23259 18470 23280 18534
rect 16108 18454 23280 18470
rect 16108 18390 16724 18454
rect 16788 18390 17443 18454
rect 17507 18390 18162 18454
rect 18226 18390 18881 18454
rect 18945 18390 19600 18454
rect 19664 18390 20319 18454
rect 20383 18390 21038 18454
rect 21102 18390 21757 18454
rect 21821 18390 22476 18454
rect 22540 18390 23195 18454
rect 23259 18390 23280 18454
rect 16108 18374 23280 18390
rect 16108 18310 16724 18374
rect 16788 18310 17443 18374
rect 17507 18310 18162 18374
rect 18226 18310 18881 18374
rect 18945 18310 19600 18374
rect 19664 18310 20319 18374
rect 20383 18310 21038 18374
rect 21102 18310 21757 18374
rect 21821 18310 22476 18374
rect 22540 18310 23195 18374
rect 23259 18310 23280 18374
rect 16108 18294 23280 18310
rect 16108 18230 16724 18294
rect 16788 18230 17443 18294
rect 17507 18230 18162 18294
rect 18226 18230 18881 18294
rect 18945 18230 19600 18294
rect 19664 18230 20319 18294
rect 20383 18230 21038 18294
rect 21102 18230 21757 18294
rect 21821 18230 22476 18294
rect 22540 18230 23195 18294
rect 23259 18230 23280 18294
rect 16108 18214 23280 18230
rect 16108 18150 16724 18214
rect 16788 18150 17443 18214
rect 17507 18150 18162 18214
rect 18226 18150 18881 18214
rect 18945 18150 19600 18214
rect 19664 18150 20319 18214
rect 20383 18150 21038 18214
rect 21102 18150 21757 18214
rect 21821 18150 22476 18214
rect 22540 18150 23195 18214
rect 23259 18150 23280 18214
rect 16108 18134 23280 18150
rect 16108 18070 16724 18134
rect 16788 18070 17443 18134
rect 17507 18070 18162 18134
rect 18226 18070 18881 18134
rect 18945 18070 19600 18134
rect 19664 18070 20319 18134
rect 20383 18070 21038 18134
rect 21102 18070 21757 18134
rect 21821 18070 22476 18134
rect 22540 18070 23195 18134
rect 23259 18070 23280 18134
rect 16108 17914 23280 18070
rect 16108 17850 16724 17914
rect 16788 17850 17443 17914
rect 17507 17850 18162 17914
rect 18226 17850 18881 17914
rect 18945 17850 19600 17914
rect 19664 17850 20319 17914
rect 20383 17850 21038 17914
rect 21102 17850 21757 17914
rect 21821 17850 22476 17914
rect 22540 17850 23195 17914
rect 23259 17850 23280 17914
rect 16108 17834 23280 17850
rect 16108 17770 16724 17834
rect 16788 17770 17443 17834
rect 17507 17770 18162 17834
rect 18226 17770 18881 17834
rect 18945 17770 19600 17834
rect 19664 17770 20319 17834
rect 20383 17770 21038 17834
rect 21102 17770 21757 17834
rect 21821 17770 22476 17834
rect 22540 17770 23195 17834
rect 23259 17770 23280 17834
rect 16108 17754 23280 17770
rect 16108 17690 16724 17754
rect 16788 17690 17443 17754
rect 17507 17690 18162 17754
rect 18226 17690 18881 17754
rect 18945 17690 19600 17754
rect 19664 17690 20319 17754
rect 20383 17690 21038 17754
rect 21102 17690 21757 17754
rect 21821 17690 22476 17754
rect 22540 17690 23195 17754
rect 23259 17690 23280 17754
rect 16108 17674 23280 17690
rect 16108 17610 16724 17674
rect 16788 17610 17443 17674
rect 17507 17610 18162 17674
rect 18226 17610 18881 17674
rect 18945 17610 19600 17674
rect 19664 17610 20319 17674
rect 20383 17610 21038 17674
rect 21102 17610 21757 17674
rect 21821 17610 22476 17674
rect 22540 17610 23195 17674
rect 23259 17610 23280 17674
rect 16108 17594 23280 17610
rect 16108 17530 16724 17594
rect 16788 17530 17443 17594
rect 17507 17530 18162 17594
rect 18226 17530 18881 17594
rect 18945 17530 19600 17594
rect 19664 17530 20319 17594
rect 20383 17530 21038 17594
rect 21102 17530 21757 17594
rect 21821 17530 22476 17594
rect 22540 17530 23195 17594
rect 23259 17530 23280 17594
rect 16108 17514 23280 17530
rect 16108 17450 16724 17514
rect 16788 17450 17443 17514
rect 17507 17450 18162 17514
rect 18226 17450 18881 17514
rect 18945 17450 19600 17514
rect 19664 17450 20319 17514
rect 20383 17450 21038 17514
rect 21102 17450 21757 17514
rect 21821 17450 22476 17514
rect 22540 17450 23195 17514
rect 23259 17450 23280 17514
rect 16108 17434 23280 17450
rect 16108 17370 16724 17434
rect 16788 17370 17443 17434
rect 17507 17370 18162 17434
rect 18226 17370 18881 17434
rect 18945 17370 19600 17434
rect 19664 17370 20319 17434
rect 20383 17370 21038 17434
rect 21102 17370 21757 17434
rect 21821 17370 22476 17434
rect 22540 17370 23195 17434
rect 23259 17370 23280 17434
rect 16108 17342 23280 17370
rect 16110 17214 16310 17242
rect 16110 17150 16138 17214
rect 16202 17210 16218 17214
rect 16202 17150 16218 17154
rect 16282 17150 16310 17214
rect 16110 17122 16310 17150
rect 900 17024 2532 17052
rect 900 16960 924 17024
rect 988 16960 1004 17024
rect 1068 16960 1084 17024
rect 1148 16960 1164 17024
rect 1228 16960 1244 17024
rect 1308 16960 1324 17024
rect 1388 16960 1404 17024
rect 1468 16960 1484 17024
rect 1548 16960 1564 17024
rect 1628 16960 1644 17024
rect 1708 16960 1724 17024
rect 1788 16960 1804 17024
rect 1868 16960 1884 17024
rect 1948 16960 1964 17024
rect 2028 16960 2044 17024
rect 2108 16960 2124 17024
rect 2188 16960 2204 17024
rect 2268 16960 2284 17024
rect 2348 16960 2364 17024
rect 2428 16960 2444 17024
rect 2508 16960 2532 17024
rect 46104 17024 47736 17052
rect 17401 17002 17467 17003
rect 17396 17000 17402 17002
rect 900 16932 2532 16960
rect 17312 16940 17402 17000
rect 17396 16938 17402 16940
rect 17466 16938 17472 17002
rect 46104 16960 46128 17024
rect 46192 16960 46208 17024
rect 46272 16960 46288 17024
rect 46352 16960 46368 17024
rect 46432 16960 46448 17024
rect 46512 16960 46528 17024
rect 46592 16960 46608 17024
rect 46672 16960 46688 17024
rect 46752 16960 46768 17024
rect 46832 16960 46848 17024
rect 46912 16960 46928 17024
rect 46992 16960 47008 17024
rect 47072 16960 47088 17024
rect 47152 16960 47168 17024
rect 47232 16960 47248 17024
rect 47312 16960 47328 17024
rect 47392 16960 47408 17024
rect 47472 16960 47488 17024
rect 47552 16960 47568 17024
rect 47632 16960 47648 17024
rect 47712 16960 47736 17024
rect 17401 16937 17467 16938
rect 46104 16932 47736 16960
rect 19604 16328 19610 16392
rect 19674 16390 19680 16392
rect 20713 16390 20779 16393
rect 19674 16388 20779 16390
rect 19674 16332 20718 16388
rect 20774 16332 20779 16388
rect 19674 16330 20779 16332
rect 19674 16328 19680 16330
rect 20713 16327 20779 16330
rect 3348 15144 4980 15172
rect 3348 15080 3372 15144
rect 3436 15080 3452 15144
rect 3516 15080 3532 15144
rect 3596 15080 3612 15144
rect 3676 15080 3692 15144
rect 3756 15080 3772 15144
rect 3836 15080 3852 15144
rect 3916 15080 3932 15144
rect 3996 15080 4012 15144
rect 4076 15080 4092 15144
rect 4156 15080 4172 15144
rect 4236 15080 4252 15144
rect 4316 15080 4332 15144
rect 4396 15080 4412 15144
rect 4476 15080 4492 15144
rect 4556 15080 4572 15144
rect 4636 15080 4652 15144
rect 4716 15080 4732 15144
rect 4796 15080 4812 15144
rect 4876 15080 4892 15144
rect 4956 15080 4980 15144
rect 3348 15052 4980 15080
rect 43656 15144 45288 15172
rect 43656 15080 43680 15144
rect 43744 15080 43760 15144
rect 43824 15080 43840 15144
rect 43904 15080 43920 15144
rect 43984 15080 44000 15144
rect 44064 15080 44080 15144
rect 44144 15080 44160 15144
rect 44224 15080 44240 15144
rect 44304 15080 44320 15144
rect 44384 15080 44400 15144
rect 44464 15080 44480 15144
rect 44544 15080 44560 15144
rect 44624 15080 44640 15144
rect 44704 15080 44720 15144
rect 44784 15080 44800 15144
rect 44864 15080 44880 15144
rect 44944 15080 44960 15144
rect 45024 15080 45040 15144
rect 45104 15080 45120 15144
rect 45184 15080 45200 15144
rect 45264 15080 45288 15144
rect 43656 15052 45288 15080
rect 16108 14870 23280 14882
rect 16108 14814 16140 14870
rect 16196 14814 16220 14870
rect 16276 14854 23280 14870
rect 16276 14814 16724 14854
rect 16108 14790 16724 14814
rect 16788 14790 17443 14854
rect 17507 14790 18162 14854
rect 18226 14790 18881 14854
rect 18945 14790 19600 14854
rect 19664 14790 20319 14854
rect 20383 14790 21038 14854
rect 21102 14790 21757 14854
rect 21821 14790 22476 14854
rect 22540 14790 23195 14854
rect 23259 14790 23280 14854
rect 16108 14774 23280 14790
rect 16108 14710 16724 14774
rect 16788 14710 17443 14774
rect 17507 14710 18162 14774
rect 18226 14710 18881 14774
rect 18945 14710 19600 14774
rect 19664 14710 20319 14774
rect 20383 14710 21038 14774
rect 21102 14710 21757 14774
rect 21821 14710 22476 14774
rect 22540 14710 23195 14774
rect 23259 14710 23280 14774
rect 16108 14694 23280 14710
rect 16108 14630 16724 14694
rect 16788 14630 17443 14694
rect 17507 14630 18162 14694
rect 18226 14630 18881 14694
rect 18945 14630 19600 14694
rect 19664 14630 20319 14694
rect 20383 14630 21038 14694
rect 21102 14630 21757 14694
rect 21821 14630 22476 14694
rect 22540 14630 23195 14694
rect 23259 14630 23280 14694
rect 16108 14614 23280 14630
rect 16108 14550 16724 14614
rect 16788 14550 17443 14614
rect 17507 14550 18162 14614
rect 18226 14550 18881 14614
rect 18945 14550 19600 14614
rect 19664 14550 20319 14614
rect 20383 14550 21038 14614
rect 21102 14550 21757 14614
rect 21821 14550 22476 14614
rect 22540 14550 23195 14614
rect 23259 14550 23280 14614
rect 16108 14534 23280 14550
rect 16108 14470 16724 14534
rect 16788 14470 17443 14534
rect 17507 14470 18162 14534
rect 18226 14470 18881 14534
rect 18945 14470 19600 14534
rect 19664 14470 20319 14534
rect 20383 14470 21038 14534
rect 21102 14470 21757 14534
rect 21821 14470 22476 14534
rect 22540 14470 23195 14534
rect 23259 14470 23280 14534
rect 16108 14454 23280 14470
rect 16108 14390 16724 14454
rect 16788 14390 17443 14454
rect 17507 14390 18162 14454
rect 18226 14390 18881 14454
rect 18945 14390 19600 14454
rect 19664 14390 20319 14454
rect 20383 14390 21038 14454
rect 21102 14390 21757 14454
rect 21821 14390 22476 14454
rect 22540 14390 23195 14454
rect 23259 14390 23280 14454
rect 16108 14374 23280 14390
rect 16108 14310 16724 14374
rect 16788 14310 17443 14374
rect 17507 14310 18162 14374
rect 18226 14310 18881 14374
rect 18945 14310 19600 14374
rect 19664 14310 20319 14374
rect 20383 14310 21038 14374
rect 21102 14310 21757 14374
rect 21821 14310 22476 14374
rect 22540 14310 23195 14374
rect 23259 14310 23280 14374
rect 16108 14154 23280 14310
rect 16108 14090 16724 14154
rect 16788 14090 17443 14154
rect 17507 14090 18162 14154
rect 18226 14090 18881 14154
rect 18945 14090 19600 14154
rect 19664 14090 20319 14154
rect 20383 14090 21038 14154
rect 21102 14090 21757 14154
rect 21821 14090 22476 14154
rect 22540 14090 23195 14154
rect 23259 14090 23280 14154
rect 16108 14074 23280 14090
rect 16108 14010 16724 14074
rect 16788 14010 17443 14074
rect 17507 14010 18162 14074
rect 18226 14010 18881 14074
rect 18945 14010 19600 14074
rect 19664 14010 20319 14074
rect 20383 14010 21038 14074
rect 21102 14010 21757 14074
rect 21821 14010 22476 14074
rect 22540 14010 23195 14074
rect 23259 14010 23280 14074
rect 16108 13994 23280 14010
rect 16108 13930 16724 13994
rect 16788 13930 17443 13994
rect 17507 13930 18162 13994
rect 18226 13930 18881 13994
rect 18945 13930 19600 13994
rect 19664 13930 20319 13994
rect 20383 13930 21038 13994
rect 21102 13930 21757 13994
rect 21821 13930 22476 13994
rect 22540 13930 23195 13994
rect 23259 13930 23280 13994
rect 16108 13914 23280 13930
rect 16108 13850 16724 13914
rect 16788 13850 17443 13914
rect 17507 13850 18162 13914
rect 18226 13850 18881 13914
rect 18945 13850 19600 13914
rect 19664 13850 20319 13914
rect 20383 13850 21038 13914
rect 21102 13850 21757 13914
rect 21821 13850 22476 13914
rect 22540 13850 23195 13914
rect 23259 13850 23280 13914
rect 16108 13834 23280 13850
rect 16108 13770 16724 13834
rect 16788 13770 17443 13834
rect 17507 13770 18162 13834
rect 18226 13770 18881 13834
rect 18945 13770 19600 13834
rect 19664 13770 20319 13834
rect 20383 13770 21038 13834
rect 21102 13770 21757 13834
rect 21821 13770 22476 13834
rect 22540 13770 23195 13834
rect 23259 13770 23280 13834
rect 16108 13754 23280 13770
rect 16108 13690 16724 13754
rect 16788 13690 17443 13754
rect 17507 13690 18162 13754
rect 18226 13690 18881 13754
rect 18945 13690 19600 13754
rect 19664 13690 20319 13754
rect 20383 13690 21038 13754
rect 21102 13690 21757 13754
rect 21821 13690 22476 13754
rect 22540 13690 23195 13754
rect 23259 13690 23280 13754
rect 16108 13674 23280 13690
rect 16108 13610 16724 13674
rect 16788 13610 17443 13674
rect 17507 13610 18162 13674
rect 18226 13610 18881 13674
rect 18945 13610 19600 13674
rect 19664 13610 20319 13674
rect 20383 13610 21038 13674
rect 21102 13610 21757 13674
rect 21821 13610 22476 13674
rect 22540 13610 23195 13674
rect 23259 13610 23280 13674
rect 16108 13582 23280 13610
rect 16110 13454 16310 13482
rect 16110 13390 16138 13454
rect 16202 13450 16218 13454
rect 16202 13390 16218 13394
rect 16282 13390 16310 13454
rect 17125 13462 17191 13465
rect 17258 13462 17264 13464
rect 17125 13460 17264 13462
rect 17125 13404 17130 13460
rect 17186 13404 17264 13460
rect 17125 13402 17264 13404
rect 17125 13399 17191 13402
rect 17258 13400 17264 13402
rect 17328 13400 17334 13464
rect 16110 13362 16310 13390
rect 900 13264 2532 13292
rect 900 13200 924 13264
rect 988 13200 1004 13264
rect 1068 13200 1084 13264
rect 1148 13200 1164 13264
rect 1228 13200 1244 13264
rect 1308 13200 1324 13264
rect 1388 13200 1404 13264
rect 1468 13200 1484 13264
rect 1548 13200 1564 13264
rect 1628 13200 1644 13264
rect 1708 13200 1724 13264
rect 1788 13200 1804 13264
rect 1868 13200 1884 13264
rect 1948 13200 1964 13264
rect 2028 13200 2044 13264
rect 2108 13200 2124 13264
rect 2188 13200 2204 13264
rect 2268 13200 2284 13264
rect 2348 13200 2364 13264
rect 2428 13200 2444 13264
rect 2508 13200 2532 13264
rect 900 13172 2532 13200
rect 46104 13264 47736 13292
rect 46104 13200 46128 13264
rect 46192 13200 46208 13264
rect 46272 13200 46288 13264
rect 46352 13200 46368 13264
rect 46432 13200 46448 13264
rect 46512 13200 46528 13264
rect 46592 13200 46608 13264
rect 46672 13200 46688 13264
rect 46752 13200 46768 13264
rect 46832 13200 46848 13264
rect 46912 13200 46928 13264
rect 46992 13200 47008 13264
rect 47072 13200 47088 13264
rect 47152 13200 47168 13264
rect 47232 13200 47248 13264
rect 47312 13200 47328 13264
rect 47392 13200 47408 13264
rect 47472 13200 47488 13264
rect 47552 13200 47568 13264
rect 47632 13200 47648 13264
rect 47712 13200 47736 13264
rect 46104 13172 47736 13200
rect 3348 11384 4980 11412
rect 3348 11320 3372 11384
rect 3436 11320 3452 11384
rect 3516 11320 3532 11384
rect 3596 11320 3612 11384
rect 3676 11320 3692 11384
rect 3756 11320 3772 11384
rect 3836 11320 3852 11384
rect 3916 11320 3932 11384
rect 3996 11320 4012 11384
rect 4076 11320 4092 11384
rect 4156 11320 4172 11384
rect 4236 11320 4252 11384
rect 4316 11320 4332 11384
rect 4396 11320 4412 11384
rect 4476 11320 4492 11384
rect 4556 11320 4572 11384
rect 4636 11320 4652 11384
rect 4716 11320 4732 11384
rect 4796 11320 4812 11384
rect 4876 11320 4892 11384
rect 4956 11320 4980 11384
rect 3348 11292 4980 11320
rect 43656 11384 45288 11412
rect 43656 11320 43680 11384
rect 43744 11320 43760 11384
rect 43824 11320 43840 11384
rect 43904 11320 43920 11384
rect 43984 11320 44000 11384
rect 44064 11320 44080 11384
rect 44144 11320 44160 11384
rect 44224 11320 44240 11384
rect 44304 11320 44320 11384
rect 44384 11320 44400 11384
rect 44464 11320 44480 11384
rect 44544 11320 44560 11384
rect 44624 11320 44640 11384
rect 44704 11320 44720 11384
rect 44784 11320 44800 11384
rect 44864 11320 44880 11384
rect 44944 11320 44960 11384
rect 45024 11320 45040 11384
rect 45104 11320 45120 11384
rect 45184 11320 45200 11384
rect 45264 11320 45288 11384
rect 43656 11292 45288 11320
rect 16108 11110 23280 11122
rect 16108 11054 16140 11110
rect 16196 11054 16220 11110
rect 16276 11094 23280 11110
rect 16276 11054 16724 11094
rect 16108 11030 16724 11054
rect 16788 11030 17443 11094
rect 17507 11030 18162 11094
rect 18226 11030 18881 11094
rect 18945 11030 19600 11094
rect 19664 11030 20319 11094
rect 20383 11030 21038 11094
rect 21102 11030 21757 11094
rect 21821 11030 22476 11094
rect 22540 11030 23195 11094
rect 23259 11030 23280 11094
rect 23468 11082 23474 11146
rect 23538 11144 23544 11146
rect 23657 11144 23723 11147
rect 23538 11142 23723 11144
rect 23538 11086 23662 11142
rect 23718 11086 23723 11142
rect 23538 11084 23723 11086
rect 23538 11082 23544 11084
rect 23657 11081 23723 11084
rect 16108 11014 23280 11030
rect 16108 10950 16724 11014
rect 16788 10950 17443 11014
rect 17507 10950 18162 11014
rect 18226 10950 18881 11014
rect 18945 10950 19600 11014
rect 19664 10950 20319 11014
rect 20383 10950 21038 11014
rect 21102 10950 21757 11014
rect 21821 10950 22476 11014
rect 22540 10950 23195 11014
rect 23259 10950 23280 11014
rect 16108 10934 23280 10950
rect 16108 10870 16724 10934
rect 16788 10870 17443 10934
rect 17507 10870 18162 10934
rect 18226 10870 18881 10934
rect 18945 10870 19600 10934
rect 19664 10870 20319 10934
rect 20383 10870 21038 10934
rect 21102 10870 21757 10934
rect 21821 10870 22476 10934
rect 22540 10870 23195 10934
rect 23259 10870 23280 10934
rect 16108 10854 23280 10870
rect 16108 10790 16724 10854
rect 16788 10790 17443 10854
rect 17507 10790 18162 10854
rect 18226 10790 18881 10854
rect 18945 10790 19600 10854
rect 19664 10790 20319 10854
rect 20383 10790 21038 10854
rect 21102 10790 21757 10854
rect 21821 10790 22476 10854
rect 22540 10790 23195 10854
rect 23259 10790 23280 10854
rect 16108 10774 23280 10790
rect 16108 10710 16724 10774
rect 16788 10710 17443 10774
rect 17507 10710 18162 10774
rect 18226 10710 18881 10774
rect 18945 10710 19600 10774
rect 19664 10710 20319 10774
rect 20383 10710 21038 10774
rect 21102 10710 21757 10774
rect 21821 10710 22476 10774
rect 22540 10710 23195 10774
rect 23259 10710 23280 10774
rect 16108 10694 23280 10710
rect 16108 10630 16724 10694
rect 16788 10630 17443 10694
rect 17507 10630 18162 10694
rect 18226 10630 18881 10694
rect 18945 10630 19600 10694
rect 19664 10630 20319 10694
rect 20383 10630 21038 10694
rect 21102 10630 21757 10694
rect 21821 10630 22476 10694
rect 22540 10630 23195 10694
rect 23259 10630 23280 10694
rect 16108 10614 23280 10630
rect 16108 10550 16724 10614
rect 16788 10550 17443 10614
rect 17507 10550 18162 10614
rect 18226 10550 18881 10614
rect 18945 10550 19600 10614
rect 19664 10550 20319 10614
rect 20383 10550 21038 10614
rect 21102 10550 21757 10614
rect 21821 10550 22476 10614
rect 22540 10550 23195 10614
rect 23259 10550 23280 10614
rect 16108 10394 23280 10550
rect 16108 10330 16724 10394
rect 16788 10330 17443 10394
rect 17507 10330 18162 10394
rect 18226 10330 18881 10394
rect 18945 10330 19600 10394
rect 19664 10330 20319 10394
rect 20383 10330 21038 10394
rect 21102 10330 21757 10394
rect 21821 10330 22476 10394
rect 22540 10330 23195 10394
rect 23259 10330 23280 10394
rect 16108 10314 23280 10330
rect 16108 10250 16724 10314
rect 16788 10250 17443 10314
rect 17507 10250 18162 10314
rect 18226 10250 18881 10314
rect 18945 10250 19600 10314
rect 19664 10250 20319 10314
rect 20383 10250 21038 10314
rect 21102 10250 21757 10314
rect 21821 10250 22476 10314
rect 22540 10250 23195 10314
rect 23259 10250 23280 10314
rect 16108 10234 23280 10250
rect 16108 10170 16724 10234
rect 16788 10170 17443 10234
rect 17507 10170 18162 10234
rect 18226 10170 18881 10234
rect 18945 10170 19600 10234
rect 19664 10170 20319 10234
rect 20383 10170 21038 10234
rect 21102 10170 21757 10234
rect 21821 10170 22476 10234
rect 22540 10170 23195 10234
rect 23259 10170 23280 10234
rect 16108 10154 23280 10170
rect 16108 10090 16724 10154
rect 16788 10090 17443 10154
rect 17507 10090 18162 10154
rect 18226 10090 18881 10154
rect 18945 10090 19600 10154
rect 19664 10090 20319 10154
rect 20383 10090 21038 10154
rect 21102 10090 21757 10154
rect 21821 10090 22476 10154
rect 22540 10090 23195 10154
rect 23259 10090 23280 10154
rect 16108 10074 23280 10090
rect 16108 10010 16724 10074
rect 16788 10010 17443 10074
rect 17507 10010 18162 10074
rect 18226 10010 18881 10074
rect 18945 10010 19600 10074
rect 19664 10010 20319 10074
rect 20383 10010 21038 10074
rect 21102 10010 21757 10074
rect 21821 10010 22476 10074
rect 22540 10010 23195 10074
rect 23259 10010 23280 10074
rect 16108 9994 23280 10010
rect 16108 9930 16724 9994
rect 16788 9930 17443 9994
rect 17507 9930 18162 9994
rect 18226 9930 18881 9994
rect 18945 9930 19600 9994
rect 19664 9930 20319 9994
rect 20383 9930 21038 9994
rect 21102 9930 21757 9994
rect 21821 9930 22476 9994
rect 22540 9930 23195 9994
rect 23259 9930 23280 9994
rect 16108 9914 23280 9930
rect 16108 9850 16724 9914
rect 16788 9850 17443 9914
rect 17507 9850 18162 9914
rect 18226 9850 18881 9914
rect 18945 9850 19600 9914
rect 19664 9850 20319 9914
rect 20383 9850 21038 9914
rect 21102 9850 21757 9914
rect 21821 9850 22476 9914
rect 22540 9850 23195 9914
rect 23259 9850 23280 9914
rect 16108 9822 23280 9850
rect 16110 9694 16310 9722
rect 16110 9630 16138 9694
rect 16202 9690 16218 9694
rect 16202 9630 16218 9634
rect 16282 9630 16310 9694
rect 16110 9602 16310 9630
rect 17125 9680 17191 9683
rect 17258 9680 17264 9682
rect 17125 9678 17264 9680
rect 17125 9622 17130 9678
rect 17186 9622 17264 9678
rect 17125 9620 17264 9622
rect 17125 9617 17191 9620
rect 17258 9618 17264 9620
rect 17328 9618 17334 9682
rect 900 9504 2532 9532
rect 900 9440 924 9504
rect 988 9440 1004 9504
rect 1068 9440 1084 9504
rect 1148 9440 1164 9504
rect 1228 9440 1244 9504
rect 1308 9440 1324 9504
rect 1388 9440 1404 9504
rect 1468 9440 1484 9504
rect 1548 9440 1564 9504
rect 1628 9440 1644 9504
rect 1708 9440 1724 9504
rect 1788 9440 1804 9504
rect 1868 9440 1884 9504
rect 1948 9440 1964 9504
rect 2028 9440 2044 9504
rect 2108 9440 2124 9504
rect 2188 9440 2204 9504
rect 2268 9440 2284 9504
rect 2348 9440 2364 9504
rect 2428 9440 2444 9504
rect 2508 9440 2532 9504
rect 900 9412 2532 9440
rect 46104 9504 47736 9532
rect 46104 9440 46128 9504
rect 46192 9440 46208 9504
rect 46272 9440 46288 9504
rect 46352 9440 46368 9504
rect 46432 9440 46448 9504
rect 46512 9440 46528 9504
rect 46592 9440 46608 9504
rect 46672 9440 46688 9504
rect 46752 9440 46768 9504
rect 46832 9440 46848 9504
rect 46912 9440 46928 9504
rect 46992 9440 47008 9504
rect 47072 9440 47088 9504
rect 47152 9440 47168 9504
rect 47232 9440 47248 9504
rect 47312 9440 47328 9504
rect 47392 9440 47408 9504
rect 47472 9440 47488 9504
rect 47552 9440 47568 9504
rect 47632 9440 47648 9504
rect 47712 9440 47736 9504
rect 46104 9412 47736 9440
rect 3348 7624 4980 7652
rect 3348 7560 3372 7624
rect 3436 7560 3452 7624
rect 3516 7560 3532 7624
rect 3596 7560 3612 7624
rect 3676 7560 3692 7624
rect 3756 7560 3772 7624
rect 3836 7560 3852 7624
rect 3916 7560 3932 7624
rect 3996 7560 4012 7624
rect 4076 7560 4092 7624
rect 4156 7560 4172 7624
rect 4236 7560 4252 7624
rect 4316 7560 4332 7624
rect 4396 7560 4412 7624
rect 4476 7560 4492 7624
rect 4556 7560 4572 7624
rect 4636 7560 4652 7624
rect 4716 7560 4732 7624
rect 4796 7560 4812 7624
rect 4876 7560 4892 7624
rect 4956 7560 4980 7624
rect 3348 7532 4980 7560
rect 43656 7624 45288 7652
rect 43656 7560 43680 7624
rect 43744 7560 43760 7624
rect 43824 7560 43840 7624
rect 43904 7560 43920 7624
rect 43984 7560 44000 7624
rect 44064 7560 44080 7624
rect 44144 7560 44160 7624
rect 44224 7560 44240 7624
rect 44304 7560 44320 7624
rect 44384 7560 44400 7624
rect 44464 7560 44480 7624
rect 44544 7560 44560 7624
rect 44624 7560 44640 7624
rect 44704 7560 44720 7624
rect 44784 7560 44800 7624
rect 44864 7560 44880 7624
rect 44944 7560 44960 7624
rect 45024 7560 45040 7624
rect 45104 7560 45120 7624
rect 45184 7560 45200 7624
rect 45264 7560 45288 7624
rect 43656 7532 45288 7560
rect 19517 6508 19583 6511
rect 25681 6508 25747 6511
rect 19517 6506 25747 6508
rect 19517 6450 19522 6506
rect 19578 6450 25686 6506
rect 25742 6450 25747 6506
rect 19517 6448 25747 6450
rect 19517 6445 19583 6448
rect 25681 6445 25747 6448
rect 17769 6142 17835 6145
rect 28349 6142 28415 6145
rect 17769 6140 28415 6142
rect 17769 6084 17774 6140
rect 17830 6084 28354 6140
rect 28410 6084 28415 6140
rect 17769 6082 28415 6084
rect 17769 6079 17835 6082
rect 28349 6079 28415 6082
rect 900 5744 2532 5772
rect 900 5680 924 5744
rect 988 5680 1004 5744
rect 1068 5680 1084 5744
rect 1148 5680 1164 5744
rect 1228 5680 1244 5744
rect 1308 5680 1324 5744
rect 1388 5680 1404 5744
rect 1468 5680 1484 5744
rect 1548 5680 1564 5744
rect 1628 5680 1644 5744
rect 1708 5680 1724 5744
rect 1788 5680 1804 5744
rect 1868 5680 1884 5744
rect 1948 5680 1964 5744
rect 2028 5680 2044 5744
rect 2108 5680 2124 5744
rect 2188 5680 2204 5744
rect 2268 5680 2284 5744
rect 2348 5680 2364 5744
rect 2428 5680 2444 5744
rect 2508 5680 2532 5744
rect 900 5652 2532 5680
rect 46104 5744 47736 5772
rect 46104 5680 46128 5744
rect 46192 5680 46208 5744
rect 46272 5680 46288 5744
rect 46352 5680 46368 5744
rect 46432 5680 46448 5744
rect 46512 5680 46528 5744
rect 46592 5680 46608 5744
rect 46672 5680 46688 5744
rect 46752 5680 46768 5744
rect 46832 5680 46848 5744
rect 46912 5680 46928 5744
rect 46992 5680 47008 5744
rect 47072 5680 47088 5744
rect 47152 5680 47168 5744
rect 47232 5680 47248 5744
rect 47312 5680 47328 5744
rect 47392 5680 47408 5744
rect 47472 5680 47488 5744
rect 47552 5680 47568 5744
rect 47632 5680 47648 5744
rect 47712 5680 47736 5744
rect 46104 5652 47736 5680
<< via3 >>
rect 3372 41460 3436 41464
rect 3372 41404 3376 41460
rect 3376 41404 3432 41460
rect 3432 41404 3436 41460
rect 3372 41400 3436 41404
rect 3452 41460 3516 41464
rect 3452 41404 3456 41460
rect 3456 41404 3512 41460
rect 3512 41404 3516 41460
rect 3452 41400 3516 41404
rect 3532 41460 3596 41464
rect 3532 41404 3536 41460
rect 3536 41404 3592 41460
rect 3592 41404 3596 41460
rect 3532 41400 3596 41404
rect 3612 41460 3676 41464
rect 3612 41404 3616 41460
rect 3616 41404 3672 41460
rect 3672 41404 3676 41460
rect 3612 41400 3676 41404
rect 3692 41460 3756 41464
rect 3692 41404 3696 41460
rect 3696 41404 3752 41460
rect 3752 41404 3756 41460
rect 3692 41400 3756 41404
rect 3772 41460 3836 41464
rect 3772 41404 3776 41460
rect 3776 41404 3832 41460
rect 3832 41404 3836 41460
rect 3772 41400 3836 41404
rect 3852 41460 3916 41464
rect 3852 41404 3856 41460
rect 3856 41404 3912 41460
rect 3912 41404 3916 41460
rect 3852 41400 3916 41404
rect 3932 41460 3996 41464
rect 3932 41404 3936 41460
rect 3936 41404 3992 41460
rect 3992 41404 3996 41460
rect 3932 41400 3996 41404
rect 4012 41460 4076 41464
rect 4012 41404 4016 41460
rect 4016 41404 4072 41460
rect 4072 41404 4076 41460
rect 4012 41400 4076 41404
rect 4092 41460 4156 41464
rect 4092 41404 4096 41460
rect 4096 41404 4152 41460
rect 4152 41404 4156 41460
rect 4092 41400 4156 41404
rect 4172 41460 4236 41464
rect 4172 41404 4176 41460
rect 4176 41404 4232 41460
rect 4232 41404 4236 41460
rect 4172 41400 4236 41404
rect 4252 41460 4316 41464
rect 4252 41404 4256 41460
rect 4256 41404 4312 41460
rect 4312 41404 4316 41460
rect 4252 41400 4316 41404
rect 4332 41460 4396 41464
rect 4332 41404 4336 41460
rect 4336 41404 4392 41460
rect 4392 41404 4396 41460
rect 4332 41400 4396 41404
rect 4412 41460 4476 41464
rect 4412 41404 4416 41460
rect 4416 41404 4472 41460
rect 4472 41404 4476 41460
rect 4412 41400 4476 41404
rect 4492 41460 4556 41464
rect 4492 41404 4496 41460
rect 4496 41404 4552 41460
rect 4552 41404 4556 41460
rect 4492 41400 4556 41404
rect 4572 41460 4636 41464
rect 4572 41404 4576 41460
rect 4576 41404 4632 41460
rect 4632 41404 4636 41460
rect 4572 41400 4636 41404
rect 4652 41460 4716 41464
rect 4652 41404 4656 41460
rect 4656 41404 4712 41460
rect 4712 41404 4716 41460
rect 4652 41400 4716 41404
rect 4732 41460 4796 41464
rect 4732 41404 4736 41460
rect 4736 41404 4792 41460
rect 4792 41404 4796 41460
rect 4732 41400 4796 41404
rect 4812 41460 4876 41464
rect 4812 41404 4816 41460
rect 4816 41404 4872 41460
rect 4872 41404 4876 41460
rect 4812 41400 4876 41404
rect 4892 41460 4956 41464
rect 4892 41404 4896 41460
rect 4896 41404 4952 41460
rect 4952 41404 4956 41460
rect 4892 41400 4956 41404
rect 12434 41398 12498 41402
rect 12434 41342 12438 41398
rect 12438 41342 12494 41398
rect 12494 41342 12498 41398
rect 12434 41338 12498 41342
rect 43680 41460 43744 41464
rect 43680 41404 43684 41460
rect 43684 41404 43740 41460
rect 43740 41404 43744 41460
rect 43680 41400 43744 41404
rect 43760 41460 43824 41464
rect 43760 41404 43764 41460
rect 43764 41404 43820 41460
rect 43820 41404 43824 41460
rect 43760 41400 43824 41404
rect 43840 41460 43904 41464
rect 43840 41404 43844 41460
rect 43844 41404 43900 41460
rect 43900 41404 43904 41460
rect 43840 41400 43904 41404
rect 43920 41460 43984 41464
rect 43920 41404 43924 41460
rect 43924 41404 43980 41460
rect 43980 41404 43984 41460
rect 43920 41400 43984 41404
rect 44000 41460 44064 41464
rect 44000 41404 44004 41460
rect 44004 41404 44060 41460
rect 44060 41404 44064 41460
rect 44000 41400 44064 41404
rect 44080 41460 44144 41464
rect 44080 41404 44084 41460
rect 44084 41404 44140 41460
rect 44140 41404 44144 41460
rect 44080 41400 44144 41404
rect 44160 41460 44224 41464
rect 44160 41404 44164 41460
rect 44164 41404 44220 41460
rect 44220 41404 44224 41460
rect 44160 41400 44224 41404
rect 44240 41460 44304 41464
rect 44240 41404 44244 41460
rect 44244 41404 44300 41460
rect 44300 41404 44304 41460
rect 44240 41400 44304 41404
rect 44320 41460 44384 41464
rect 44320 41404 44324 41460
rect 44324 41404 44380 41460
rect 44380 41404 44384 41460
rect 44320 41400 44384 41404
rect 44400 41460 44464 41464
rect 44400 41404 44404 41460
rect 44404 41404 44460 41460
rect 44460 41404 44464 41460
rect 44400 41400 44464 41404
rect 44480 41460 44544 41464
rect 44480 41404 44484 41460
rect 44484 41404 44540 41460
rect 44540 41404 44544 41460
rect 44480 41400 44544 41404
rect 44560 41460 44624 41464
rect 44560 41404 44564 41460
rect 44564 41404 44620 41460
rect 44620 41404 44624 41460
rect 44560 41400 44624 41404
rect 44640 41460 44704 41464
rect 44640 41404 44644 41460
rect 44644 41404 44700 41460
rect 44700 41404 44704 41460
rect 44640 41400 44704 41404
rect 44720 41460 44784 41464
rect 44720 41404 44724 41460
rect 44724 41404 44780 41460
rect 44780 41404 44784 41460
rect 44720 41400 44784 41404
rect 44800 41460 44864 41464
rect 44800 41404 44804 41460
rect 44804 41404 44860 41460
rect 44860 41404 44864 41460
rect 44800 41400 44864 41404
rect 44880 41460 44944 41464
rect 44880 41404 44884 41460
rect 44884 41404 44940 41460
rect 44940 41404 44944 41460
rect 44880 41400 44944 41404
rect 44960 41460 45024 41464
rect 44960 41404 44964 41460
rect 44964 41404 45020 41460
rect 45020 41404 45024 41460
rect 44960 41400 45024 41404
rect 45040 41460 45104 41464
rect 45040 41404 45044 41460
rect 45044 41404 45100 41460
rect 45100 41404 45104 41460
rect 45040 41400 45104 41404
rect 45120 41460 45184 41464
rect 45120 41404 45124 41460
rect 45124 41404 45180 41460
rect 45180 41404 45184 41460
rect 45120 41400 45184 41404
rect 45200 41460 45264 41464
rect 45200 41404 45204 41460
rect 45204 41404 45260 41460
rect 45260 41404 45264 41460
rect 45200 41400 45264 41404
rect 7414 41110 7478 41174
rect 8133 41110 8197 41174
rect 8852 41110 8916 41174
rect 9571 41110 9635 41174
rect 10290 41110 10354 41174
rect 11009 41110 11073 41174
rect 11728 41110 11792 41174
rect 12447 41110 12511 41174
rect 13166 41110 13230 41174
rect 13885 41110 13949 41174
rect 7414 41030 7478 41094
rect 8133 41030 8197 41094
rect 8852 41030 8916 41094
rect 9571 41030 9635 41094
rect 10290 41030 10354 41094
rect 11009 41030 11073 41094
rect 11728 41030 11792 41094
rect 12447 41030 12511 41094
rect 13166 41030 13230 41094
rect 13885 41030 13949 41094
rect 7414 40950 7478 41014
rect 8133 40950 8197 41014
rect 8852 40950 8916 41014
rect 9571 40950 9635 41014
rect 10290 40950 10354 41014
rect 11009 40950 11073 41014
rect 11728 40950 11792 41014
rect 12447 40950 12511 41014
rect 13166 40950 13230 41014
rect 13885 40950 13949 41014
rect 7414 40870 7478 40934
rect 8133 40870 8197 40934
rect 8852 40870 8916 40934
rect 9571 40870 9635 40934
rect 10290 40870 10354 40934
rect 11009 40870 11073 40934
rect 11728 40870 11792 40934
rect 12447 40870 12511 40934
rect 13166 40870 13230 40934
rect 13885 40870 13949 40934
rect 7414 40790 7478 40854
rect 8133 40790 8197 40854
rect 8852 40790 8916 40854
rect 9571 40790 9635 40854
rect 10290 40790 10354 40854
rect 11009 40790 11073 40854
rect 11728 40790 11792 40854
rect 12447 40790 12511 40854
rect 13166 40790 13230 40854
rect 13885 40790 13949 40854
rect 7414 40710 7478 40774
rect 8133 40710 8197 40774
rect 8852 40710 8916 40774
rect 9571 40710 9635 40774
rect 10290 40710 10354 40774
rect 11009 40710 11073 40774
rect 11728 40710 11792 40774
rect 12447 40710 12511 40774
rect 13166 40710 13230 40774
rect 13885 40710 13949 40774
rect 7414 40630 7478 40694
rect 8133 40630 8197 40694
rect 8852 40630 8916 40694
rect 9571 40630 9635 40694
rect 10290 40630 10354 40694
rect 11009 40630 11073 40694
rect 11728 40630 11792 40694
rect 12447 40630 12511 40694
rect 13166 40630 13230 40694
rect 13885 40630 13949 40694
rect 7414 40410 7478 40474
rect 8133 40410 8197 40474
rect 8852 40410 8916 40474
rect 9571 40410 9635 40474
rect 10290 40410 10354 40474
rect 11009 40410 11073 40474
rect 11728 40410 11792 40474
rect 12447 40410 12511 40474
rect 13166 40410 13230 40474
rect 13885 40410 13949 40474
rect 7414 40330 7478 40394
rect 8133 40330 8197 40394
rect 8852 40330 8916 40394
rect 9571 40330 9635 40394
rect 10290 40330 10354 40394
rect 11009 40330 11073 40394
rect 11728 40330 11792 40394
rect 12447 40330 12511 40394
rect 13166 40330 13230 40394
rect 13885 40330 13949 40394
rect 7414 40250 7478 40314
rect 8133 40250 8197 40314
rect 8852 40250 8916 40314
rect 9571 40250 9635 40314
rect 10290 40250 10354 40314
rect 11009 40250 11073 40314
rect 11728 40250 11792 40314
rect 12447 40250 12511 40314
rect 13166 40250 13230 40314
rect 13885 40250 13949 40314
rect 7414 40170 7478 40234
rect 8133 40170 8197 40234
rect 8852 40170 8916 40234
rect 9571 40170 9635 40234
rect 10290 40170 10354 40234
rect 11009 40170 11073 40234
rect 11728 40170 11792 40234
rect 12447 40170 12511 40234
rect 13166 40170 13230 40234
rect 13885 40170 13949 40234
rect 7414 40090 7478 40154
rect 8133 40090 8197 40154
rect 8852 40090 8916 40154
rect 9571 40090 9635 40154
rect 10290 40090 10354 40154
rect 11009 40090 11073 40154
rect 11728 40090 11792 40154
rect 12447 40090 12511 40154
rect 13166 40090 13230 40154
rect 13885 40090 13949 40154
rect 7414 40010 7478 40074
rect 8133 40010 8197 40074
rect 8852 40010 8916 40074
rect 9571 40010 9635 40074
rect 10290 40010 10354 40074
rect 11009 40010 11073 40074
rect 11728 40010 11792 40074
rect 12447 40010 12511 40074
rect 13166 40010 13230 40074
rect 13885 40010 13949 40074
rect 7414 39930 7478 39994
rect 8133 39930 8197 39994
rect 8852 39930 8916 39994
rect 9571 39930 9635 39994
rect 10290 39930 10354 39994
rect 11009 39930 11073 39994
rect 11728 39930 11792 39994
rect 12447 39930 12511 39994
rect 13166 39930 13230 39994
rect 13885 39930 13949 39994
rect 6828 39770 6892 39774
rect 6908 39770 6972 39774
rect 6828 39714 6872 39770
rect 6872 39714 6892 39770
rect 6908 39714 6928 39770
rect 6928 39714 6972 39770
rect 6828 39710 6892 39714
rect 6908 39710 6972 39714
rect 13676 39630 13740 39694
rect 27614 39690 27678 39694
rect 27614 39634 27618 39690
rect 27618 39634 27674 39690
rect 27674 39634 27678 39690
rect 27614 39630 27678 39634
rect 924 39580 988 39584
rect 924 39524 928 39580
rect 928 39524 984 39580
rect 984 39524 988 39580
rect 924 39520 988 39524
rect 1004 39580 1068 39584
rect 1004 39524 1008 39580
rect 1008 39524 1064 39580
rect 1064 39524 1068 39580
rect 1004 39520 1068 39524
rect 1084 39580 1148 39584
rect 1084 39524 1088 39580
rect 1088 39524 1144 39580
rect 1144 39524 1148 39580
rect 1084 39520 1148 39524
rect 1164 39580 1228 39584
rect 1164 39524 1168 39580
rect 1168 39524 1224 39580
rect 1224 39524 1228 39580
rect 1164 39520 1228 39524
rect 1244 39580 1308 39584
rect 1244 39524 1248 39580
rect 1248 39524 1304 39580
rect 1304 39524 1308 39580
rect 1244 39520 1308 39524
rect 1324 39580 1388 39584
rect 1324 39524 1328 39580
rect 1328 39524 1384 39580
rect 1384 39524 1388 39580
rect 1324 39520 1388 39524
rect 1404 39580 1468 39584
rect 1404 39524 1408 39580
rect 1408 39524 1464 39580
rect 1464 39524 1468 39580
rect 1404 39520 1468 39524
rect 1484 39580 1548 39584
rect 1484 39524 1488 39580
rect 1488 39524 1544 39580
rect 1544 39524 1548 39580
rect 1484 39520 1548 39524
rect 1564 39580 1628 39584
rect 1564 39524 1568 39580
rect 1568 39524 1624 39580
rect 1624 39524 1628 39580
rect 1564 39520 1628 39524
rect 1644 39580 1708 39584
rect 1644 39524 1648 39580
rect 1648 39524 1704 39580
rect 1704 39524 1708 39580
rect 1644 39520 1708 39524
rect 1724 39580 1788 39584
rect 1724 39524 1728 39580
rect 1728 39524 1784 39580
rect 1784 39524 1788 39580
rect 1724 39520 1788 39524
rect 1804 39580 1868 39584
rect 1804 39524 1808 39580
rect 1808 39524 1864 39580
rect 1864 39524 1868 39580
rect 1804 39520 1868 39524
rect 1884 39580 1948 39584
rect 1884 39524 1888 39580
rect 1888 39524 1944 39580
rect 1944 39524 1948 39580
rect 1884 39520 1948 39524
rect 1964 39580 2028 39584
rect 1964 39524 1968 39580
rect 1968 39524 2024 39580
rect 2024 39524 2028 39580
rect 1964 39520 2028 39524
rect 2044 39580 2108 39584
rect 2044 39524 2048 39580
rect 2048 39524 2104 39580
rect 2104 39524 2108 39580
rect 2044 39520 2108 39524
rect 2124 39580 2188 39584
rect 2124 39524 2128 39580
rect 2128 39524 2184 39580
rect 2184 39524 2188 39580
rect 2124 39520 2188 39524
rect 2204 39580 2268 39584
rect 2204 39524 2208 39580
rect 2208 39524 2264 39580
rect 2264 39524 2268 39580
rect 2204 39520 2268 39524
rect 2284 39580 2348 39584
rect 2284 39524 2288 39580
rect 2288 39524 2344 39580
rect 2344 39524 2348 39580
rect 2284 39520 2348 39524
rect 2364 39580 2428 39584
rect 2364 39524 2368 39580
rect 2368 39524 2424 39580
rect 2424 39524 2428 39580
rect 2364 39520 2428 39524
rect 2444 39580 2508 39584
rect 2444 39524 2448 39580
rect 2448 39524 2504 39580
rect 2504 39524 2508 39580
rect 2444 39520 2508 39524
rect 46128 39580 46192 39584
rect 46128 39524 46132 39580
rect 46132 39524 46188 39580
rect 46188 39524 46192 39580
rect 46128 39520 46192 39524
rect 46208 39580 46272 39584
rect 46208 39524 46212 39580
rect 46212 39524 46268 39580
rect 46268 39524 46272 39580
rect 46208 39520 46272 39524
rect 46288 39580 46352 39584
rect 46288 39524 46292 39580
rect 46292 39524 46348 39580
rect 46348 39524 46352 39580
rect 46288 39520 46352 39524
rect 46368 39580 46432 39584
rect 46368 39524 46372 39580
rect 46372 39524 46428 39580
rect 46428 39524 46432 39580
rect 46368 39520 46432 39524
rect 46448 39580 46512 39584
rect 46448 39524 46452 39580
rect 46452 39524 46508 39580
rect 46508 39524 46512 39580
rect 46448 39520 46512 39524
rect 46528 39580 46592 39584
rect 46528 39524 46532 39580
rect 46532 39524 46588 39580
rect 46588 39524 46592 39580
rect 46528 39520 46592 39524
rect 46608 39580 46672 39584
rect 46608 39524 46612 39580
rect 46612 39524 46668 39580
rect 46668 39524 46672 39580
rect 46608 39520 46672 39524
rect 46688 39580 46752 39584
rect 46688 39524 46692 39580
rect 46692 39524 46748 39580
rect 46748 39524 46752 39580
rect 46688 39520 46752 39524
rect 46768 39580 46832 39584
rect 46768 39524 46772 39580
rect 46772 39524 46828 39580
rect 46828 39524 46832 39580
rect 46768 39520 46832 39524
rect 46848 39580 46912 39584
rect 46848 39524 46852 39580
rect 46852 39524 46908 39580
rect 46908 39524 46912 39580
rect 46848 39520 46912 39524
rect 46928 39580 46992 39584
rect 46928 39524 46932 39580
rect 46932 39524 46988 39580
rect 46988 39524 46992 39580
rect 46928 39520 46992 39524
rect 47008 39580 47072 39584
rect 47008 39524 47012 39580
rect 47012 39524 47068 39580
rect 47068 39524 47072 39580
rect 47008 39520 47072 39524
rect 47088 39580 47152 39584
rect 47088 39524 47092 39580
rect 47092 39524 47148 39580
rect 47148 39524 47152 39580
rect 47088 39520 47152 39524
rect 47168 39580 47232 39584
rect 47168 39524 47172 39580
rect 47172 39524 47228 39580
rect 47228 39524 47232 39580
rect 47168 39520 47232 39524
rect 47248 39580 47312 39584
rect 47248 39524 47252 39580
rect 47252 39524 47308 39580
rect 47308 39524 47312 39580
rect 47248 39520 47312 39524
rect 47328 39580 47392 39584
rect 47328 39524 47332 39580
rect 47332 39524 47388 39580
rect 47388 39524 47392 39580
rect 47328 39520 47392 39524
rect 47408 39580 47472 39584
rect 47408 39524 47412 39580
rect 47412 39524 47468 39580
rect 47468 39524 47472 39580
rect 47408 39520 47472 39524
rect 47488 39580 47552 39584
rect 47488 39524 47492 39580
rect 47492 39524 47548 39580
rect 47548 39524 47552 39580
rect 47488 39520 47552 39524
rect 47568 39580 47632 39584
rect 47568 39524 47572 39580
rect 47572 39524 47628 39580
rect 47628 39524 47632 39580
rect 47568 39520 47632 39524
rect 47648 39580 47712 39584
rect 47648 39524 47652 39580
rect 47652 39524 47708 39580
rect 47708 39524 47712 39580
rect 47648 39520 47712 39524
rect 3372 37700 3436 37704
rect 3372 37644 3376 37700
rect 3376 37644 3432 37700
rect 3432 37644 3436 37700
rect 3372 37640 3436 37644
rect 3452 37700 3516 37704
rect 3452 37644 3456 37700
rect 3456 37644 3512 37700
rect 3512 37644 3516 37700
rect 3452 37640 3516 37644
rect 3532 37700 3596 37704
rect 3532 37644 3536 37700
rect 3536 37644 3592 37700
rect 3592 37644 3596 37700
rect 3532 37640 3596 37644
rect 3612 37700 3676 37704
rect 3612 37644 3616 37700
rect 3616 37644 3672 37700
rect 3672 37644 3676 37700
rect 3612 37640 3676 37644
rect 3692 37700 3756 37704
rect 3692 37644 3696 37700
rect 3696 37644 3752 37700
rect 3752 37644 3756 37700
rect 3692 37640 3756 37644
rect 3772 37700 3836 37704
rect 3772 37644 3776 37700
rect 3776 37644 3832 37700
rect 3832 37644 3836 37700
rect 3772 37640 3836 37644
rect 3852 37700 3916 37704
rect 3852 37644 3856 37700
rect 3856 37644 3912 37700
rect 3912 37644 3916 37700
rect 3852 37640 3916 37644
rect 3932 37700 3996 37704
rect 3932 37644 3936 37700
rect 3936 37644 3992 37700
rect 3992 37644 3996 37700
rect 3932 37640 3996 37644
rect 4012 37700 4076 37704
rect 4012 37644 4016 37700
rect 4016 37644 4072 37700
rect 4072 37644 4076 37700
rect 4012 37640 4076 37644
rect 4092 37700 4156 37704
rect 4092 37644 4096 37700
rect 4096 37644 4152 37700
rect 4152 37644 4156 37700
rect 4092 37640 4156 37644
rect 4172 37700 4236 37704
rect 4172 37644 4176 37700
rect 4176 37644 4232 37700
rect 4232 37644 4236 37700
rect 4172 37640 4236 37644
rect 4252 37700 4316 37704
rect 4252 37644 4256 37700
rect 4256 37644 4312 37700
rect 4312 37644 4316 37700
rect 4252 37640 4316 37644
rect 4332 37700 4396 37704
rect 4332 37644 4336 37700
rect 4336 37644 4392 37700
rect 4392 37644 4396 37700
rect 4332 37640 4396 37644
rect 4412 37700 4476 37704
rect 4412 37644 4416 37700
rect 4416 37644 4472 37700
rect 4472 37644 4476 37700
rect 4412 37640 4476 37644
rect 4492 37700 4556 37704
rect 4492 37644 4496 37700
rect 4496 37644 4552 37700
rect 4552 37644 4556 37700
rect 4492 37640 4556 37644
rect 4572 37700 4636 37704
rect 4572 37644 4576 37700
rect 4576 37644 4632 37700
rect 4632 37644 4636 37700
rect 4572 37640 4636 37644
rect 4652 37700 4716 37704
rect 4652 37644 4656 37700
rect 4656 37644 4712 37700
rect 4712 37644 4716 37700
rect 4652 37640 4716 37644
rect 4732 37700 4796 37704
rect 4732 37644 4736 37700
rect 4736 37644 4792 37700
rect 4792 37644 4796 37700
rect 4732 37640 4796 37644
rect 4812 37700 4876 37704
rect 4812 37644 4816 37700
rect 4816 37644 4872 37700
rect 4872 37644 4876 37700
rect 4812 37640 4876 37644
rect 4892 37700 4956 37704
rect 4892 37644 4896 37700
rect 4896 37644 4952 37700
rect 4952 37644 4956 37700
rect 4892 37640 4956 37644
rect 43680 37700 43744 37704
rect 43680 37644 43684 37700
rect 43684 37644 43740 37700
rect 43740 37644 43744 37700
rect 43680 37640 43744 37644
rect 43760 37700 43824 37704
rect 43760 37644 43764 37700
rect 43764 37644 43820 37700
rect 43820 37644 43824 37700
rect 43760 37640 43824 37644
rect 43840 37700 43904 37704
rect 43840 37644 43844 37700
rect 43844 37644 43900 37700
rect 43900 37644 43904 37700
rect 43840 37640 43904 37644
rect 43920 37700 43984 37704
rect 43920 37644 43924 37700
rect 43924 37644 43980 37700
rect 43980 37644 43984 37700
rect 43920 37640 43984 37644
rect 44000 37700 44064 37704
rect 44000 37644 44004 37700
rect 44004 37644 44060 37700
rect 44060 37644 44064 37700
rect 44000 37640 44064 37644
rect 44080 37700 44144 37704
rect 44080 37644 44084 37700
rect 44084 37644 44140 37700
rect 44140 37644 44144 37700
rect 44080 37640 44144 37644
rect 44160 37700 44224 37704
rect 44160 37644 44164 37700
rect 44164 37644 44220 37700
rect 44220 37644 44224 37700
rect 44160 37640 44224 37644
rect 44240 37700 44304 37704
rect 44240 37644 44244 37700
rect 44244 37644 44300 37700
rect 44300 37644 44304 37700
rect 44240 37640 44304 37644
rect 44320 37700 44384 37704
rect 44320 37644 44324 37700
rect 44324 37644 44380 37700
rect 44380 37644 44384 37700
rect 44320 37640 44384 37644
rect 44400 37700 44464 37704
rect 44400 37644 44404 37700
rect 44404 37644 44460 37700
rect 44460 37644 44464 37700
rect 44400 37640 44464 37644
rect 44480 37700 44544 37704
rect 44480 37644 44484 37700
rect 44484 37644 44540 37700
rect 44540 37644 44544 37700
rect 44480 37640 44544 37644
rect 44560 37700 44624 37704
rect 44560 37644 44564 37700
rect 44564 37644 44620 37700
rect 44620 37644 44624 37700
rect 44560 37640 44624 37644
rect 44640 37700 44704 37704
rect 44640 37644 44644 37700
rect 44644 37644 44700 37700
rect 44700 37644 44704 37700
rect 44640 37640 44704 37644
rect 44720 37700 44784 37704
rect 44720 37644 44724 37700
rect 44724 37644 44780 37700
rect 44780 37644 44784 37700
rect 44720 37640 44784 37644
rect 44800 37700 44864 37704
rect 44800 37644 44804 37700
rect 44804 37644 44860 37700
rect 44860 37644 44864 37700
rect 44800 37640 44864 37644
rect 44880 37700 44944 37704
rect 44880 37644 44884 37700
rect 44884 37644 44940 37700
rect 44940 37644 44944 37700
rect 44880 37640 44944 37644
rect 44960 37700 45024 37704
rect 44960 37644 44964 37700
rect 44964 37644 45020 37700
rect 45020 37644 45024 37700
rect 44960 37640 45024 37644
rect 45040 37700 45104 37704
rect 45040 37644 45044 37700
rect 45044 37644 45100 37700
rect 45100 37644 45104 37700
rect 45040 37640 45104 37644
rect 45120 37700 45184 37704
rect 45120 37644 45124 37700
rect 45124 37644 45180 37700
rect 45180 37644 45184 37700
rect 45120 37640 45184 37644
rect 45200 37700 45264 37704
rect 45200 37644 45204 37700
rect 45204 37644 45260 37700
rect 45260 37644 45264 37700
rect 45200 37640 45264 37644
rect 12986 37616 13050 37620
rect 12986 37560 12990 37616
rect 12990 37560 13046 37616
rect 13046 37560 13050 37616
rect 12986 37556 13050 37560
rect 16850 37616 16914 37620
rect 16850 37560 16854 37616
rect 16854 37560 16910 37616
rect 16910 37560 16914 37616
rect 16850 37556 16914 37560
rect 27890 37616 27954 37620
rect 27890 37560 27894 37616
rect 27894 37560 27950 37616
rect 27950 37560 27954 37616
rect 27890 37556 27954 37560
rect 6532 37350 6596 37414
rect 7251 37350 7315 37414
rect 7970 37350 8034 37414
rect 8689 37350 8753 37414
rect 9408 37350 9472 37414
rect 10127 37350 10191 37414
rect 10846 37350 10910 37414
rect 11565 37350 11629 37414
rect 12284 37350 12348 37414
rect 13003 37350 13067 37414
rect 6532 37270 6596 37334
rect 7251 37270 7315 37334
rect 7970 37270 8034 37334
rect 8689 37270 8753 37334
rect 9408 37270 9472 37334
rect 10127 37270 10191 37334
rect 10846 37270 10910 37334
rect 11565 37270 11629 37334
rect 12284 37270 12348 37334
rect 13003 37270 13067 37334
rect 6532 37190 6596 37254
rect 7251 37190 7315 37254
rect 7970 37190 8034 37254
rect 8689 37190 8753 37254
rect 9408 37190 9472 37254
rect 10127 37190 10191 37254
rect 10846 37190 10910 37254
rect 11565 37190 11629 37254
rect 12284 37190 12348 37254
rect 13003 37190 13067 37254
rect 6532 37110 6596 37174
rect 7251 37110 7315 37174
rect 7970 37110 8034 37174
rect 8689 37110 8753 37174
rect 9408 37110 9472 37174
rect 10127 37110 10191 37174
rect 10846 37110 10910 37174
rect 11565 37110 11629 37174
rect 12284 37110 12348 37174
rect 13003 37110 13067 37174
rect 6532 37030 6596 37094
rect 7251 37030 7315 37094
rect 7970 37030 8034 37094
rect 8689 37030 8753 37094
rect 9408 37030 9472 37094
rect 10127 37030 10191 37094
rect 10846 37030 10910 37094
rect 11565 37030 11629 37094
rect 12284 37030 12348 37094
rect 13003 37030 13067 37094
rect 6532 36950 6596 37014
rect 7251 36950 7315 37014
rect 7970 36950 8034 37014
rect 8689 36950 8753 37014
rect 9408 36950 9472 37014
rect 10127 36950 10191 37014
rect 10846 36950 10910 37014
rect 11565 36950 11629 37014
rect 12284 36950 12348 37014
rect 13003 36950 13067 37014
rect 6532 36870 6596 36934
rect 7251 36870 7315 36934
rect 7970 36870 8034 36934
rect 8689 36870 8753 36934
rect 9408 36870 9472 36934
rect 10127 36870 10191 36934
rect 10846 36870 10910 36934
rect 11565 36870 11629 36934
rect 12284 36870 12348 36934
rect 13003 36870 13067 36934
rect 6532 36650 6596 36714
rect 7251 36650 7315 36714
rect 7970 36650 8034 36714
rect 8689 36650 8753 36714
rect 9408 36650 9472 36714
rect 10127 36650 10191 36714
rect 10846 36650 10910 36714
rect 11565 36650 11629 36714
rect 12284 36650 12348 36714
rect 13003 36650 13067 36714
rect 6532 36570 6596 36634
rect 7251 36570 7315 36634
rect 7970 36570 8034 36634
rect 8689 36570 8753 36634
rect 9408 36570 9472 36634
rect 10127 36570 10191 36634
rect 10846 36570 10910 36634
rect 11565 36570 11629 36634
rect 12284 36570 12348 36634
rect 13003 36570 13067 36634
rect 6532 36490 6596 36554
rect 7251 36490 7315 36554
rect 7970 36490 8034 36554
rect 8689 36490 8753 36554
rect 9408 36490 9472 36554
rect 10127 36490 10191 36554
rect 10846 36490 10910 36554
rect 11565 36490 11629 36554
rect 12284 36490 12348 36554
rect 13003 36490 13067 36554
rect 6532 36410 6596 36474
rect 7251 36410 7315 36474
rect 7970 36410 8034 36474
rect 8689 36410 8753 36474
rect 9408 36410 9472 36474
rect 10127 36410 10191 36474
rect 10846 36410 10910 36474
rect 11565 36410 11629 36474
rect 12284 36410 12348 36474
rect 13003 36410 13067 36474
rect 6532 36330 6596 36394
rect 7251 36330 7315 36394
rect 7970 36330 8034 36394
rect 8689 36330 8753 36394
rect 9408 36330 9472 36394
rect 10127 36330 10191 36394
rect 10846 36330 10910 36394
rect 11565 36330 11629 36394
rect 12284 36330 12348 36394
rect 13003 36330 13067 36394
rect 6532 36250 6596 36314
rect 7251 36250 7315 36314
rect 7970 36250 8034 36314
rect 8689 36250 8753 36314
rect 9408 36250 9472 36314
rect 10127 36250 10191 36314
rect 10846 36250 10910 36314
rect 11565 36250 11629 36314
rect 12284 36250 12348 36314
rect 13003 36250 13067 36314
rect 6532 36170 6596 36234
rect 7251 36170 7315 36234
rect 7970 36170 8034 36234
rect 8689 36170 8753 36234
rect 9408 36170 9472 36234
rect 10127 36170 10191 36234
rect 10846 36170 10910 36234
rect 11565 36170 11629 36234
rect 12284 36170 12348 36234
rect 13003 36170 13067 36234
rect 13980 37350 14044 37414
rect 14699 37350 14763 37414
rect 15418 37350 15482 37414
rect 16137 37350 16201 37414
rect 16856 37350 16920 37414
rect 17575 37350 17639 37414
rect 18294 37350 18358 37414
rect 19013 37350 19077 37414
rect 19732 37350 19796 37414
rect 20451 37350 20515 37414
rect 13980 37270 14044 37334
rect 14699 37270 14763 37334
rect 15418 37270 15482 37334
rect 16137 37270 16201 37334
rect 16856 37270 16920 37334
rect 17575 37270 17639 37334
rect 18294 37270 18358 37334
rect 19013 37270 19077 37334
rect 19732 37270 19796 37334
rect 20451 37270 20515 37334
rect 13980 37190 14044 37254
rect 14699 37190 14763 37254
rect 15418 37190 15482 37254
rect 16137 37190 16201 37254
rect 16856 37190 16920 37254
rect 17575 37190 17639 37254
rect 18294 37190 18358 37254
rect 19013 37190 19077 37254
rect 19732 37190 19796 37254
rect 20451 37190 20515 37254
rect 13980 37110 14044 37174
rect 14699 37110 14763 37174
rect 15418 37110 15482 37174
rect 16137 37110 16201 37174
rect 16856 37110 16920 37174
rect 17575 37110 17639 37174
rect 18294 37110 18358 37174
rect 19013 37110 19077 37174
rect 19732 37110 19796 37174
rect 20451 37110 20515 37174
rect 13980 37030 14044 37094
rect 14699 37030 14763 37094
rect 15418 37030 15482 37094
rect 16137 37030 16201 37094
rect 16856 37030 16920 37094
rect 17575 37030 17639 37094
rect 18294 37030 18358 37094
rect 19013 37030 19077 37094
rect 19732 37030 19796 37094
rect 20451 37030 20515 37094
rect 13980 36950 14044 37014
rect 14699 36950 14763 37014
rect 15418 36950 15482 37014
rect 16137 36950 16201 37014
rect 16856 36950 16920 37014
rect 17575 36950 17639 37014
rect 18294 36950 18358 37014
rect 19013 36950 19077 37014
rect 19732 36950 19796 37014
rect 20451 36950 20515 37014
rect 13980 36870 14044 36934
rect 14699 36870 14763 36934
rect 15418 36870 15482 36934
rect 16137 36870 16201 36934
rect 16856 36870 16920 36934
rect 17575 36870 17639 36934
rect 18294 36870 18358 36934
rect 19013 36870 19077 36934
rect 19732 36870 19796 36934
rect 20451 36870 20515 36934
rect 13980 36650 14044 36714
rect 14699 36650 14763 36714
rect 15418 36650 15482 36714
rect 16137 36650 16201 36714
rect 16856 36650 16920 36714
rect 17575 36650 17639 36714
rect 18294 36650 18358 36714
rect 19013 36650 19077 36714
rect 19732 36650 19796 36714
rect 20451 36650 20515 36714
rect 13980 36570 14044 36634
rect 14699 36570 14763 36634
rect 15418 36570 15482 36634
rect 16137 36570 16201 36634
rect 16856 36570 16920 36634
rect 17575 36570 17639 36634
rect 18294 36570 18358 36634
rect 19013 36570 19077 36634
rect 19732 36570 19796 36634
rect 20451 36570 20515 36634
rect 13980 36490 14044 36554
rect 14699 36490 14763 36554
rect 15418 36490 15482 36554
rect 16137 36490 16201 36554
rect 16856 36490 16920 36554
rect 17575 36490 17639 36554
rect 18294 36490 18358 36554
rect 19013 36490 19077 36554
rect 19732 36490 19796 36554
rect 20451 36490 20515 36554
rect 13980 36410 14044 36474
rect 14699 36410 14763 36474
rect 15418 36410 15482 36474
rect 16137 36410 16201 36474
rect 16856 36410 16920 36474
rect 17575 36410 17639 36474
rect 18294 36410 18358 36474
rect 19013 36410 19077 36474
rect 19732 36410 19796 36474
rect 20451 36410 20515 36474
rect 13980 36330 14044 36394
rect 14699 36330 14763 36394
rect 15418 36330 15482 36394
rect 16137 36330 16201 36394
rect 16856 36330 16920 36394
rect 17575 36330 17639 36394
rect 18294 36330 18358 36394
rect 19013 36330 19077 36394
rect 19732 36330 19796 36394
rect 20451 36330 20515 36394
rect 13980 36250 14044 36314
rect 14699 36250 14763 36314
rect 15418 36250 15482 36314
rect 16137 36250 16201 36314
rect 16856 36250 16920 36314
rect 17575 36250 17639 36314
rect 18294 36250 18358 36314
rect 19013 36250 19077 36314
rect 19732 36250 19796 36314
rect 20451 36250 20515 36314
rect 13980 36170 14044 36234
rect 14699 36170 14763 36234
rect 15418 36170 15482 36234
rect 16137 36170 16201 36234
rect 16856 36170 16920 36234
rect 17575 36170 17639 36234
rect 18294 36170 18358 36234
rect 19013 36170 19077 36234
rect 19732 36170 19796 36234
rect 20451 36170 20515 36234
rect 21428 37350 21492 37414
rect 22147 37350 22211 37414
rect 22866 37350 22930 37414
rect 23585 37350 23649 37414
rect 24304 37350 24368 37414
rect 25023 37350 25087 37414
rect 25742 37350 25806 37414
rect 26461 37350 26525 37414
rect 27180 37350 27244 37414
rect 27899 37350 27963 37414
rect 21428 37270 21492 37334
rect 22147 37270 22211 37334
rect 22866 37270 22930 37334
rect 23585 37270 23649 37334
rect 24304 37270 24368 37334
rect 25023 37270 25087 37334
rect 25742 37270 25806 37334
rect 26461 37270 26525 37334
rect 27180 37270 27244 37334
rect 27899 37270 27963 37334
rect 21428 37190 21492 37254
rect 22147 37190 22211 37254
rect 22866 37190 22930 37254
rect 23585 37190 23649 37254
rect 24304 37190 24368 37254
rect 25023 37190 25087 37254
rect 25742 37190 25806 37254
rect 26461 37190 26525 37254
rect 27180 37190 27244 37254
rect 27899 37190 27963 37254
rect 21428 37110 21492 37174
rect 22147 37110 22211 37174
rect 22866 37110 22930 37174
rect 23585 37110 23649 37174
rect 24304 37110 24368 37174
rect 25023 37110 25087 37174
rect 25742 37110 25806 37174
rect 26461 37110 26525 37174
rect 27180 37110 27244 37174
rect 27899 37110 27963 37174
rect 21428 37030 21492 37094
rect 22147 37030 22211 37094
rect 22866 37030 22930 37094
rect 23585 37030 23649 37094
rect 24304 37030 24368 37094
rect 25023 37030 25087 37094
rect 25742 37030 25806 37094
rect 26461 37030 26525 37094
rect 27180 37030 27244 37094
rect 27899 37030 27963 37094
rect 21428 36950 21492 37014
rect 22147 36950 22211 37014
rect 22866 36950 22930 37014
rect 23585 36950 23649 37014
rect 24304 36950 24368 37014
rect 25023 36950 25087 37014
rect 25742 36950 25806 37014
rect 26461 36950 26525 37014
rect 27180 36950 27244 37014
rect 27899 36950 27963 37014
rect 21428 36870 21492 36934
rect 22147 36870 22211 36934
rect 22866 36870 22930 36934
rect 23585 36870 23649 36934
rect 24304 36870 24368 36934
rect 25023 36870 25087 36934
rect 25742 36870 25806 36934
rect 26461 36870 26525 36934
rect 27180 36870 27244 36934
rect 27899 36870 27963 36934
rect 21428 36650 21492 36714
rect 22147 36650 22211 36714
rect 22866 36650 22930 36714
rect 23585 36650 23649 36714
rect 24304 36650 24368 36714
rect 25023 36650 25087 36714
rect 25742 36650 25806 36714
rect 26461 36650 26525 36714
rect 27180 36650 27244 36714
rect 27899 36650 27963 36714
rect 21428 36570 21492 36634
rect 22147 36570 22211 36634
rect 22866 36570 22930 36634
rect 23585 36570 23649 36634
rect 24304 36570 24368 36634
rect 25023 36570 25087 36634
rect 25742 36570 25806 36634
rect 26461 36570 26525 36634
rect 27180 36570 27244 36634
rect 27899 36570 27963 36634
rect 21428 36490 21492 36554
rect 22147 36490 22211 36554
rect 22866 36490 22930 36554
rect 23585 36490 23649 36554
rect 24304 36490 24368 36554
rect 25023 36490 25087 36554
rect 25742 36490 25806 36554
rect 26461 36490 26525 36554
rect 27180 36490 27244 36554
rect 27899 36490 27963 36554
rect 21428 36410 21492 36474
rect 22147 36410 22211 36474
rect 22866 36410 22930 36474
rect 23585 36410 23649 36474
rect 24304 36410 24368 36474
rect 25023 36410 25087 36474
rect 25742 36410 25806 36474
rect 26461 36410 26525 36474
rect 27180 36410 27244 36474
rect 27899 36410 27963 36474
rect 21428 36330 21492 36394
rect 22147 36330 22211 36394
rect 22866 36330 22930 36394
rect 23585 36330 23649 36394
rect 24304 36330 24368 36394
rect 25023 36330 25087 36394
rect 25742 36330 25806 36394
rect 26461 36330 26525 36394
rect 27180 36330 27244 36394
rect 27899 36330 27963 36394
rect 21428 36250 21492 36314
rect 22147 36250 22211 36314
rect 22866 36250 22930 36314
rect 23585 36250 23649 36314
rect 24304 36250 24368 36314
rect 25023 36250 25087 36314
rect 25742 36250 25806 36314
rect 26461 36250 26525 36314
rect 27180 36250 27244 36314
rect 27899 36250 27963 36314
rect 21428 36170 21492 36234
rect 22147 36170 22211 36234
rect 22866 36170 22930 36234
rect 23585 36170 23649 36234
rect 24304 36170 24368 36234
rect 25023 36170 25087 36234
rect 25742 36170 25806 36234
rect 26461 36170 26525 36234
rect 27180 36170 27244 36234
rect 27899 36170 27963 36234
rect 5946 36010 6010 36014
rect 6026 36010 6090 36014
rect 5946 35954 5990 36010
rect 5990 35954 6010 36010
rect 6026 35954 6046 36010
rect 6046 35954 6090 36010
rect 5946 35950 6010 35954
rect 6026 35950 6090 35954
rect 13394 36010 13458 36014
rect 13474 36010 13538 36014
rect 13394 35954 13438 36010
rect 13438 35954 13458 36010
rect 13474 35954 13494 36010
rect 13494 35954 13538 36010
rect 13394 35950 13458 35954
rect 13474 35950 13538 35954
rect 20842 36010 20906 36014
rect 20922 36010 20986 36014
rect 20842 35954 20886 36010
rect 20886 35954 20906 36010
rect 20922 35954 20942 36010
rect 20942 35954 20986 36010
rect 20842 35950 20906 35954
rect 20922 35950 20986 35954
rect 924 35820 988 35824
rect 924 35764 928 35820
rect 928 35764 984 35820
rect 984 35764 988 35820
rect 924 35760 988 35764
rect 1004 35820 1068 35824
rect 1004 35764 1008 35820
rect 1008 35764 1064 35820
rect 1064 35764 1068 35820
rect 1004 35760 1068 35764
rect 1084 35820 1148 35824
rect 1084 35764 1088 35820
rect 1088 35764 1144 35820
rect 1144 35764 1148 35820
rect 1084 35760 1148 35764
rect 1164 35820 1228 35824
rect 1164 35764 1168 35820
rect 1168 35764 1224 35820
rect 1224 35764 1228 35820
rect 1164 35760 1228 35764
rect 1244 35820 1308 35824
rect 1244 35764 1248 35820
rect 1248 35764 1304 35820
rect 1304 35764 1308 35820
rect 1244 35760 1308 35764
rect 1324 35820 1388 35824
rect 1324 35764 1328 35820
rect 1328 35764 1384 35820
rect 1384 35764 1388 35820
rect 1324 35760 1388 35764
rect 1404 35820 1468 35824
rect 1404 35764 1408 35820
rect 1408 35764 1464 35820
rect 1464 35764 1468 35820
rect 1404 35760 1468 35764
rect 1484 35820 1548 35824
rect 1484 35764 1488 35820
rect 1488 35764 1544 35820
rect 1544 35764 1548 35820
rect 1484 35760 1548 35764
rect 1564 35820 1628 35824
rect 1564 35764 1568 35820
rect 1568 35764 1624 35820
rect 1624 35764 1628 35820
rect 1564 35760 1628 35764
rect 1644 35820 1708 35824
rect 1644 35764 1648 35820
rect 1648 35764 1704 35820
rect 1704 35764 1708 35820
rect 1644 35760 1708 35764
rect 1724 35820 1788 35824
rect 1724 35764 1728 35820
rect 1728 35764 1784 35820
rect 1784 35764 1788 35820
rect 1724 35760 1788 35764
rect 1804 35820 1868 35824
rect 1804 35764 1808 35820
rect 1808 35764 1864 35820
rect 1864 35764 1868 35820
rect 1804 35760 1868 35764
rect 1884 35820 1948 35824
rect 1884 35764 1888 35820
rect 1888 35764 1944 35820
rect 1944 35764 1948 35820
rect 1884 35760 1948 35764
rect 1964 35820 2028 35824
rect 1964 35764 1968 35820
rect 1968 35764 2024 35820
rect 2024 35764 2028 35820
rect 1964 35760 2028 35764
rect 2044 35820 2108 35824
rect 2044 35764 2048 35820
rect 2048 35764 2104 35820
rect 2104 35764 2108 35820
rect 2044 35760 2108 35764
rect 2124 35820 2188 35824
rect 2124 35764 2128 35820
rect 2128 35764 2184 35820
rect 2184 35764 2188 35820
rect 2124 35760 2188 35764
rect 2204 35820 2268 35824
rect 2204 35764 2208 35820
rect 2208 35764 2264 35820
rect 2264 35764 2268 35820
rect 2204 35760 2268 35764
rect 2284 35820 2348 35824
rect 2284 35764 2288 35820
rect 2288 35764 2344 35820
rect 2344 35764 2348 35820
rect 2284 35760 2348 35764
rect 2364 35820 2428 35824
rect 2364 35764 2368 35820
rect 2368 35764 2424 35820
rect 2424 35764 2428 35820
rect 2364 35760 2428 35764
rect 2444 35820 2508 35824
rect 2444 35764 2448 35820
rect 2448 35764 2504 35820
rect 2504 35764 2508 35820
rect 2444 35760 2508 35764
rect 46128 35820 46192 35824
rect 46128 35764 46132 35820
rect 46132 35764 46188 35820
rect 46188 35764 46192 35820
rect 46128 35760 46192 35764
rect 46208 35820 46272 35824
rect 46208 35764 46212 35820
rect 46212 35764 46268 35820
rect 46268 35764 46272 35820
rect 46208 35760 46272 35764
rect 46288 35820 46352 35824
rect 46288 35764 46292 35820
rect 46292 35764 46348 35820
rect 46348 35764 46352 35820
rect 46288 35760 46352 35764
rect 46368 35820 46432 35824
rect 46368 35764 46372 35820
rect 46372 35764 46428 35820
rect 46428 35764 46432 35820
rect 46368 35760 46432 35764
rect 46448 35820 46512 35824
rect 46448 35764 46452 35820
rect 46452 35764 46508 35820
rect 46508 35764 46512 35820
rect 46448 35760 46512 35764
rect 46528 35820 46592 35824
rect 46528 35764 46532 35820
rect 46532 35764 46588 35820
rect 46588 35764 46592 35820
rect 46528 35760 46592 35764
rect 46608 35820 46672 35824
rect 46608 35764 46612 35820
rect 46612 35764 46668 35820
rect 46668 35764 46672 35820
rect 46608 35760 46672 35764
rect 46688 35820 46752 35824
rect 46688 35764 46692 35820
rect 46692 35764 46748 35820
rect 46748 35764 46752 35820
rect 46688 35760 46752 35764
rect 46768 35820 46832 35824
rect 46768 35764 46772 35820
rect 46772 35764 46828 35820
rect 46828 35764 46832 35820
rect 46768 35760 46832 35764
rect 46848 35820 46912 35824
rect 46848 35764 46852 35820
rect 46852 35764 46908 35820
rect 46908 35764 46912 35820
rect 46848 35760 46912 35764
rect 46928 35820 46992 35824
rect 46928 35764 46932 35820
rect 46932 35764 46988 35820
rect 46988 35764 46992 35820
rect 46928 35760 46992 35764
rect 47008 35820 47072 35824
rect 47008 35764 47012 35820
rect 47012 35764 47068 35820
rect 47068 35764 47072 35820
rect 47008 35760 47072 35764
rect 47088 35820 47152 35824
rect 47088 35764 47092 35820
rect 47092 35764 47148 35820
rect 47148 35764 47152 35820
rect 47088 35760 47152 35764
rect 47168 35820 47232 35824
rect 47168 35764 47172 35820
rect 47172 35764 47228 35820
rect 47228 35764 47232 35820
rect 47168 35760 47232 35764
rect 47248 35820 47312 35824
rect 47248 35764 47252 35820
rect 47252 35764 47308 35820
rect 47308 35764 47312 35820
rect 47248 35760 47312 35764
rect 47328 35820 47392 35824
rect 47328 35764 47332 35820
rect 47332 35764 47388 35820
rect 47388 35764 47392 35820
rect 47328 35760 47392 35764
rect 47408 35820 47472 35824
rect 47408 35764 47412 35820
rect 47412 35764 47468 35820
rect 47468 35764 47472 35820
rect 47408 35760 47472 35764
rect 47488 35820 47552 35824
rect 47488 35764 47492 35820
rect 47492 35764 47548 35820
rect 47548 35764 47552 35820
rect 47488 35760 47552 35764
rect 47568 35820 47632 35824
rect 47568 35764 47572 35820
rect 47572 35764 47628 35820
rect 47628 35764 47632 35820
rect 47568 35760 47632 35764
rect 47648 35820 47712 35824
rect 47648 35764 47652 35820
rect 47652 35764 47708 35820
rect 47708 35764 47712 35820
rect 47648 35760 47712 35764
rect 3372 33940 3436 33944
rect 3372 33884 3376 33940
rect 3376 33884 3432 33940
rect 3432 33884 3436 33940
rect 3372 33880 3436 33884
rect 3452 33940 3516 33944
rect 3452 33884 3456 33940
rect 3456 33884 3512 33940
rect 3512 33884 3516 33940
rect 3452 33880 3516 33884
rect 3532 33940 3596 33944
rect 3532 33884 3536 33940
rect 3536 33884 3592 33940
rect 3592 33884 3596 33940
rect 3532 33880 3596 33884
rect 3612 33940 3676 33944
rect 3612 33884 3616 33940
rect 3616 33884 3672 33940
rect 3672 33884 3676 33940
rect 3612 33880 3676 33884
rect 3692 33940 3756 33944
rect 3692 33884 3696 33940
rect 3696 33884 3752 33940
rect 3752 33884 3756 33940
rect 3692 33880 3756 33884
rect 3772 33940 3836 33944
rect 3772 33884 3776 33940
rect 3776 33884 3832 33940
rect 3832 33884 3836 33940
rect 3772 33880 3836 33884
rect 3852 33940 3916 33944
rect 3852 33884 3856 33940
rect 3856 33884 3912 33940
rect 3912 33884 3916 33940
rect 3852 33880 3916 33884
rect 3932 33940 3996 33944
rect 3932 33884 3936 33940
rect 3936 33884 3992 33940
rect 3992 33884 3996 33940
rect 3932 33880 3996 33884
rect 4012 33940 4076 33944
rect 4012 33884 4016 33940
rect 4016 33884 4072 33940
rect 4072 33884 4076 33940
rect 4012 33880 4076 33884
rect 4092 33940 4156 33944
rect 4092 33884 4096 33940
rect 4096 33884 4152 33940
rect 4152 33884 4156 33940
rect 4092 33880 4156 33884
rect 4172 33940 4236 33944
rect 4172 33884 4176 33940
rect 4176 33884 4232 33940
rect 4232 33884 4236 33940
rect 4172 33880 4236 33884
rect 4252 33940 4316 33944
rect 4252 33884 4256 33940
rect 4256 33884 4312 33940
rect 4312 33884 4316 33940
rect 4252 33880 4316 33884
rect 4332 33940 4396 33944
rect 4332 33884 4336 33940
rect 4336 33884 4392 33940
rect 4392 33884 4396 33940
rect 4332 33880 4396 33884
rect 4412 33940 4476 33944
rect 4412 33884 4416 33940
rect 4416 33884 4472 33940
rect 4472 33884 4476 33940
rect 4412 33880 4476 33884
rect 4492 33940 4556 33944
rect 4492 33884 4496 33940
rect 4496 33884 4552 33940
rect 4552 33884 4556 33940
rect 4492 33880 4556 33884
rect 4572 33940 4636 33944
rect 4572 33884 4576 33940
rect 4576 33884 4632 33940
rect 4632 33884 4636 33940
rect 4572 33880 4636 33884
rect 4652 33940 4716 33944
rect 4652 33884 4656 33940
rect 4656 33884 4712 33940
rect 4712 33884 4716 33940
rect 4652 33880 4716 33884
rect 4732 33940 4796 33944
rect 4732 33884 4736 33940
rect 4736 33884 4792 33940
rect 4792 33884 4796 33940
rect 4732 33880 4796 33884
rect 4812 33940 4876 33944
rect 4812 33884 4816 33940
rect 4816 33884 4872 33940
rect 4872 33884 4876 33940
rect 4812 33880 4876 33884
rect 4892 33940 4956 33944
rect 4892 33884 4896 33940
rect 4896 33884 4952 33940
rect 4952 33884 4956 33940
rect 4892 33880 4956 33884
rect 43680 33940 43744 33944
rect 43680 33884 43684 33940
rect 43684 33884 43740 33940
rect 43740 33884 43744 33940
rect 43680 33880 43744 33884
rect 43760 33940 43824 33944
rect 43760 33884 43764 33940
rect 43764 33884 43820 33940
rect 43820 33884 43824 33940
rect 43760 33880 43824 33884
rect 43840 33940 43904 33944
rect 43840 33884 43844 33940
rect 43844 33884 43900 33940
rect 43900 33884 43904 33940
rect 43840 33880 43904 33884
rect 43920 33940 43984 33944
rect 43920 33884 43924 33940
rect 43924 33884 43980 33940
rect 43980 33884 43984 33940
rect 43920 33880 43984 33884
rect 44000 33940 44064 33944
rect 44000 33884 44004 33940
rect 44004 33884 44060 33940
rect 44060 33884 44064 33940
rect 44000 33880 44064 33884
rect 44080 33940 44144 33944
rect 44080 33884 44084 33940
rect 44084 33884 44140 33940
rect 44140 33884 44144 33940
rect 44080 33880 44144 33884
rect 44160 33940 44224 33944
rect 44160 33884 44164 33940
rect 44164 33884 44220 33940
rect 44220 33884 44224 33940
rect 44160 33880 44224 33884
rect 44240 33940 44304 33944
rect 44240 33884 44244 33940
rect 44244 33884 44300 33940
rect 44300 33884 44304 33940
rect 44240 33880 44304 33884
rect 44320 33940 44384 33944
rect 44320 33884 44324 33940
rect 44324 33884 44380 33940
rect 44380 33884 44384 33940
rect 44320 33880 44384 33884
rect 44400 33940 44464 33944
rect 44400 33884 44404 33940
rect 44404 33884 44460 33940
rect 44460 33884 44464 33940
rect 44400 33880 44464 33884
rect 44480 33940 44544 33944
rect 44480 33884 44484 33940
rect 44484 33884 44540 33940
rect 44540 33884 44544 33940
rect 44480 33880 44544 33884
rect 44560 33940 44624 33944
rect 44560 33884 44564 33940
rect 44564 33884 44620 33940
rect 44620 33884 44624 33940
rect 44560 33880 44624 33884
rect 44640 33940 44704 33944
rect 44640 33884 44644 33940
rect 44644 33884 44700 33940
rect 44700 33884 44704 33940
rect 44640 33880 44704 33884
rect 44720 33940 44784 33944
rect 44720 33884 44724 33940
rect 44724 33884 44780 33940
rect 44780 33884 44784 33940
rect 44720 33880 44784 33884
rect 44800 33940 44864 33944
rect 44800 33884 44804 33940
rect 44804 33884 44860 33940
rect 44860 33884 44864 33940
rect 44800 33880 44864 33884
rect 44880 33940 44944 33944
rect 44880 33884 44884 33940
rect 44884 33884 44940 33940
rect 44940 33884 44944 33940
rect 44880 33880 44944 33884
rect 44960 33940 45024 33944
rect 44960 33884 44964 33940
rect 44964 33884 45020 33940
rect 45020 33884 45024 33940
rect 44960 33880 45024 33884
rect 45040 33940 45104 33944
rect 45040 33884 45044 33940
rect 45044 33884 45100 33940
rect 45100 33884 45104 33940
rect 45040 33880 45104 33884
rect 45120 33940 45184 33944
rect 45120 33884 45124 33940
rect 45124 33884 45180 33940
rect 45180 33884 45184 33940
rect 45120 33880 45184 33884
rect 45200 33940 45264 33944
rect 45200 33884 45204 33940
rect 45204 33884 45260 33940
rect 45260 33884 45264 33940
rect 45200 33880 45264 33884
rect 10088 33774 10152 33838
rect 7218 33590 7282 33654
rect 7937 33590 8001 33654
rect 8656 33590 8720 33654
rect 9375 33590 9439 33654
rect 10094 33590 10158 33654
rect 10813 33590 10877 33654
rect 11532 33590 11596 33654
rect 12251 33590 12315 33654
rect 12970 33590 13034 33654
rect 13689 33590 13753 33654
rect 7218 33510 7282 33574
rect 7937 33510 8001 33574
rect 8656 33510 8720 33574
rect 9375 33510 9439 33574
rect 10094 33510 10158 33574
rect 10813 33510 10877 33574
rect 11532 33510 11596 33574
rect 12251 33510 12315 33574
rect 12970 33510 13034 33574
rect 13689 33510 13753 33574
rect 7218 33430 7282 33494
rect 7937 33430 8001 33494
rect 8656 33430 8720 33494
rect 9375 33430 9439 33494
rect 10094 33430 10158 33494
rect 10813 33430 10877 33494
rect 11532 33430 11596 33494
rect 12251 33430 12315 33494
rect 12970 33430 13034 33494
rect 13689 33430 13753 33494
rect 7218 33350 7282 33414
rect 7937 33350 8001 33414
rect 8656 33350 8720 33414
rect 9375 33350 9439 33414
rect 10094 33350 10158 33414
rect 10813 33350 10877 33414
rect 11532 33350 11596 33414
rect 12251 33350 12315 33414
rect 12970 33350 13034 33414
rect 13689 33350 13753 33414
rect 7218 33270 7282 33334
rect 7937 33270 8001 33334
rect 8656 33270 8720 33334
rect 9375 33270 9439 33334
rect 10094 33270 10158 33334
rect 10813 33270 10877 33334
rect 11532 33270 11596 33334
rect 12251 33270 12315 33334
rect 12970 33270 13034 33334
rect 13689 33270 13753 33334
rect 7218 33190 7282 33254
rect 7937 33190 8001 33254
rect 8656 33190 8720 33254
rect 9375 33190 9439 33254
rect 10094 33190 10158 33254
rect 10813 33190 10877 33254
rect 11532 33190 11596 33254
rect 12251 33190 12315 33254
rect 12970 33190 13034 33254
rect 13689 33190 13753 33254
rect 7218 33110 7282 33174
rect 7937 33110 8001 33174
rect 8656 33110 8720 33174
rect 9375 33110 9439 33174
rect 10094 33110 10158 33174
rect 10813 33110 10877 33174
rect 11532 33110 11596 33174
rect 12251 33110 12315 33174
rect 12970 33110 13034 33174
rect 13689 33110 13753 33174
rect 7218 32890 7282 32954
rect 7937 32890 8001 32954
rect 8656 32890 8720 32954
rect 9375 32890 9439 32954
rect 10094 32890 10158 32954
rect 10813 32890 10877 32954
rect 11532 32890 11596 32954
rect 12251 32890 12315 32954
rect 12970 32890 13034 32954
rect 13689 32890 13753 32954
rect 7218 32810 7282 32874
rect 7937 32810 8001 32874
rect 8656 32810 8720 32874
rect 9375 32810 9439 32874
rect 10094 32810 10158 32874
rect 10813 32810 10877 32874
rect 11532 32810 11596 32874
rect 12251 32810 12315 32874
rect 12970 32810 13034 32874
rect 13689 32810 13753 32874
rect 7218 32730 7282 32794
rect 7937 32730 8001 32794
rect 8656 32730 8720 32794
rect 9375 32730 9439 32794
rect 10094 32730 10158 32794
rect 10813 32730 10877 32794
rect 11532 32730 11596 32794
rect 12251 32730 12315 32794
rect 12970 32730 13034 32794
rect 13689 32730 13753 32794
rect 7218 32650 7282 32714
rect 7937 32650 8001 32714
rect 8656 32650 8720 32714
rect 9375 32650 9439 32714
rect 10094 32650 10158 32714
rect 10813 32650 10877 32714
rect 11532 32650 11596 32714
rect 12251 32650 12315 32714
rect 12970 32650 13034 32714
rect 13689 32650 13753 32714
rect 7218 32570 7282 32634
rect 7937 32570 8001 32634
rect 8656 32570 8720 32634
rect 9375 32570 9439 32634
rect 10094 32570 10158 32634
rect 10813 32570 10877 32634
rect 11532 32570 11596 32634
rect 12251 32570 12315 32634
rect 12970 32570 13034 32634
rect 13689 32570 13753 32634
rect 7218 32490 7282 32554
rect 7937 32490 8001 32554
rect 8656 32490 8720 32554
rect 9375 32490 9439 32554
rect 10094 32490 10158 32554
rect 10813 32490 10877 32554
rect 11532 32490 11596 32554
rect 12251 32490 12315 32554
rect 12970 32490 13034 32554
rect 13689 32490 13753 32554
rect 7218 32410 7282 32474
rect 7937 32410 8001 32474
rect 8656 32410 8720 32474
rect 9375 32410 9439 32474
rect 10094 32410 10158 32474
rect 10813 32410 10877 32474
rect 11532 32410 11596 32474
rect 12251 32410 12315 32474
rect 12970 32410 13034 32474
rect 13689 32410 13753 32474
rect 6632 32250 6696 32254
rect 6712 32250 6776 32254
rect 6632 32194 6676 32250
rect 6676 32194 6696 32250
rect 6712 32194 6732 32250
rect 6732 32194 6776 32250
rect 6632 32190 6696 32194
rect 6712 32190 6776 32194
rect 13538 32188 13602 32252
rect 924 32060 988 32064
rect 924 32004 928 32060
rect 928 32004 984 32060
rect 984 32004 988 32060
rect 924 32000 988 32004
rect 1004 32060 1068 32064
rect 1004 32004 1008 32060
rect 1008 32004 1064 32060
rect 1064 32004 1068 32060
rect 1004 32000 1068 32004
rect 1084 32060 1148 32064
rect 1084 32004 1088 32060
rect 1088 32004 1144 32060
rect 1144 32004 1148 32060
rect 1084 32000 1148 32004
rect 1164 32060 1228 32064
rect 1164 32004 1168 32060
rect 1168 32004 1224 32060
rect 1224 32004 1228 32060
rect 1164 32000 1228 32004
rect 1244 32060 1308 32064
rect 1244 32004 1248 32060
rect 1248 32004 1304 32060
rect 1304 32004 1308 32060
rect 1244 32000 1308 32004
rect 1324 32060 1388 32064
rect 1324 32004 1328 32060
rect 1328 32004 1384 32060
rect 1384 32004 1388 32060
rect 1324 32000 1388 32004
rect 1404 32060 1468 32064
rect 1404 32004 1408 32060
rect 1408 32004 1464 32060
rect 1464 32004 1468 32060
rect 1404 32000 1468 32004
rect 1484 32060 1548 32064
rect 1484 32004 1488 32060
rect 1488 32004 1544 32060
rect 1544 32004 1548 32060
rect 1484 32000 1548 32004
rect 1564 32060 1628 32064
rect 1564 32004 1568 32060
rect 1568 32004 1624 32060
rect 1624 32004 1628 32060
rect 1564 32000 1628 32004
rect 1644 32060 1708 32064
rect 1644 32004 1648 32060
rect 1648 32004 1704 32060
rect 1704 32004 1708 32060
rect 1644 32000 1708 32004
rect 1724 32060 1788 32064
rect 1724 32004 1728 32060
rect 1728 32004 1784 32060
rect 1784 32004 1788 32060
rect 1724 32000 1788 32004
rect 1804 32060 1868 32064
rect 1804 32004 1808 32060
rect 1808 32004 1864 32060
rect 1864 32004 1868 32060
rect 1804 32000 1868 32004
rect 1884 32060 1948 32064
rect 1884 32004 1888 32060
rect 1888 32004 1944 32060
rect 1944 32004 1948 32060
rect 1884 32000 1948 32004
rect 1964 32060 2028 32064
rect 1964 32004 1968 32060
rect 1968 32004 2024 32060
rect 2024 32004 2028 32060
rect 1964 32000 2028 32004
rect 2044 32060 2108 32064
rect 2044 32004 2048 32060
rect 2048 32004 2104 32060
rect 2104 32004 2108 32060
rect 2044 32000 2108 32004
rect 2124 32060 2188 32064
rect 2124 32004 2128 32060
rect 2128 32004 2184 32060
rect 2184 32004 2188 32060
rect 2124 32000 2188 32004
rect 2204 32060 2268 32064
rect 2204 32004 2208 32060
rect 2208 32004 2264 32060
rect 2264 32004 2268 32060
rect 2204 32000 2268 32004
rect 2284 32060 2348 32064
rect 2284 32004 2288 32060
rect 2288 32004 2344 32060
rect 2344 32004 2348 32060
rect 2284 32000 2348 32004
rect 2364 32060 2428 32064
rect 2364 32004 2368 32060
rect 2368 32004 2424 32060
rect 2424 32004 2428 32060
rect 2364 32000 2428 32004
rect 2444 32060 2508 32064
rect 2444 32004 2448 32060
rect 2448 32004 2504 32060
rect 2504 32004 2508 32060
rect 2444 32000 2508 32004
rect 46128 32060 46192 32064
rect 46128 32004 46132 32060
rect 46132 32004 46188 32060
rect 46188 32004 46192 32060
rect 46128 32000 46192 32004
rect 46208 32060 46272 32064
rect 46208 32004 46212 32060
rect 46212 32004 46268 32060
rect 46268 32004 46272 32060
rect 46208 32000 46272 32004
rect 46288 32060 46352 32064
rect 46288 32004 46292 32060
rect 46292 32004 46348 32060
rect 46348 32004 46352 32060
rect 46288 32000 46352 32004
rect 46368 32060 46432 32064
rect 46368 32004 46372 32060
rect 46372 32004 46428 32060
rect 46428 32004 46432 32060
rect 46368 32000 46432 32004
rect 46448 32060 46512 32064
rect 46448 32004 46452 32060
rect 46452 32004 46508 32060
rect 46508 32004 46512 32060
rect 46448 32000 46512 32004
rect 46528 32060 46592 32064
rect 46528 32004 46532 32060
rect 46532 32004 46588 32060
rect 46588 32004 46592 32060
rect 46528 32000 46592 32004
rect 46608 32060 46672 32064
rect 46608 32004 46612 32060
rect 46612 32004 46668 32060
rect 46668 32004 46672 32060
rect 46608 32000 46672 32004
rect 46688 32060 46752 32064
rect 46688 32004 46692 32060
rect 46692 32004 46748 32060
rect 46748 32004 46752 32060
rect 46688 32000 46752 32004
rect 46768 32060 46832 32064
rect 46768 32004 46772 32060
rect 46772 32004 46828 32060
rect 46828 32004 46832 32060
rect 46768 32000 46832 32004
rect 46848 32060 46912 32064
rect 46848 32004 46852 32060
rect 46852 32004 46908 32060
rect 46908 32004 46912 32060
rect 46848 32000 46912 32004
rect 46928 32060 46992 32064
rect 46928 32004 46932 32060
rect 46932 32004 46988 32060
rect 46988 32004 46992 32060
rect 46928 32000 46992 32004
rect 47008 32060 47072 32064
rect 47008 32004 47012 32060
rect 47012 32004 47068 32060
rect 47068 32004 47072 32060
rect 47008 32000 47072 32004
rect 47088 32060 47152 32064
rect 47088 32004 47092 32060
rect 47092 32004 47148 32060
rect 47148 32004 47152 32060
rect 47088 32000 47152 32004
rect 47168 32060 47232 32064
rect 47168 32004 47172 32060
rect 47172 32004 47228 32060
rect 47228 32004 47232 32060
rect 47168 32000 47232 32004
rect 47248 32060 47312 32064
rect 47248 32004 47252 32060
rect 47252 32004 47308 32060
rect 47308 32004 47312 32060
rect 47248 32000 47312 32004
rect 47328 32060 47392 32064
rect 47328 32004 47332 32060
rect 47332 32004 47388 32060
rect 47388 32004 47392 32060
rect 47328 32000 47392 32004
rect 47408 32060 47472 32064
rect 47408 32004 47412 32060
rect 47412 32004 47468 32060
rect 47468 32004 47472 32060
rect 47408 32000 47472 32004
rect 47488 32060 47552 32064
rect 47488 32004 47492 32060
rect 47492 32004 47548 32060
rect 47548 32004 47552 32060
rect 47488 32000 47552 32004
rect 47568 32060 47632 32064
rect 47568 32004 47572 32060
rect 47572 32004 47628 32060
rect 47628 32004 47632 32060
rect 47568 32000 47632 32004
rect 47648 32060 47712 32064
rect 47648 32004 47652 32060
rect 47652 32004 47708 32060
rect 47708 32004 47712 32060
rect 47648 32000 47712 32004
rect 3372 30180 3436 30184
rect 3372 30124 3376 30180
rect 3376 30124 3432 30180
rect 3432 30124 3436 30180
rect 3372 30120 3436 30124
rect 3452 30180 3516 30184
rect 3452 30124 3456 30180
rect 3456 30124 3512 30180
rect 3512 30124 3516 30180
rect 3452 30120 3516 30124
rect 3532 30180 3596 30184
rect 3532 30124 3536 30180
rect 3536 30124 3592 30180
rect 3592 30124 3596 30180
rect 3532 30120 3596 30124
rect 3612 30180 3676 30184
rect 3612 30124 3616 30180
rect 3616 30124 3672 30180
rect 3672 30124 3676 30180
rect 3612 30120 3676 30124
rect 3692 30180 3756 30184
rect 3692 30124 3696 30180
rect 3696 30124 3752 30180
rect 3752 30124 3756 30180
rect 3692 30120 3756 30124
rect 3772 30180 3836 30184
rect 3772 30124 3776 30180
rect 3776 30124 3832 30180
rect 3832 30124 3836 30180
rect 3772 30120 3836 30124
rect 3852 30180 3916 30184
rect 3852 30124 3856 30180
rect 3856 30124 3912 30180
rect 3912 30124 3916 30180
rect 3852 30120 3916 30124
rect 3932 30180 3996 30184
rect 3932 30124 3936 30180
rect 3936 30124 3992 30180
rect 3992 30124 3996 30180
rect 3932 30120 3996 30124
rect 4012 30180 4076 30184
rect 4012 30124 4016 30180
rect 4016 30124 4072 30180
rect 4072 30124 4076 30180
rect 4012 30120 4076 30124
rect 4092 30180 4156 30184
rect 4092 30124 4096 30180
rect 4096 30124 4152 30180
rect 4152 30124 4156 30180
rect 4092 30120 4156 30124
rect 4172 30180 4236 30184
rect 4172 30124 4176 30180
rect 4176 30124 4232 30180
rect 4232 30124 4236 30180
rect 4172 30120 4236 30124
rect 4252 30180 4316 30184
rect 4252 30124 4256 30180
rect 4256 30124 4312 30180
rect 4312 30124 4316 30180
rect 4252 30120 4316 30124
rect 4332 30180 4396 30184
rect 4332 30124 4336 30180
rect 4336 30124 4392 30180
rect 4392 30124 4396 30180
rect 4332 30120 4396 30124
rect 4412 30180 4476 30184
rect 4412 30124 4416 30180
rect 4416 30124 4472 30180
rect 4472 30124 4476 30180
rect 4412 30120 4476 30124
rect 4492 30180 4556 30184
rect 4492 30124 4496 30180
rect 4496 30124 4552 30180
rect 4552 30124 4556 30180
rect 4492 30120 4556 30124
rect 4572 30180 4636 30184
rect 4572 30124 4576 30180
rect 4576 30124 4632 30180
rect 4632 30124 4636 30180
rect 4572 30120 4636 30124
rect 4652 30180 4716 30184
rect 4652 30124 4656 30180
rect 4656 30124 4712 30180
rect 4712 30124 4716 30180
rect 4652 30120 4716 30124
rect 4732 30180 4796 30184
rect 4732 30124 4736 30180
rect 4736 30124 4792 30180
rect 4792 30124 4796 30180
rect 4732 30120 4796 30124
rect 4812 30180 4876 30184
rect 4812 30124 4816 30180
rect 4816 30124 4872 30180
rect 4872 30124 4876 30180
rect 4812 30120 4876 30124
rect 4892 30180 4956 30184
rect 4892 30124 4896 30180
rect 4896 30124 4952 30180
rect 4952 30124 4956 30180
rect 4892 30120 4956 30124
rect 43680 30180 43744 30184
rect 43680 30124 43684 30180
rect 43684 30124 43740 30180
rect 43740 30124 43744 30180
rect 43680 30120 43744 30124
rect 43760 30180 43824 30184
rect 43760 30124 43764 30180
rect 43764 30124 43820 30180
rect 43820 30124 43824 30180
rect 43760 30120 43824 30124
rect 43840 30180 43904 30184
rect 43840 30124 43844 30180
rect 43844 30124 43900 30180
rect 43900 30124 43904 30180
rect 43840 30120 43904 30124
rect 43920 30180 43984 30184
rect 43920 30124 43924 30180
rect 43924 30124 43980 30180
rect 43980 30124 43984 30180
rect 43920 30120 43984 30124
rect 44000 30180 44064 30184
rect 44000 30124 44004 30180
rect 44004 30124 44060 30180
rect 44060 30124 44064 30180
rect 44000 30120 44064 30124
rect 44080 30180 44144 30184
rect 44080 30124 44084 30180
rect 44084 30124 44140 30180
rect 44140 30124 44144 30180
rect 44080 30120 44144 30124
rect 44160 30180 44224 30184
rect 44160 30124 44164 30180
rect 44164 30124 44220 30180
rect 44220 30124 44224 30180
rect 44160 30120 44224 30124
rect 44240 30180 44304 30184
rect 44240 30124 44244 30180
rect 44244 30124 44300 30180
rect 44300 30124 44304 30180
rect 44240 30120 44304 30124
rect 44320 30180 44384 30184
rect 44320 30124 44324 30180
rect 44324 30124 44380 30180
rect 44380 30124 44384 30180
rect 44320 30120 44384 30124
rect 44400 30180 44464 30184
rect 44400 30124 44404 30180
rect 44404 30124 44460 30180
rect 44460 30124 44464 30180
rect 44400 30120 44464 30124
rect 44480 30180 44544 30184
rect 44480 30124 44484 30180
rect 44484 30124 44540 30180
rect 44540 30124 44544 30180
rect 44480 30120 44544 30124
rect 44560 30180 44624 30184
rect 44560 30124 44564 30180
rect 44564 30124 44620 30180
rect 44620 30124 44624 30180
rect 44560 30120 44624 30124
rect 44640 30180 44704 30184
rect 44640 30124 44644 30180
rect 44644 30124 44700 30180
rect 44700 30124 44704 30180
rect 44640 30120 44704 30124
rect 44720 30180 44784 30184
rect 44720 30124 44724 30180
rect 44724 30124 44780 30180
rect 44780 30124 44784 30180
rect 44720 30120 44784 30124
rect 44800 30180 44864 30184
rect 44800 30124 44804 30180
rect 44804 30124 44860 30180
rect 44860 30124 44864 30180
rect 44800 30120 44864 30124
rect 44880 30180 44944 30184
rect 44880 30124 44884 30180
rect 44884 30124 44940 30180
rect 44940 30124 44944 30180
rect 44880 30120 44944 30124
rect 44960 30180 45024 30184
rect 44960 30124 44964 30180
rect 44964 30124 45020 30180
rect 45020 30124 45024 30180
rect 44960 30120 45024 30124
rect 45040 30180 45104 30184
rect 45040 30124 45044 30180
rect 45044 30124 45100 30180
rect 45100 30124 45104 30180
rect 45040 30120 45104 30124
rect 45120 30180 45184 30184
rect 45120 30124 45124 30180
rect 45124 30124 45180 30180
rect 45180 30124 45184 30180
rect 45120 30120 45184 30124
rect 45200 30180 45264 30184
rect 45200 30124 45204 30180
rect 45204 30124 45260 30180
rect 45260 30124 45264 30180
rect 45200 30120 45264 30124
rect 18920 28588 18984 28592
rect 18920 28532 18934 28588
rect 18934 28532 18984 28588
rect 18920 28528 18984 28532
rect 924 28300 988 28304
rect 924 28244 928 28300
rect 928 28244 984 28300
rect 984 28244 988 28300
rect 924 28240 988 28244
rect 1004 28300 1068 28304
rect 1004 28244 1008 28300
rect 1008 28244 1064 28300
rect 1064 28244 1068 28300
rect 1004 28240 1068 28244
rect 1084 28300 1148 28304
rect 1084 28244 1088 28300
rect 1088 28244 1144 28300
rect 1144 28244 1148 28300
rect 1084 28240 1148 28244
rect 1164 28300 1228 28304
rect 1164 28244 1168 28300
rect 1168 28244 1224 28300
rect 1224 28244 1228 28300
rect 1164 28240 1228 28244
rect 1244 28300 1308 28304
rect 1244 28244 1248 28300
rect 1248 28244 1304 28300
rect 1304 28244 1308 28300
rect 1244 28240 1308 28244
rect 1324 28300 1388 28304
rect 1324 28244 1328 28300
rect 1328 28244 1384 28300
rect 1384 28244 1388 28300
rect 1324 28240 1388 28244
rect 1404 28300 1468 28304
rect 1404 28244 1408 28300
rect 1408 28244 1464 28300
rect 1464 28244 1468 28300
rect 1404 28240 1468 28244
rect 1484 28300 1548 28304
rect 1484 28244 1488 28300
rect 1488 28244 1544 28300
rect 1544 28244 1548 28300
rect 1484 28240 1548 28244
rect 1564 28300 1628 28304
rect 1564 28244 1568 28300
rect 1568 28244 1624 28300
rect 1624 28244 1628 28300
rect 1564 28240 1628 28244
rect 1644 28300 1708 28304
rect 1644 28244 1648 28300
rect 1648 28244 1704 28300
rect 1704 28244 1708 28300
rect 1644 28240 1708 28244
rect 1724 28300 1788 28304
rect 1724 28244 1728 28300
rect 1728 28244 1784 28300
rect 1784 28244 1788 28300
rect 1724 28240 1788 28244
rect 1804 28300 1868 28304
rect 1804 28244 1808 28300
rect 1808 28244 1864 28300
rect 1864 28244 1868 28300
rect 1804 28240 1868 28244
rect 1884 28300 1948 28304
rect 1884 28244 1888 28300
rect 1888 28244 1944 28300
rect 1944 28244 1948 28300
rect 1884 28240 1948 28244
rect 1964 28300 2028 28304
rect 1964 28244 1968 28300
rect 1968 28244 2024 28300
rect 2024 28244 2028 28300
rect 1964 28240 2028 28244
rect 2044 28300 2108 28304
rect 2044 28244 2048 28300
rect 2048 28244 2104 28300
rect 2104 28244 2108 28300
rect 2044 28240 2108 28244
rect 2124 28300 2188 28304
rect 2124 28244 2128 28300
rect 2128 28244 2184 28300
rect 2184 28244 2188 28300
rect 2124 28240 2188 28244
rect 2204 28300 2268 28304
rect 2204 28244 2208 28300
rect 2208 28244 2264 28300
rect 2264 28244 2268 28300
rect 2204 28240 2268 28244
rect 2284 28300 2348 28304
rect 2284 28244 2288 28300
rect 2288 28244 2344 28300
rect 2344 28244 2348 28300
rect 2284 28240 2348 28244
rect 2364 28300 2428 28304
rect 2364 28244 2368 28300
rect 2368 28244 2424 28300
rect 2424 28244 2428 28300
rect 2364 28240 2428 28244
rect 2444 28300 2508 28304
rect 2444 28244 2448 28300
rect 2448 28244 2504 28300
rect 2504 28244 2508 28300
rect 2444 28240 2508 28244
rect 46128 28300 46192 28304
rect 46128 28244 46132 28300
rect 46132 28244 46188 28300
rect 46188 28244 46192 28300
rect 46128 28240 46192 28244
rect 46208 28300 46272 28304
rect 46208 28244 46212 28300
rect 46212 28244 46268 28300
rect 46268 28244 46272 28300
rect 46208 28240 46272 28244
rect 46288 28300 46352 28304
rect 46288 28244 46292 28300
rect 46292 28244 46348 28300
rect 46348 28244 46352 28300
rect 46288 28240 46352 28244
rect 46368 28300 46432 28304
rect 46368 28244 46372 28300
rect 46372 28244 46428 28300
rect 46428 28244 46432 28300
rect 46368 28240 46432 28244
rect 46448 28300 46512 28304
rect 46448 28244 46452 28300
rect 46452 28244 46508 28300
rect 46508 28244 46512 28300
rect 46448 28240 46512 28244
rect 46528 28300 46592 28304
rect 46528 28244 46532 28300
rect 46532 28244 46588 28300
rect 46588 28244 46592 28300
rect 46528 28240 46592 28244
rect 46608 28300 46672 28304
rect 46608 28244 46612 28300
rect 46612 28244 46668 28300
rect 46668 28244 46672 28300
rect 46608 28240 46672 28244
rect 46688 28300 46752 28304
rect 46688 28244 46692 28300
rect 46692 28244 46748 28300
rect 46748 28244 46752 28300
rect 46688 28240 46752 28244
rect 46768 28300 46832 28304
rect 46768 28244 46772 28300
rect 46772 28244 46828 28300
rect 46828 28244 46832 28300
rect 46768 28240 46832 28244
rect 46848 28300 46912 28304
rect 46848 28244 46852 28300
rect 46852 28244 46908 28300
rect 46908 28244 46912 28300
rect 46848 28240 46912 28244
rect 46928 28300 46992 28304
rect 46928 28244 46932 28300
rect 46932 28244 46988 28300
rect 46988 28244 46992 28300
rect 46928 28240 46992 28244
rect 47008 28300 47072 28304
rect 47008 28244 47012 28300
rect 47012 28244 47068 28300
rect 47068 28244 47072 28300
rect 47008 28240 47072 28244
rect 47088 28300 47152 28304
rect 47088 28244 47092 28300
rect 47092 28244 47148 28300
rect 47148 28244 47152 28300
rect 47088 28240 47152 28244
rect 47168 28300 47232 28304
rect 47168 28244 47172 28300
rect 47172 28244 47228 28300
rect 47228 28244 47232 28300
rect 47168 28240 47232 28244
rect 47248 28300 47312 28304
rect 47248 28244 47252 28300
rect 47252 28244 47308 28300
rect 47308 28244 47312 28300
rect 47248 28240 47312 28244
rect 47328 28300 47392 28304
rect 47328 28244 47332 28300
rect 47332 28244 47388 28300
rect 47388 28244 47392 28300
rect 47328 28240 47392 28244
rect 47408 28300 47472 28304
rect 47408 28244 47412 28300
rect 47412 28244 47468 28300
rect 47468 28244 47472 28300
rect 47408 28240 47472 28244
rect 47488 28300 47552 28304
rect 47488 28244 47492 28300
rect 47492 28244 47548 28300
rect 47548 28244 47552 28300
rect 47488 28240 47552 28244
rect 47568 28300 47632 28304
rect 47568 28244 47572 28300
rect 47572 28244 47628 28300
rect 47628 28244 47632 28300
rect 47568 28240 47632 28244
rect 47648 28300 47712 28304
rect 47648 28244 47652 28300
rect 47652 28244 47708 28300
rect 47708 28244 47712 28300
rect 47648 28240 47712 28244
rect 3372 26420 3436 26424
rect 3372 26364 3376 26420
rect 3376 26364 3432 26420
rect 3432 26364 3436 26420
rect 3372 26360 3436 26364
rect 3452 26420 3516 26424
rect 3452 26364 3456 26420
rect 3456 26364 3512 26420
rect 3512 26364 3516 26420
rect 3452 26360 3516 26364
rect 3532 26420 3596 26424
rect 3532 26364 3536 26420
rect 3536 26364 3592 26420
rect 3592 26364 3596 26420
rect 3532 26360 3596 26364
rect 3612 26420 3676 26424
rect 3612 26364 3616 26420
rect 3616 26364 3672 26420
rect 3672 26364 3676 26420
rect 3612 26360 3676 26364
rect 3692 26420 3756 26424
rect 3692 26364 3696 26420
rect 3696 26364 3752 26420
rect 3752 26364 3756 26420
rect 3692 26360 3756 26364
rect 3772 26420 3836 26424
rect 3772 26364 3776 26420
rect 3776 26364 3832 26420
rect 3832 26364 3836 26420
rect 3772 26360 3836 26364
rect 3852 26420 3916 26424
rect 3852 26364 3856 26420
rect 3856 26364 3912 26420
rect 3912 26364 3916 26420
rect 3852 26360 3916 26364
rect 3932 26420 3996 26424
rect 3932 26364 3936 26420
rect 3936 26364 3992 26420
rect 3992 26364 3996 26420
rect 3932 26360 3996 26364
rect 4012 26420 4076 26424
rect 4012 26364 4016 26420
rect 4016 26364 4072 26420
rect 4072 26364 4076 26420
rect 4012 26360 4076 26364
rect 4092 26420 4156 26424
rect 4092 26364 4096 26420
rect 4096 26364 4152 26420
rect 4152 26364 4156 26420
rect 4092 26360 4156 26364
rect 4172 26420 4236 26424
rect 4172 26364 4176 26420
rect 4176 26364 4232 26420
rect 4232 26364 4236 26420
rect 4172 26360 4236 26364
rect 4252 26420 4316 26424
rect 4252 26364 4256 26420
rect 4256 26364 4312 26420
rect 4312 26364 4316 26420
rect 4252 26360 4316 26364
rect 4332 26420 4396 26424
rect 4332 26364 4336 26420
rect 4336 26364 4392 26420
rect 4392 26364 4396 26420
rect 4332 26360 4396 26364
rect 4412 26420 4476 26424
rect 4412 26364 4416 26420
rect 4416 26364 4472 26420
rect 4472 26364 4476 26420
rect 4412 26360 4476 26364
rect 4492 26420 4556 26424
rect 4492 26364 4496 26420
rect 4496 26364 4552 26420
rect 4552 26364 4556 26420
rect 4492 26360 4556 26364
rect 4572 26420 4636 26424
rect 4572 26364 4576 26420
rect 4576 26364 4632 26420
rect 4632 26364 4636 26420
rect 4572 26360 4636 26364
rect 4652 26420 4716 26424
rect 4652 26364 4656 26420
rect 4656 26364 4712 26420
rect 4712 26364 4716 26420
rect 4652 26360 4716 26364
rect 4732 26420 4796 26424
rect 4732 26364 4736 26420
rect 4736 26364 4792 26420
rect 4792 26364 4796 26420
rect 4732 26360 4796 26364
rect 4812 26420 4876 26424
rect 4812 26364 4816 26420
rect 4816 26364 4872 26420
rect 4872 26364 4876 26420
rect 4812 26360 4876 26364
rect 4892 26420 4956 26424
rect 4892 26364 4896 26420
rect 4896 26364 4952 26420
rect 4952 26364 4956 26420
rect 4892 26360 4956 26364
rect 43680 26420 43744 26424
rect 43680 26364 43684 26420
rect 43684 26364 43740 26420
rect 43740 26364 43744 26420
rect 43680 26360 43744 26364
rect 43760 26420 43824 26424
rect 43760 26364 43764 26420
rect 43764 26364 43820 26420
rect 43820 26364 43824 26420
rect 43760 26360 43824 26364
rect 43840 26420 43904 26424
rect 43840 26364 43844 26420
rect 43844 26364 43900 26420
rect 43900 26364 43904 26420
rect 43840 26360 43904 26364
rect 43920 26420 43984 26424
rect 43920 26364 43924 26420
rect 43924 26364 43980 26420
rect 43980 26364 43984 26420
rect 43920 26360 43984 26364
rect 44000 26420 44064 26424
rect 44000 26364 44004 26420
rect 44004 26364 44060 26420
rect 44060 26364 44064 26420
rect 44000 26360 44064 26364
rect 44080 26420 44144 26424
rect 44080 26364 44084 26420
rect 44084 26364 44140 26420
rect 44140 26364 44144 26420
rect 44080 26360 44144 26364
rect 44160 26420 44224 26424
rect 44160 26364 44164 26420
rect 44164 26364 44220 26420
rect 44220 26364 44224 26420
rect 44160 26360 44224 26364
rect 44240 26420 44304 26424
rect 44240 26364 44244 26420
rect 44244 26364 44300 26420
rect 44300 26364 44304 26420
rect 44240 26360 44304 26364
rect 44320 26420 44384 26424
rect 44320 26364 44324 26420
rect 44324 26364 44380 26420
rect 44380 26364 44384 26420
rect 44320 26360 44384 26364
rect 44400 26420 44464 26424
rect 44400 26364 44404 26420
rect 44404 26364 44460 26420
rect 44460 26364 44464 26420
rect 44400 26360 44464 26364
rect 44480 26420 44544 26424
rect 44480 26364 44484 26420
rect 44484 26364 44540 26420
rect 44540 26364 44544 26420
rect 44480 26360 44544 26364
rect 44560 26420 44624 26424
rect 44560 26364 44564 26420
rect 44564 26364 44620 26420
rect 44620 26364 44624 26420
rect 44560 26360 44624 26364
rect 44640 26420 44704 26424
rect 44640 26364 44644 26420
rect 44644 26364 44700 26420
rect 44700 26364 44704 26420
rect 44640 26360 44704 26364
rect 44720 26420 44784 26424
rect 44720 26364 44724 26420
rect 44724 26364 44780 26420
rect 44780 26364 44784 26420
rect 44720 26360 44784 26364
rect 44800 26420 44864 26424
rect 44800 26364 44804 26420
rect 44804 26364 44860 26420
rect 44860 26364 44864 26420
rect 44800 26360 44864 26364
rect 44880 26420 44944 26424
rect 44880 26364 44884 26420
rect 44884 26364 44940 26420
rect 44940 26364 44944 26420
rect 44880 26360 44944 26364
rect 44960 26420 45024 26424
rect 44960 26364 44964 26420
rect 44964 26364 45020 26420
rect 45020 26364 45024 26420
rect 44960 26360 45024 26364
rect 45040 26420 45104 26424
rect 45040 26364 45044 26420
rect 45044 26364 45100 26420
rect 45100 26364 45104 26420
rect 45040 26360 45104 26364
rect 45120 26420 45184 26424
rect 45120 26364 45124 26420
rect 45124 26364 45180 26420
rect 45180 26364 45184 26420
rect 45120 26360 45184 26364
rect 45200 26420 45264 26424
rect 45200 26364 45204 26420
rect 45204 26364 45260 26420
rect 45260 26364 45264 26420
rect 45200 26360 45264 26364
rect 16038 26070 16102 26134
rect 16757 26070 16821 26134
rect 17476 26070 17540 26134
rect 18195 26070 18259 26134
rect 18914 26070 18978 26134
rect 19633 26070 19697 26134
rect 20352 26070 20416 26134
rect 21071 26070 21135 26134
rect 21790 26070 21854 26134
rect 22509 26070 22573 26134
rect 16038 25990 16102 26054
rect 16757 25990 16821 26054
rect 17476 25990 17540 26054
rect 18195 25990 18259 26054
rect 18914 25990 18978 26054
rect 19633 25990 19697 26054
rect 20352 25990 20416 26054
rect 21071 25990 21135 26054
rect 21790 25990 21854 26054
rect 22509 25990 22573 26054
rect 16038 25910 16102 25974
rect 16757 25910 16821 25974
rect 17476 25910 17540 25974
rect 18195 25910 18259 25974
rect 18914 25910 18978 25974
rect 19633 25910 19697 25974
rect 20352 25910 20416 25974
rect 21071 25910 21135 25974
rect 21790 25910 21854 25974
rect 22509 25910 22573 25974
rect 16038 25830 16102 25894
rect 16757 25830 16821 25894
rect 17476 25830 17540 25894
rect 18195 25830 18259 25894
rect 18914 25830 18978 25894
rect 19633 25830 19697 25894
rect 20352 25830 20416 25894
rect 21071 25830 21135 25894
rect 21790 25830 21854 25894
rect 22509 25830 22573 25894
rect 16038 25750 16102 25814
rect 16757 25750 16821 25814
rect 17476 25750 17540 25814
rect 18195 25750 18259 25814
rect 18914 25750 18978 25814
rect 19633 25750 19697 25814
rect 20352 25750 20416 25814
rect 21071 25750 21135 25814
rect 21790 25750 21854 25814
rect 22509 25750 22573 25814
rect 16038 25670 16102 25734
rect 16757 25670 16821 25734
rect 17476 25670 17540 25734
rect 18195 25670 18259 25734
rect 18914 25670 18978 25734
rect 19633 25670 19697 25734
rect 20352 25670 20416 25734
rect 21071 25670 21135 25734
rect 21790 25670 21854 25734
rect 22509 25670 22573 25734
rect 16038 25590 16102 25654
rect 16757 25590 16821 25654
rect 17476 25590 17540 25654
rect 18195 25590 18259 25654
rect 18914 25590 18978 25654
rect 19633 25590 19697 25654
rect 20352 25590 20416 25654
rect 21071 25590 21135 25654
rect 21790 25590 21854 25654
rect 22509 25590 22573 25654
rect 16038 25370 16102 25434
rect 16757 25370 16821 25434
rect 17476 25370 17540 25434
rect 18195 25370 18259 25434
rect 18914 25370 18978 25434
rect 19633 25370 19697 25434
rect 20352 25370 20416 25434
rect 21071 25370 21135 25434
rect 21790 25370 21854 25434
rect 22509 25370 22573 25434
rect 16038 25290 16102 25354
rect 16757 25290 16821 25354
rect 17476 25290 17540 25354
rect 18195 25290 18259 25354
rect 18914 25290 18978 25354
rect 19633 25290 19697 25354
rect 20352 25290 20416 25354
rect 21071 25290 21135 25354
rect 21790 25290 21854 25354
rect 22509 25290 22573 25354
rect 16038 25210 16102 25274
rect 16757 25210 16821 25274
rect 17476 25210 17540 25274
rect 18195 25210 18259 25274
rect 18914 25210 18978 25274
rect 19633 25210 19697 25274
rect 20352 25210 20416 25274
rect 21071 25210 21135 25274
rect 21790 25210 21854 25274
rect 22509 25210 22573 25274
rect 16038 25130 16102 25194
rect 16757 25130 16821 25194
rect 17476 25130 17540 25194
rect 18195 25130 18259 25194
rect 18914 25130 18978 25194
rect 19633 25130 19697 25194
rect 20352 25130 20416 25194
rect 21071 25130 21135 25194
rect 21790 25130 21854 25194
rect 22509 25130 22573 25194
rect 16038 25050 16102 25114
rect 16757 25050 16821 25114
rect 17476 25050 17540 25114
rect 18195 25050 18259 25114
rect 18914 25050 18978 25114
rect 19633 25050 19697 25114
rect 20352 25050 20416 25114
rect 21071 25050 21135 25114
rect 21790 25050 21854 25114
rect 22509 25050 22573 25114
rect 16038 24970 16102 25034
rect 16757 24970 16821 25034
rect 17476 24970 17540 25034
rect 18195 24970 18259 25034
rect 18914 24970 18978 25034
rect 19633 24970 19697 25034
rect 20352 24970 20416 25034
rect 21071 24970 21135 25034
rect 21790 24970 21854 25034
rect 22509 24970 22573 25034
rect 22784 24990 22848 25054
rect 16038 24890 16102 24954
rect 16757 24890 16821 24954
rect 17476 24890 17540 24954
rect 18195 24890 18259 24954
rect 18914 24890 18978 24954
rect 19633 24890 19697 24954
rect 20352 24890 20416 24954
rect 21071 24890 21135 24954
rect 21790 24890 21854 24954
rect 22509 24890 22573 24954
rect 15452 24730 15516 24734
rect 15532 24730 15596 24734
rect 15452 24674 15496 24730
rect 15496 24674 15516 24730
rect 15532 24674 15552 24730
rect 15552 24674 15596 24730
rect 15452 24670 15516 24674
rect 15532 24670 15596 24674
rect 924 24540 988 24544
rect 924 24484 928 24540
rect 928 24484 984 24540
rect 984 24484 988 24540
rect 924 24480 988 24484
rect 1004 24540 1068 24544
rect 1004 24484 1008 24540
rect 1008 24484 1064 24540
rect 1064 24484 1068 24540
rect 1004 24480 1068 24484
rect 1084 24540 1148 24544
rect 1084 24484 1088 24540
rect 1088 24484 1144 24540
rect 1144 24484 1148 24540
rect 1084 24480 1148 24484
rect 1164 24540 1228 24544
rect 1164 24484 1168 24540
rect 1168 24484 1224 24540
rect 1224 24484 1228 24540
rect 1164 24480 1228 24484
rect 1244 24540 1308 24544
rect 1244 24484 1248 24540
rect 1248 24484 1304 24540
rect 1304 24484 1308 24540
rect 1244 24480 1308 24484
rect 1324 24540 1388 24544
rect 1324 24484 1328 24540
rect 1328 24484 1384 24540
rect 1384 24484 1388 24540
rect 1324 24480 1388 24484
rect 1404 24540 1468 24544
rect 1404 24484 1408 24540
rect 1408 24484 1464 24540
rect 1464 24484 1468 24540
rect 1404 24480 1468 24484
rect 1484 24540 1548 24544
rect 1484 24484 1488 24540
rect 1488 24484 1544 24540
rect 1544 24484 1548 24540
rect 1484 24480 1548 24484
rect 1564 24540 1628 24544
rect 1564 24484 1568 24540
rect 1568 24484 1624 24540
rect 1624 24484 1628 24540
rect 1564 24480 1628 24484
rect 1644 24540 1708 24544
rect 1644 24484 1648 24540
rect 1648 24484 1704 24540
rect 1704 24484 1708 24540
rect 1644 24480 1708 24484
rect 1724 24540 1788 24544
rect 1724 24484 1728 24540
rect 1728 24484 1784 24540
rect 1784 24484 1788 24540
rect 1724 24480 1788 24484
rect 1804 24540 1868 24544
rect 1804 24484 1808 24540
rect 1808 24484 1864 24540
rect 1864 24484 1868 24540
rect 1804 24480 1868 24484
rect 1884 24540 1948 24544
rect 1884 24484 1888 24540
rect 1888 24484 1944 24540
rect 1944 24484 1948 24540
rect 1884 24480 1948 24484
rect 1964 24540 2028 24544
rect 1964 24484 1968 24540
rect 1968 24484 2024 24540
rect 2024 24484 2028 24540
rect 1964 24480 2028 24484
rect 2044 24540 2108 24544
rect 2044 24484 2048 24540
rect 2048 24484 2104 24540
rect 2104 24484 2108 24540
rect 2044 24480 2108 24484
rect 2124 24540 2188 24544
rect 2124 24484 2128 24540
rect 2128 24484 2184 24540
rect 2184 24484 2188 24540
rect 2124 24480 2188 24484
rect 2204 24540 2268 24544
rect 2204 24484 2208 24540
rect 2208 24484 2264 24540
rect 2264 24484 2268 24540
rect 2204 24480 2268 24484
rect 2284 24540 2348 24544
rect 2284 24484 2288 24540
rect 2288 24484 2344 24540
rect 2344 24484 2348 24540
rect 2284 24480 2348 24484
rect 2364 24540 2428 24544
rect 2364 24484 2368 24540
rect 2368 24484 2424 24540
rect 2424 24484 2428 24540
rect 2364 24480 2428 24484
rect 2444 24540 2508 24544
rect 2444 24484 2448 24540
rect 2448 24484 2504 24540
rect 2504 24484 2508 24540
rect 2444 24480 2508 24484
rect 15470 24562 15534 24566
rect 15470 24506 15474 24562
rect 15474 24506 15530 24562
rect 15530 24506 15534 24562
rect 15470 24502 15534 24506
rect 46128 24540 46192 24544
rect 46128 24484 46132 24540
rect 46132 24484 46188 24540
rect 46188 24484 46192 24540
rect 46128 24480 46192 24484
rect 46208 24540 46272 24544
rect 46208 24484 46212 24540
rect 46212 24484 46268 24540
rect 46268 24484 46272 24540
rect 46208 24480 46272 24484
rect 46288 24540 46352 24544
rect 46288 24484 46292 24540
rect 46292 24484 46348 24540
rect 46348 24484 46352 24540
rect 46288 24480 46352 24484
rect 46368 24540 46432 24544
rect 46368 24484 46372 24540
rect 46372 24484 46428 24540
rect 46428 24484 46432 24540
rect 46368 24480 46432 24484
rect 46448 24540 46512 24544
rect 46448 24484 46452 24540
rect 46452 24484 46508 24540
rect 46508 24484 46512 24540
rect 46448 24480 46512 24484
rect 46528 24540 46592 24544
rect 46528 24484 46532 24540
rect 46532 24484 46588 24540
rect 46588 24484 46592 24540
rect 46528 24480 46592 24484
rect 46608 24540 46672 24544
rect 46608 24484 46612 24540
rect 46612 24484 46668 24540
rect 46668 24484 46672 24540
rect 46608 24480 46672 24484
rect 46688 24540 46752 24544
rect 46688 24484 46692 24540
rect 46692 24484 46748 24540
rect 46748 24484 46752 24540
rect 46688 24480 46752 24484
rect 46768 24540 46832 24544
rect 46768 24484 46772 24540
rect 46772 24484 46828 24540
rect 46828 24484 46832 24540
rect 46768 24480 46832 24484
rect 46848 24540 46912 24544
rect 46848 24484 46852 24540
rect 46852 24484 46908 24540
rect 46908 24484 46912 24540
rect 46848 24480 46912 24484
rect 46928 24540 46992 24544
rect 46928 24484 46932 24540
rect 46932 24484 46988 24540
rect 46988 24484 46992 24540
rect 46928 24480 46992 24484
rect 47008 24540 47072 24544
rect 47008 24484 47012 24540
rect 47012 24484 47068 24540
rect 47068 24484 47072 24540
rect 47008 24480 47072 24484
rect 47088 24540 47152 24544
rect 47088 24484 47092 24540
rect 47092 24484 47148 24540
rect 47148 24484 47152 24540
rect 47088 24480 47152 24484
rect 47168 24540 47232 24544
rect 47168 24484 47172 24540
rect 47172 24484 47228 24540
rect 47228 24484 47232 24540
rect 47168 24480 47232 24484
rect 47248 24540 47312 24544
rect 47248 24484 47252 24540
rect 47252 24484 47308 24540
rect 47308 24484 47312 24540
rect 47248 24480 47312 24484
rect 47328 24540 47392 24544
rect 47328 24484 47332 24540
rect 47332 24484 47388 24540
rect 47388 24484 47392 24540
rect 47328 24480 47392 24484
rect 47408 24540 47472 24544
rect 47408 24484 47412 24540
rect 47412 24484 47468 24540
rect 47468 24484 47472 24540
rect 47408 24480 47472 24484
rect 47488 24540 47552 24544
rect 47488 24484 47492 24540
rect 47492 24484 47548 24540
rect 47548 24484 47552 24540
rect 47488 24480 47552 24484
rect 47568 24540 47632 24544
rect 47568 24484 47572 24540
rect 47572 24484 47628 24540
rect 47628 24484 47632 24540
rect 47568 24480 47632 24484
rect 47648 24540 47712 24544
rect 47648 24484 47652 24540
rect 47652 24484 47708 24540
rect 47708 24484 47712 24540
rect 47648 24480 47712 24484
rect 3372 22660 3436 22664
rect 3372 22604 3376 22660
rect 3376 22604 3432 22660
rect 3432 22604 3436 22660
rect 3372 22600 3436 22604
rect 3452 22660 3516 22664
rect 3452 22604 3456 22660
rect 3456 22604 3512 22660
rect 3512 22604 3516 22660
rect 3452 22600 3516 22604
rect 3532 22660 3596 22664
rect 3532 22604 3536 22660
rect 3536 22604 3592 22660
rect 3592 22604 3596 22660
rect 3532 22600 3596 22604
rect 3612 22660 3676 22664
rect 3612 22604 3616 22660
rect 3616 22604 3672 22660
rect 3672 22604 3676 22660
rect 3612 22600 3676 22604
rect 3692 22660 3756 22664
rect 3692 22604 3696 22660
rect 3696 22604 3752 22660
rect 3752 22604 3756 22660
rect 3692 22600 3756 22604
rect 3772 22660 3836 22664
rect 3772 22604 3776 22660
rect 3776 22604 3832 22660
rect 3832 22604 3836 22660
rect 3772 22600 3836 22604
rect 3852 22660 3916 22664
rect 3852 22604 3856 22660
rect 3856 22604 3912 22660
rect 3912 22604 3916 22660
rect 3852 22600 3916 22604
rect 3932 22660 3996 22664
rect 3932 22604 3936 22660
rect 3936 22604 3992 22660
rect 3992 22604 3996 22660
rect 3932 22600 3996 22604
rect 4012 22660 4076 22664
rect 4012 22604 4016 22660
rect 4016 22604 4072 22660
rect 4072 22604 4076 22660
rect 4012 22600 4076 22604
rect 4092 22660 4156 22664
rect 4092 22604 4096 22660
rect 4096 22604 4152 22660
rect 4152 22604 4156 22660
rect 4092 22600 4156 22604
rect 4172 22660 4236 22664
rect 4172 22604 4176 22660
rect 4176 22604 4232 22660
rect 4232 22604 4236 22660
rect 4172 22600 4236 22604
rect 4252 22660 4316 22664
rect 4252 22604 4256 22660
rect 4256 22604 4312 22660
rect 4312 22604 4316 22660
rect 4252 22600 4316 22604
rect 4332 22660 4396 22664
rect 4332 22604 4336 22660
rect 4336 22604 4392 22660
rect 4392 22604 4396 22660
rect 4332 22600 4396 22604
rect 4412 22660 4476 22664
rect 4412 22604 4416 22660
rect 4416 22604 4472 22660
rect 4472 22604 4476 22660
rect 4412 22600 4476 22604
rect 4492 22660 4556 22664
rect 4492 22604 4496 22660
rect 4496 22604 4552 22660
rect 4552 22604 4556 22660
rect 4492 22600 4556 22604
rect 4572 22660 4636 22664
rect 4572 22604 4576 22660
rect 4576 22604 4632 22660
rect 4632 22604 4636 22660
rect 4572 22600 4636 22604
rect 4652 22660 4716 22664
rect 4652 22604 4656 22660
rect 4656 22604 4712 22660
rect 4712 22604 4716 22660
rect 4652 22600 4716 22604
rect 4732 22660 4796 22664
rect 4732 22604 4736 22660
rect 4736 22604 4792 22660
rect 4792 22604 4796 22660
rect 4732 22600 4796 22604
rect 4812 22660 4876 22664
rect 4812 22604 4816 22660
rect 4816 22604 4872 22660
rect 4872 22604 4876 22660
rect 4812 22600 4876 22604
rect 4892 22660 4956 22664
rect 4892 22604 4896 22660
rect 4896 22604 4952 22660
rect 4952 22604 4956 22660
rect 4892 22600 4956 22604
rect 14228 22550 14292 22614
rect 43680 22660 43744 22664
rect 43680 22604 43684 22660
rect 43684 22604 43740 22660
rect 43740 22604 43744 22660
rect 43680 22600 43744 22604
rect 43760 22660 43824 22664
rect 43760 22604 43764 22660
rect 43764 22604 43820 22660
rect 43820 22604 43824 22660
rect 43760 22600 43824 22604
rect 43840 22660 43904 22664
rect 43840 22604 43844 22660
rect 43844 22604 43900 22660
rect 43900 22604 43904 22660
rect 43840 22600 43904 22604
rect 43920 22660 43984 22664
rect 43920 22604 43924 22660
rect 43924 22604 43980 22660
rect 43980 22604 43984 22660
rect 43920 22600 43984 22604
rect 44000 22660 44064 22664
rect 44000 22604 44004 22660
rect 44004 22604 44060 22660
rect 44060 22604 44064 22660
rect 44000 22600 44064 22604
rect 44080 22660 44144 22664
rect 44080 22604 44084 22660
rect 44084 22604 44140 22660
rect 44140 22604 44144 22660
rect 44080 22600 44144 22604
rect 44160 22660 44224 22664
rect 44160 22604 44164 22660
rect 44164 22604 44220 22660
rect 44220 22604 44224 22660
rect 44160 22600 44224 22604
rect 44240 22660 44304 22664
rect 44240 22604 44244 22660
rect 44244 22604 44300 22660
rect 44300 22604 44304 22660
rect 44240 22600 44304 22604
rect 44320 22660 44384 22664
rect 44320 22604 44324 22660
rect 44324 22604 44380 22660
rect 44380 22604 44384 22660
rect 44320 22600 44384 22604
rect 44400 22660 44464 22664
rect 44400 22604 44404 22660
rect 44404 22604 44460 22660
rect 44460 22604 44464 22660
rect 44400 22600 44464 22604
rect 44480 22660 44544 22664
rect 44480 22604 44484 22660
rect 44484 22604 44540 22660
rect 44540 22604 44544 22660
rect 44480 22600 44544 22604
rect 44560 22660 44624 22664
rect 44560 22604 44564 22660
rect 44564 22604 44620 22660
rect 44620 22604 44624 22660
rect 44560 22600 44624 22604
rect 44640 22660 44704 22664
rect 44640 22604 44644 22660
rect 44644 22604 44700 22660
rect 44700 22604 44704 22660
rect 44640 22600 44704 22604
rect 44720 22660 44784 22664
rect 44720 22604 44724 22660
rect 44724 22604 44780 22660
rect 44780 22604 44784 22660
rect 44720 22600 44784 22604
rect 44800 22660 44864 22664
rect 44800 22604 44804 22660
rect 44804 22604 44860 22660
rect 44860 22604 44864 22660
rect 44800 22600 44864 22604
rect 44880 22660 44944 22664
rect 44880 22604 44884 22660
rect 44884 22604 44940 22660
rect 44940 22604 44944 22660
rect 44880 22600 44944 22604
rect 44960 22660 45024 22664
rect 44960 22604 44964 22660
rect 44964 22604 45020 22660
rect 45020 22604 45024 22660
rect 44960 22600 45024 22604
rect 45040 22660 45104 22664
rect 45040 22604 45044 22660
rect 45044 22604 45100 22660
rect 45100 22604 45104 22660
rect 45040 22600 45104 22604
rect 45120 22660 45184 22664
rect 45120 22604 45124 22660
rect 45124 22604 45180 22660
rect 45180 22604 45184 22660
rect 45120 22600 45184 22604
rect 45200 22660 45264 22664
rect 45200 22604 45204 22660
rect 45204 22604 45260 22660
rect 45260 22604 45264 22660
rect 45200 22600 45264 22604
rect 14176 22310 14240 22374
rect 14895 22310 14959 22374
rect 15614 22310 15678 22374
rect 16333 22310 16397 22374
rect 17052 22310 17116 22374
rect 17771 22310 17835 22374
rect 18490 22310 18554 22374
rect 19209 22310 19273 22374
rect 19928 22310 19992 22374
rect 20647 22310 20711 22374
rect 14176 22230 14240 22294
rect 14895 22230 14959 22294
rect 15614 22230 15678 22294
rect 16333 22230 16397 22294
rect 17052 22230 17116 22294
rect 17771 22230 17835 22294
rect 18490 22230 18554 22294
rect 19209 22230 19273 22294
rect 19928 22230 19992 22294
rect 20647 22230 20711 22294
rect 14176 22150 14240 22214
rect 14895 22150 14959 22214
rect 15614 22150 15678 22214
rect 16333 22150 16397 22214
rect 17052 22150 17116 22214
rect 17771 22150 17835 22214
rect 18490 22150 18554 22214
rect 19209 22150 19273 22214
rect 19928 22150 19992 22214
rect 20647 22150 20711 22214
rect 14176 22070 14240 22134
rect 14895 22070 14959 22134
rect 15614 22070 15678 22134
rect 16333 22070 16397 22134
rect 17052 22070 17116 22134
rect 17771 22070 17835 22134
rect 18490 22070 18554 22134
rect 19209 22070 19273 22134
rect 19928 22070 19992 22134
rect 20647 22070 20711 22134
rect 14176 21990 14240 22054
rect 14895 21990 14959 22054
rect 15614 21990 15678 22054
rect 16333 21990 16397 22054
rect 17052 21990 17116 22054
rect 17771 21990 17835 22054
rect 18490 21990 18554 22054
rect 19209 21990 19273 22054
rect 19928 21990 19992 22054
rect 20647 21990 20711 22054
rect 14176 21910 14240 21974
rect 14895 21910 14959 21974
rect 15614 21910 15678 21974
rect 16333 21910 16397 21974
rect 17052 21910 17116 21974
rect 17771 21910 17835 21974
rect 18490 21910 18554 21974
rect 19209 21910 19273 21974
rect 19928 21910 19992 21974
rect 20647 21910 20711 21974
rect 14176 21830 14240 21894
rect 14895 21830 14959 21894
rect 15614 21830 15678 21894
rect 16333 21830 16397 21894
rect 17052 21830 17116 21894
rect 17771 21830 17835 21894
rect 18490 21830 18554 21894
rect 19209 21830 19273 21894
rect 19928 21830 19992 21894
rect 20647 21830 20711 21894
rect 14176 21610 14240 21674
rect 14895 21610 14959 21674
rect 15614 21610 15678 21674
rect 16333 21610 16397 21674
rect 17052 21610 17116 21674
rect 17771 21610 17835 21674
rect 18490 21610 18554 21674
rect 19209 21610 19273 21674
rect 19928 21610 19992 21674
rect 20647 21610 20711 21674
rect 14176 21530 14240 21594
rect 14895 21530 14959 21594
rect 15614 21530 15678 21594
rect 16333 21530 16397 21594
rect 17052 21530 17116 21594
rect 17771 21530 17835 21594
rect 18490 21530 18554 21594
rect 19209 21530 19273 21594
rect 19928 21530 19992 21594
rect 20647 21530 20711 21594
rect 20852 21634 20916 21638
rect 20852 21578 20902 21634
rect 20902 21578 20916 21634
rect 20852 21574 20916 21578
rect 14176 21450 14240 21514
rect 14895 21450 14959 21514
rect 15614 21450 15678 21514
rect 16333 21450 16397 21514
rect 17052 21450 17116 21514
rect 17771 21450 17835 21514
rect 18490 21450 18554 21514
rect 19209 21450 19273 21514
rect 19928 21450 19992 21514
rect 20647 21450 20711 21514
rect 14176 21370 14240 21434
rect 14895 21370 14959 21434
rect 15614 21370 15678 21434
rect 16333 21370 16397 21434
rect 17052 21370 17116 21434
rect 17771 21370 17835 21434
rect 18490 21370 18554 21434
rect 19209 21370 19273 21434
rect 19928 21370 19992 21434
rect 20647 21370 20711 21434
rect 14176 21290 14240 21354
rect 14895 21290 14959 21354
rect 15614 21290 15678 21354
rect 16333 21290 16397 21354
rect 17052 21290 17116 21354
rect 17771 21290 17835 21354
rect 18490 21290 18554 21354
rect 19209 21290 19273 21354
rect 19928 21290 19992 21354
rect 20647 21290 20711 21354
rect 14176 21210 14240 21274
rect 14895 21210 14959 21274
rect 15614 21210 15678 21274
rect 16333 21210 16397 21274
rect 17052 21210 17116 21274
rect 17771 21210 17835 21274
rect 18490 21210 18554 21274
rect 19209 21210 19273 21274
rect 19928 21210 19992 21274
rect 20647 21210 20711 21274
rect 14176 21130 14240 21194
rect 14895 21130 14959 21194
rect 15614 21130 15678 21194
rect 16333 21130 16397 21194
rect 17052 21130 17116 21194
rect 17771 21130 17835 21194
rect 18490 21130 18554 21194
rect 19209 21130 19273 21194
rect 19928 21130 19992 21194
rect 20647 21130 20711 21194
rect 13590 20970 13654 20974
rect 13670 20970 13734 20974
rect 13590 20914 13634 20970
rect 13634 20914 13654 20970
rect 13670 20914 13690 20970
rect 13690 20914 13734 20970
rect 13590 20910 13654 20914
rect 13670 20910 13734 20914
rect 14090 20902 14154 20906
rect 14090 20846 14094 20902
rect 14094 20846 14150 20902
rect 14150 20846 14154 20902
rect 14090 20842 14154 20846
rect 924 20780 988 20784
rect 924 20724 928 20780
rect 928 20724 984 20780
rect 984 20724 988 20780
rect 924 20720 988 20724
rect 1004 20780 1068 20784
rect 1004 20724 1008 20780
rect 1008 20724 1064 20780
rect 1064 20724 1068 20780
rect 1004 20720 1068 20724
rect 1084 20780 1148 20784
rect 1084 20724 1088 20780
rect 1088 20724 1144 20780
rect 1144 20724 1148 20780
rect 1084 20720 1148 20724
rect 1164 20780 1228 20784
rect 1164 20724 1168 20780
rect 1168 20724 1224 20780
rect 1224 20724 1228 20780
rect 1164 20720 1228 20724
rect 1244 20780 1308 20784
rect 1244 20724 1248 20780
rect 1248 20724 1304 20780
rect 1304 20724 1308 20780
rect 1244 20720 1308 20724
rect 1324 20780 1388 20784
rect 1324 20724 1328 20780
rect 1328 20724 1384 20780
rect 1384 20724 1388 20780
rect 1324 20720 1388 20724
rect 1404 20780 1468 20784
rect 1404 20724 1408 20780
rect 1408 20724 1464 20780
rect 1464 20724 1468 20780
rect 1404 20720 1468 20724
rect 1484 20780 1548 20784
rect 1484 20724 1488 20780
rect 1488 20724 1544 20780
rect 1544 20724 1548 20780
rect 1484 20720 1548 20724
rect 1564 20780 1628 20784
rect 1564 20724 1568 20780
rect 1568 20724 1624 20780
rect 1624 20724 1628 20780
rect 1564 20720 1628 20724
rect 1644 20780 1708 20784
rect 1644 20724 1648 20780
rect 1648 20724 1704 20780
rect 1704 20724 1708 20780
rect 1644 20720 1708 20724
rect 1724 20780 1788 20784
rect 1724 20724 1728 20780
rect 1728 20724 1784 20780
rect 1784 20724 1788 20780
rect 1724 20720 1788 20724
rect 1804 20780 1868 20784
rect 1804 20724 1808 20780
rect 1808 20724 1864 20780
rect 1864 20724 1868 20780
rect 1804 20720 1868 20724
rect 1884 20780 1948 20784
rect 1884 20724 1888 20780
rect 1888 20724 1944 20780
rect 1944 20724 1948 20780
rect 1884 20720 1948 20724
rect 1964 20780 2028 20784
rect 1964 20724 1968 20780
rect 1968 20724 2024 20780
rect 2024 20724 2028 20780
rect 1964 20720 2028 20724
rect 2044 20780 2108 20784
rect 2044 20724 2048 20780
rect 2048 20724 2104 20780
rect 2104 20724 2108 20780
rect 2044 20720 2108 20724
rect 2124 20780 2188 20784
rect 2124 20724 2128 20780
rect 2128 20724 2184 20780
rect 2184 20724 2188 20780
rect 2124 20720 2188 20724
rect 2204 20780 2268 20784
rect 2204 20724 2208 20780
rect 2208 20724 2264 20780
rect 2264 20724 2268 20780
rect 2204 20720 2268 20724
rect 2284 20780 2348 20784
rect 2284 20724 2288 20780
rect 2288 20724 2344 20780
rect 2344 20724 2348 20780
rect 2284 20720 2348 20724
rect 2364 20780 2428 20784
rect 2364 20724 2368 20780
rect 2368 20724 2424 20780
rect 2424 20724 2428 20780
rect 2364 20720 2428 20724
rect 2444 20780 2508 20784
rect 2444 20724 2448 20780
rect 2448 20724 2504 20780
rect 2504 20724 2508 20780
rect 2444 20720 2508 20724
rect 46128 20780 46192 20784
rect 46128 20724 46132 20780
rect 46132 20724 46188 20780
rect 46188 20724 46192 20780
rect 46128 20720 46192 20724
rect 46208 20780 46272 20784
rect 46208 20724 46212 20780
rect 46212 20724 46268 20780
rect 46268 20724 46272 20780
rect 46208 20720 46272 20724
rect 46288 20780 46352 20784
rect 46288 20724 46292 20780
rect 46292 20724 46348 20780
rect 46348 20724 46352 20780
rect 46288 20720 46352 20724
rect 46368 20780 46432 20784
rect 46368 20724 46372 20780
rect 46372 20724 46428 20780
rect 46428 20724 46432 20780
rect 46368 20720 46432 20724
rect 46448 20780 46512 20784
rect 46448 20724 46452 20780
rect 46452 20724 46508 20780
rect 46508 20724 46512 20780
rect 46448 20720 46512 20724
rect 46528 20780 46592 20784
rect 46528 20724 46532 20780
rect 46532 20724 46588 20780
rect 46588 20724 46592 20780
rect 46528 20720 46592 20724
rect 46608 20780 46672 20784
rect 46608 20724 46612 20780
rect 46612 20724 46668 20780
rect 46668 20724 46672 20780
rect 46608 20720 46672 20724
rect 46688 20780 46752 20784
rect 46688 20724 46692 20780
rect 46692 20724 46748 20780
rect 46748 20724 46752 20780
rect 46688 20720 46752 20724
rect 46768 20780 46832 20784
rect 46768 20724 46772 20780
rect 46772 20724 46828 20780
rect 46828 20724 46832 20780
rect 46768 20720 46832 20724
rect 46848 20780 46912 20784
rect 46848 20724 46852 20780
rect 46852 20724 46908 20780
rect 46908 20724 46912 20780
rect 46848 20720 46912 20724
rect 46928 20780 46992 20784
rect 46928 20724 46932 20780
rect 46932 20724 46988 20780
rect 46988 20724 46992 20780
rect 46928 20720 46992 20724
rect 47008 20780 47072 20784
rect 47008 20724 47012 20780
rect 47012 20724 47068 20780
rect 47068 20724 47072 20780
rect 47008 20720 47072 20724
rect 47088 20780 47152 20784
rect 47088 20724 47092 20780
rect 47092 20724 47148 20780
rect 47148 20724 47152 20780
rect 47088 20720 47152 20724
rect 47168 20780 47232 20784
rect 47168 20724 47172 20780
rect 47172 20724 47228 20780
rect 47228 20724 47232 20780
rect 47168 20720 47232 20724
rect 47248 20780 47312 20784
rect 47248 20724 47252 20780
rect 47252 20724 47308 20780
rect 47308 20724 47312 20780
rect 47248 20720 47312 20724
rect 47328 20780 47392 20784
rect 47328 20724 47332 20780
rect 47332 20724 47388 20780
rect 47388 20724 47392 20780
rect 47328 20720 47392 20724
rect 47408 20780 47472 20784
rect 47408 20724 47412 20780
rect 47412 20724 47468 20780
rect 47468 20724 47472 20780
rect 47408 20720 47472 20724
rect 47488 20780 47552 20784
rect 47488 20724 47492 20780
rect 47492 20724 47548 20780
rect 47548 20724 47552 20780
rect 47488 20720 47552 20724
rect 47568 20780 47632 20784
rect 47568 20724 47572 20780
rect 47572 20724 47628 20780
rect 47628 20724 47632 20780
rect 47568 20720 47632 20724
rect 47648 20780 47712 20784
rect 47648 20724 47652 20780
rect 47652 20724 47708 20780
rect 47708 20724 47712 20780
rect 47648 20720 47712 20724
rect 3372 18900 3436 18904
rect 3372 18844 3376 18900
rect 3376 18844 3432 18900
rect 3432 18844 3436 18900
rect 3372 18840 3436 18844
rect 3452 18900 3516 18904
rect 3452 18844 3456 18900
rect 3456 18844 3512 18900
rect 3512 18844 3516 18900
rect 3452 18840 3516 18844
rect 3532 18900 3596 18904
rect 3532 18844 3536 18900
rect 3536 18844 3592 18900
rect 3592 18844 3596 18900
rect 3532 18840 3596 18844
rect 3612 18900 3676 18904
rect 3612 18844 3616 18900
rect 3616 18844 3672 18900
rect 3672 18844 3676 18900
rect 3612 18840 3676 18844
rect 3692 18900 3756 18904
rect 3692 18844 3696 18900
rect 3696 18844 3752 18900
rect 3752 18844 3756 18900
rect 3692 18840 3756 18844
rect 3772 18900 3836 18904
rect 3772 18844 3776 18900
rect 3776 18844 3832 18900
rect 3832 18844 3836 18900
rect 3772 18840 3836 18844
rect 3852 18900 3916 18904
rect 3852 18844 3856 18900
rect 3856 18844 3912 18900
rect 3912 18844 3916 18900
rect 3852 18840 3916 18844
rect 3932 18900 3996 18904
rect 3932 18844 3936 18900
rect 3936 18844 3992 18900
rect 3992 18844 3996 18900
rect 3932 18840 3996 18844
rect 4012 18900 4076 18904
rect 4012 18844 4016 18900
rect 4016 18844 4072 18900
rect 4072 18844 4076 18900
rect 4012 18840 4076 18844
rect 4092 18900 4156 18904
rect 4092 18844 4096 18900
rect 4096 18844 4152 18900
rect 4152 18844 4156 18900
rect 4092 18840 4156 18844
rect 4172 18900 4236 18904
rect 4172 18844 4176 18900
rect 4176 18844 4232 18900
rect 4232 18844 4236 18900
rect 4172 18840 4236 18844
rect 4252 18900 4316 18904
rect 4252 18844 4256 18900
rect 4256 18844 4312 18900
rect 4312 18844 4316 18900
rect 4252 18840 4316 18844
rect 4332 18900 4396 18904
rect 4332 18844 4336 18900
rect 4336 18844 4392 18900
rect 4392 18844 4396 18900
rect 4332 18840 4396 18844
rect 4412 18900 4476 18904
rect 4412 18844 4416 18900
rect 4416 18844 4472 18900
rect 4472 18844 4476 18900
rect 4412 18840 4476 18844
rect 4492 18900 4556 18904
rect 4492 18844 4496 18900
rect 4496 18844 4552 18900
rect 4552 18844 4556 18900
rect 4492 18840 4556 18844
rect 4572 18900 4636 18904
rect 4572 18844 4576 18900
rect 4576 18844 4632 18900
rect 4632 18844 4636 18900
rect 4572 18840 4636 18844
rect 4652 18900 4716 18904
rect 4652 18844 4656 18900
rect 4656 18844 4712 18900
rect 4712 18844 4716 18900
rect 4652 18840 4716 18844
rect 4732 18900 4796 18904
rect 4732 18844 4736 18900
rect 4736 18844 4792 18900
rect 4792 18844 4796 18900
rect 4732 18840 4796 18844
rect 4812 18900 4876 18904
rect 4812 18844 4816 18900
rect 4816 18844 4872 18900
rect 4872 18844 4876 18900
rect 4812 18840 4876 18844
rect 4892 18900 4956 18904
rect 4892 18844 4896 18900
rect 4896 18844 4952 18900
rect 4952 18844 4956 18900
rect 4892 18840 4956 18844
rect 20990 18890 21054 18954
rect 43680 18900 43744 18904
rect 43680 18844 43684 18900
rect 43684 18844 43740 18900
rect 43740 18844 43744 18900
rect 43680 18840 43744 18844
rect 43760 18900 43824 18904
rect 43760 18844 43764 18900
rect 43764 18844 43820 18900
rect 43820 18844 43824 18900
rect 43760 18840 43824 18844
rect 43840 18900 43904 18904
rect 43840 18844 43844 18900
rect 43844 18844 43900 18900
rect 43900 18844 43904 18900
rect 43840 18840 43904 18844
rect 43920 18900 43984 18904
rect 43920 18844 43924 18900
rect 43924 18844 43980 18900
rect 43980 18844 43984 18900
rect 43920 18840 43984 18844
rect 44000 18900 44064 18904
rect 44000 18844 44004 18900
rect 44004 18844 44060 18900
rect 44060 18844 44064 18900
rect 44000 18840 44064 18844
rect 44080 18900 44144 18904
rect 44080 18844 44084 18900
rect 44084 18844 44140 18900
rect 44140 18844 44144 18900
rect 44080 18840 44144 18844
rect 44160 18900 44224 18904
rect 44160 18844 44164 18900
rect 44164 18844 44220 18900
rect 44220 18844 44224 18900
rect 44160 18840 44224 18844
rect 44240 18900 44304 18904
rect 44240 18844 44244 18900
rect 44244 18844 44300 18900
rect 44300 18844 44304 18900
rect 44240 18840 44304 18844
rect 44320 18900 44384 18904
rect 44320 18844 44324 18900
rect 44324 18844 44380 18900
rect 44380 18844 44384 18900
rect 44320 18840 44384 18844
rect 44400 18900 44464 18904
rect 44400 18844 44404 18900
rect 44404 18844 44460 18900
rect 44460 18844 44464 18900
rect 44400 18840 44464 18844
rect 44480 18900 44544 18904
rect 44480 18844 44484 18900
rect 44484 18844 44540 18900
rect 44540 18844 44544 18900
rect 44480 18840 44544 18844
rect 44560 18900 44624 18904
rect 44560 18844 44564 18900
rect 44564 18844 44620 18900
rect 44620 18844 44624 18900
rect 44560 18840 44624 18844
rect 44640 18900 44704 18904
rect 44640 18844 44644 18900
rect 44644 18844 44700 18900
rect 44700 18844 44704 18900
rect 44640 18840 44704 18844
rect 44720 18900 44784 18904
rect 44720 18844 44724 18900
rect 44724 18844 44780 18900
rect 44780 18844 44784 18900
rect 44720 18840 44784 18844
rect 44800 18900 44864 18904
rect 44800 18844 44804 18900
rect 44804 18844 44860 18900
rect 44860 18844 44864 18900
rect 44800 18840 44864 18844
rect 44880 18900 44944 18904
rect 44880 18844 44884 18900
rect 44884 18844 44940 18900
rect 44940 18844 44944 18900
rect 44880 18840 44944 18844
rect 44960 18900 45024 18904
rect 44960 18844 44964 18900
rect 44964 18844 45020 18900
rect 45020 18844 45024 18900
rect 44960 18840 45024 18844
rect 45040 18900 45104 18904
rect 45040 18844 45044 18900
rect 45044 18844 45100 18900
rect 45100 18844 45104 18900
rect 45040 18840 45104 18844
rect 45120 18900 45184 18904
rect 45120 18844 45124 18900
rect 45124 18844 45180 18900
rect 45180 18844 45184 18900
rect 45120 18840 45184 18844
rect 45200 18900 45264 18904
rect 45200 18844 45204 18900
rect 45204 18844 45260 18900
rect 45260 18844 45264 18900
rect 45200 18840 45264 18844
rect 16724 18550 16788 18614
rect 17443 18550 17507 18614
rect 18162 18550 18226 18614
rect 18881 18550 18945 18614
rect 19600 18550 19664 18614
rect 20319 18550 20383 18614
rect 21038 18550 21102 18614
rect 21757 18550 21821 18614
rect 22476 18550 22540 18614
rect 23195 18550 23259 18614
rect 16724 18470 16788 18534
rect 17443 18470 17507 18534
rect 18162 18470 18226 18534
rect 18881 18470 18945 18534
rect 19600 18470 19664 18534
rect 20319 18470 20383 18534
rect 21038 18470 21102 18534
rect 21757 18470 21821 18534
rect 22476 18470 22540 18534
rect 23195 18470 23259 18534
rect 16724 18390 16788 18454
rect 17443 18390 17507 18454
rect 18162 18390 18226 18454
rect 18881 18390 18945 18454
rect 19600 18390 19664 18454
rect 20319 18390 20383 18454
rect 21038 18390 21102 18454
rect 21757 18390 21821 18454
rect 22476 18390 22540 18454
rect 23195 18390 23259 18454
rect 16724 18310 16788 18374
rect 17443 18310 17507 18374
rect 18162 18310 18226 18374
rect 18881 18310 18945 18374
rect 19600 18310 19664 18374
rect 20319 18310 20383 18374
rect 21038 18310 21102 18374
rect 21757 18310 21821 18374
rect 22476 18310 22540 18374
rect 23195 18310 23259 18374
rect 16724 18230 16788 18294
rect 17443 18230 17507 18294
rect 18162 18230 18226 18294
rect 18881 18230 18945 18294
rect 19600 18230 19664 18294
rect 20319 18230 20383 18294
rect 21038 18230 21102 18294
rect 21757 18230 21821 18294
rect 22476 18230 22540 18294
rect 23195 18230 23259 18294
rect 16724 18150 16788 18214
rect 17443 18150 17507 18214
rect 18162 18150 18226 18214
rect 18881 18150 18945 18214
rect 19600 18150 19664 18214
rect 20319 18150 20383 18214
rect 21038 18150 21102 18214
rect 21757 18150 21821 18214
rect 22476 18150 22540 18214
rect 23195 18150 23259 18214
rect 16724 18070 16788 18134
rect 17443 18070 17507 18134
rect 18162 18070 18226 18134
rect 18881 18070 18945 18134
rect 19600 18070 19664 18134
rect 20319 18070 20383 18134
rect 21038 18070 21102 18134
rect 21757 18070 21821 18134
rect 22476 18070 22540 18134
rect 23195 18070 23259 18134
rect 16724 17850 16788 17914
rect 17443 17850 17507 17914
rect 18162 17850 18226 17914
rect 18881 17850 18945 17914
rect 19600 17850 19664 17914
rect 20319 17850 20383 17914
rect 21038 17850 21102 17914
rect 21757 17850 21821 17914
rect 22476 17850 22540 17914
rect 23195 17850 23259 17914
rect 16724 17770 16788 17834
rect 17443 17770 17507 17834
rect 18162 17770 18226 17834
rect 18881 17770 18945 17834
rect 19600 17770 19664 17834
rect 20319 17770 20383 17834
rect 21038 17770 21102 17834
rect 21757 17770 21821 17834
rect 22476 17770 22540 17834
rect 23195 17770 23259 17834
rect 16724 17690 16788 17754
rect 17443 17690 17507 17754
rect 18162 17690 18226 17754
rect 18881 17690 18945 17754
rect 19600 17690 19664 17754
rect 20319 17690 20383 17754
rect 21038 17690 21102 17754
rect 21757 17690 21821 17754
rect 22476 17690 22540 17754
rect 23195 17690 23259 17754
rect 16724 17610 16788 17674
rect 17443 17610 17507 17674
rect 18162 17610 18226 17674
rect 18881 17610 18945 17674
rect 19600 17610 19664 17674
rect 20319 17610 20383 17674
rect 21038 17610 21102 17674
rect 21757 17610 21821 17674
rect 22476 17610 22540 17674
rect 23195 17610 23259 17674
rect 16724 17530 16788 17594
rect 17443 17530 17507 17594
rect 18162 17530 18226 17594
rect 18881 17530 18945 17594
rect 19600 17530 19664 17594
rect 20319 17530 20383 17594
rect 21038 17530 21102 17594
rect 21757 17530 21821 17594
rect 22476 17530 22540 17594
rect 23195 17530 23259 17594
rect 16724 17450 16788 17514
rect 17443 17450 17507 17514
rect 18162 17450 18226 17514
rect 18881 17450 18945 17514
rect 19600 17450 19664 17514
rect 20319 17450 20383 17514
rect 21038 17450 21102 17514
rect 21757 17450 21821 17514
rect 22476 17450 22540 17514
rect 23195 17450 23259 17514
rect 16724 17370 16788 17434
rect 17443 17370 17507 17434
rect 18162 17370 18226 17434
rect 18881 17370 18945 17434
rect 19600 17370 19664 17434
rect 20319 17370 20383 17434
rect 21038 17370 21102 17434
rect 21757 17370 21821 17434
rect 22476 17370 22540 17434
rect 23195 17370 23259 17434
rect 16138 17210 16202 17214
rect 16218 17210 16282 17214
rect 16138 17154 16182 17210
rect 16182 17154 16202 17210
rect 16218 17154 16238 17210
rect 16238 17154 16282 17210
rect 16138 17150 16202 17154
rect 16218 17150 16282 17154
rect 924 17020 988 17024
rect 924 16964 928 17020
rect 928 16964 984 17020
rect 984 16964 988 17020
rect 924 16960 988 16964
rect 1004 17020 1068 17024
rect 1004 16964 1008 17020
rect 1008 16964 1064 17020
rect 1064 16964 1068 17020
rect 1004 16960 1068 16964
rect 1084 17020 1148 17024
rect 1084 16964 1088 17020
rect 1088 16964 1144 17020
rect 1144 16964 1148 17020
rect 1084 16960 1148 16964
rect 1164 17020 1228 17024
rect 1164 16964 1168 17020
rect 1168 16964 1224 17020
rect 1224 16964 1228 17020
rect 1164 16960 1228 16964
rect 1244 17020 1308 17024
rect 1244 16964 1248 17020
rect 1248 16964 1304 17020
rect 1304 16964 1308 17020
rect 1244 16960 1308 16964
rect 1324 17020 1388 17024
rect 1324 16964 1328 17020
rect 1328 16964 1384 17020
rect 1384 16964 1388 17020
rect 1324 16960 1388 16964
rect 1404 17020 1468 17024
rect 1404 16964 1408 17020
rect 1408 16964 1464 17020
rect 1464 16964 1468 17020
rect 1404 16960 1468 16964
rect 1484 17020 1548 17024
rect 1484 16964 1488 17020
rect 1488 16964 1544 17020
rect 1544 16964 1548 17020
rect 1484 16960 1548 16964
rect 1564 17020 1628 17024
rect 1564 16964 1568 17020
rect 1568 16964 1624 17020
rect 1624 16964 1628 17020
rect 1564 16960 1628 16964
rect 1644 17020 1708 17024
rect 1644 16964 1648 17020
rect 1648 16964 1704 17020
rect 1704 16964 1708 17020
rect 1644 16960 1708 16964
rect 1724 17020 1788 17024
rect 1724 16964 1728 17020
rect 1728 16964 1784 17020
rect 1784 16964 1788 17020
rect 1724 16960 1788 16964
rect 1804 17020 1868 17024
rect 1804 16964 1808 17020
rect 1808 16964 1864 17020
rect 1864 16964 1868 17020
rect 1804 16960 1868 16964
rect 1884 17020 1948 17024
rect 1884 16964 1888 17020
rect 1888 16964 1944 17020
rect 1944 16964 1948 17020
rect 1884 16960 1948 16964
rect 1964 17020 2028 17024
rect 1964 16964 1968 17020
rect 1968 16964 2024 17020
rect 2024 16964 2028 17020
rect 1964 16960 2028 16964
rect 2044 17020 2108 17024
rect 2044 16964 2048 17020
rect 2048 16964 2104 17020
rect 2104 16964 2108 17020
rect 2044 16960 2108 16964
rect 2124 17020 2188 17024
rect 2124 16964 2128 17020
rect 2128 16964 2184 17020
rect 2184 16964 2188 17020
rect 2124 16960 2188 16964
rect 2204 17020 2268 17024
rect 2204 16964 2208 17020
rect 2208 16964 2264 17020
rect 2264 16964 2268 17020
rect 2204 16960 2268 16964
rect 2284 17020 2348 17024
rect 2284 16964 2288 17020
rect 2288 16964 2344 17020
rect 2344 16964 2348 17020
rect 2284 16960 2348 16964
rect 2364 17020 2428 17024
rect 2364 16964 2368 17020
rect 2368 16964 2424 17020
rect 2424 16964 2428 17020
rect 2364 16960 2428 16964
rect 2444 17020 2508 17024
rect 2444 16964 2448 17020
rect 2448 16964 2504 17020
rect 2504 16964 2508 17020
rect 2444 16960 2508 16964
rect 17402 16998 17466 17002
rect 17402 16942 17406 16998
rect 17406 16942 17462 16998
rect 17462 16942 17466 16998
rect 17402 16938 17466 16942
rect 46128 17020 46192 17024
rect 46128 16964 46132 17020
rect 46132 16964 46188 17020
rect 46188 16964 46192 17020
rect 46128 16960 46192 16964
rect 46208 17020 46272 17024
rect 46208 16964 46212 17020
rect 46212 16964 46268 17020
rect 46268 16964 46272 17020
rect 46208 16960 46272 16964
rect 46288 17020 46352 17024
rect 46288 16964 46292 17020
rect 46292 16964 46348 17020
rect 46348 16964 46352 17020
rect 46288 16960 46352 16964
rect 46368 17020 46432 17024
rect 46368 16964 46372 17020
rect 46372 16964 46428 17020
rect 46428 16964 46432 17020
rect 46368 16960 46432 16964
rect 46448 17020 46512 17024
rect 46448 16964 46452 17020
rect 46452 16964 46508 17020
rect 46508 16964 46512 17020
rect 46448 16960 46512 16964
rect 46528 17020 46592 17024
rect 46528 16964 46532 17020
rect 46532 16964 46588 17020
rect 46588 16964 46592 17020
rect 46528 16960 46592 16964
rect 46608 17020 46672 17024
rect 46608 16964 46612 17020
rect 46612 16964 46668 17020
rect 46668 16964 46672 17020
rect 46608 16960 46672 16964
rect 46688 17020 46752 17024
rect 46688 16964 46692 17020
rect 46692 16964 46748 17020
rect 46748 16964 46752 17020
rect 46688 16960 46752 16964
rect 46768 17020 46832 17024
rect 46768 16964 46772 17020
rect 46772 16964 46828 17020
rect 46828 16964 46832 17020
rect 46768 16960 46832 16964
rect 46848 17020 46912 17024
rect 46848 16964 46852 17020
rect 46852 16964 46908 17020
rect 46908 16964 46912 17020
rect 46848 16960 46912 16964
rect 46928 17020 46992 17024
rect 46928 16964 46932 17020
rect 46932 16964 46988 17020
rect 46988 16964 46992 17020
rect 46928 16960 46992 16964
rect 47008 17020 47072 17024
rect 47008 16964 47012 17020
rect 47012 16964 47068 17020
rect 47068 16964 47072 17020
rect 47008 16960 47072 16964
rect 47088 17020 47152 17024
rect 47088 16964 47092 17020
rect 47092 16964 47148 17020
rect 47148 16964 47152 17020
rect 47088 16960 47152 16964
rect 47168 17020 47232 17024
rect 47168 16964 47172 17020
rect 47172 16964 47228 17020
rect 47228 16964 47232 17020
rect 47168 16960 47232 16964
rect 47248 17020 47312 17024
rect 47248 16964 47252 17020
rect 47252 16964 47308 17020
rect 47308 16964 47312 17020
rect 47248 16960 47312 16964
rect 47328 17020 47392 17024
rect 47328 16964 47332 17020
rect 47332 16964 47388 17020
rect 47388 16964 47392 17020
rect 47328 16960 47392 16964
rect 47408 17020 47472 17024
rect 47408 16964 47412 17020
rect 47412 16964 47468 17020
rect 47468 16964 47472 17020
rect 47408 16960 47472 16964
rect 47488 17020 47552 17024
rect 47488 16964 47492 17020
rect 47492 16964 47548 17020
rect 47548 16964 47552 17020
rect 47488 16960 47552 16964
rect 47568 17020 47632 17024
rect 47568 16964 47572 17020
rect 47572 16964 47628 17020
rect 47628 16964 47632 17020
rect 47568 16960 47632 16964
rect 47648 17020 47712 17024
rect 47648 16964 47652 17020
rect 47652 16964 47708 17020
rect 47708 16964 47712 17020
rect 47648 16960 47712 16964
rect 19610 16328 19674 16392
rect 3372 15140 3436 15144
rect 3372 15084 3376 15140
rect 3376 15084 3432 15140
rect 3432 15084 3436 15140
rect 3372 15080 3436 15084
rect 3452 15140 3516 15144
rect 3452 15084 3456 15140
rect 3456 15084 3512 15140
rect 3512 15084 3516 15140
rect 3452 15080 3516 15084
rect 3532 15140 3596 15144
rect 3532 15084 3536 15140
rect 3536 15084 3592 15140
rect 3592 15084 3596 15140
rect 3532 15080 3596 15084
rect 3612 15140 3676 15144
rect 3612 15084 3616 15140
rect 3616 15084 3672 15140
rect 3672 15084 3676 15140
rect 3612 15080 3676 15084
rect 3692 15140 3756 15144
rect 3692 15084 3696 15140
rect 3696 15084 3752 15140
rect 3752 15084 3756 15140
rect 3692 15080 3756 15084
rect 3772 15140 3836 15144
rect 3772 15084 3776 15140
rect 3776 15084 3832 15140
rect 3832 15084 3836 15140
rect 3772 15080 3836 15084
rect 3852 15140 3916 15144
rect 3852 15084 3856 15140
rect 3856 15084 3912 15140
rect 3912 15084 3916 15140
rect 3852 15080 3916 15084
rect 3932 15140 3996 15144
rect 3932 15084 3936 15140
rect 3936 15084 3992 15140
rect 3992 15084 3996 15140
rect 3932 15080 3996 15084
rect 4012 15140 4076 15144
rect 4012 15084 4016 15140
rect 4016 15084 4072 15140
rect 4072 15084 4076 15140
rect 4012 15080 4076 15084
rect 4092 15140 4156 15144
rect 4092 15084 4096 15140
rect 4096 15084 4152 15140
rect 4152 15084 4156 15140
rect 4092 15080 4156 15084
rect 4172 15140 4236 15144
rect 4172 15084 4176 15140
rect 4176 15084 4232 15140
rect 4232 15084 4236 15140
rect 4172 15080 4236 15084
rect 4252 15140 4316 15144
rect 4252 15084 4256 15140
rect 4256 15084 4312 15140
rect 4312 15084 4316 15140
rect 4252 15080 4316 15084
rect 4332 15140 4396 15144
rect 4332 15084 4336 15140
rect 4336 15084 4392 15140
rect 4392 15084 4396 15140
rect 4332 15080 4396 15084
rect 4412 15140 4476 15144
rect 4412 15084 4416 15140
rect 4416 15084 4472 15140
rect 4472 15084 4476 15140
rect 4412 15080 4476 15084
rect 4492 15140 4556 15144
rect 4492 15084 4496 15140
rect 4496 15084 4552 15140
rect 4552 15084 4556 15140
rect 4492 15080 4556 15084
rect 4572 15140 4636 15144
rect 4572 15084 4576 15140
rect 4576 15084 4632 15140
rect 4632 15084 4636 15140
rect 4572 15080 4636 15084
rect 4652 15140 4716 15144
rect 4652 15084 4656 15140
rect 4656 15084 4712 15140
rect 4712 15084 4716 15140
rect 4652 15080 4716 15084
rect 4732 15140 4796 15144
rect 4732 15084 4736 15140
rect 4736 15084 4792 15140
rect 4792 15084 4796 15140
rect 4732 15080 4796 15084
rect 4812 15140 4876 15144
rect 4812 15084 4816 15140
rect 4816 15084 4872 15140
rect 4872 15084 4876 15140
rect 4812 15080 4876 15084
rect 4892 15140 4956 15144
rect 4892 15084 4896 15140
rect 4896 15084 4952 15140
rect 4952 15084 4956 15140
rect 4892 15080 4956 15084
rect 43680 15140 43744 15144
rect 43680 15084 43684 15140
rect 43684 15084 43740 15140
rect 43740 15084 43744 15140
rect 43680 15080 43744 15084
rect 43760 15140 43824 15144
rect 43760 15084 43764 15140
rect 43764 15084 43820 15140
rect 43820 15084 43824 15140
rect 43760 15080 43824 15084
rect 43840 15140 43904 15144
rect 43840 15084 43844 15140
rect 43844 15084 43900 15140
rect 43900 15084 43904 15140
rect 43840 15080 43904 15084
rect 43920 15140 43984 15144
rect 43920 15084 43924 15140
rect 43924 15084 43980 15140
rect 43980 15084 43984 15140
rect 43920 15080 43984 15084
rect 44000 15140 44064 15144
rect 44000 15084 44004 15140
rect 44004 15084 44060 15140
rect 44060 15084 44064 15140
rect 44000 15080 44064 15084
rect 44080 15140 44144 15144
rect 44080 15084 44084 15140
rect 44084 15084 44140 15140
rect 44140 15084 44144 15140
rect 44080 15080 44144 15084
rect 44160 15140 44224 15144
rect 44160 15084 44164 15140
rect 44164 15084 44220 15140
rect 44220 15084 44224 15140
rect 44160 15080 44224 15084
rect 44240 15140 44304 15144
rect 44240 15084 44244 15140
rect 44244 15084 44300 15140
rect 44300 15084 44304 15140
rect 44240 15080 44304 15084
rect 44320 15140 44384 15144
rect 44320 15084 44324 15140
rect 44324 15084 44380 15140
rect 44380 15084 44384 15140
rect 44320 15080 44384 15084
rect 44400 15140 44464 15144
rect 44400 15084 44404 15140
rect 44404 15084 44460 15140
rect 44460 15084 44464 15140
rect 44400 15080 44464 15084
rect 44480 15140 44544 15144
rect 44480 15084 44484 15140
rect 44484 15084 44540 15140
rect 44540 15084 44544 15140
rect 44480 15080 44544 15084
rect 44560 15140 44624 15144
rect 44560 15084 44564 15140
rect 44564 15084 44620 15140
rect 44620 15084 44624 15140
rect 44560 15080 44624 15084
rect 44640 15140 44704 15144
rect 44640 15084 44644 15140
rect 44644 15084 44700 15140
rect 44700 15084 44704 15140
rect 44640 15080 44704 15084
rect 44720 15140 44784 15144
rect 44720 15084 44724 15140
rect 44724 15084 44780 15140
rect 44780 15084 44784 15140
rect 44720 15080 44784 15084
rect 44800 15140 44864 15144
rect 44800 15084 44804 15140
rect 44804 15084 44860 15140
rect 44860 15084 44864 15140
rect 44800 15080 44864 15084
rect 44880 15140 44944 15144
rect 44880 15084 44884 15140
rect 44884 15084 44940 15140
rect 44940 15084 44944 15140
rect 44880 15080 44944 15084
rect 44960 15140 45024 15144
rect 44960 15084 44964 15140
rect 44964 15084 45020 15140
rect 45020 15084 45024 15140
rect 44960 15080 45024 15084
rect 45040 15140 45104 15144
rect 45040 15084 45044 15140
rect 45044 15084 45100 15140
rect 45100 15084 45104 15140
rect 45040 15080 45104 15084
rect 45120 15140 45184 15144
rect 45120 15084 45124 15140
rect 45124 15084 45180 15140
rect 45180 15084 45184 15140
rect 45120 15080 45184 15084
rect 45200 15140 45264 15144
rect 45200 15084 45204 15140
rect 45204 15084 45260 15140
rect 45260 15084 45264 15140
rect 45200 15080 45264 15084
rect 16724 14790 16788 14854
rect 17443 14790 17507 14854
rect 18162 14790 18226 14854
rect 18881 14790 18945 14854
rect 19600 14790 19664 14854
rect 20319 14790 20383 14854
rect 21038 14790 21102 14854
rect 21757 14790 21821 14854
rect 22476 14790 22540 14854
rect 23195 14790 23259 14854
rect 16724 14710 16788 14774
rect 17443 14710 17507 14774
rect 18162 14710 18226 14774
rect 18881 14710 18945 14774
rect 19600 14710 19664 14774
rect 20319 14710 20383 14774
rect 21038 14710 21102 14774
rect 21757 14710 21821 14774
rect 22476 14710 22540 14774
rect 23195 14710 23259 14774
rect 16724 14630 16788 14694
rect 17443 14630 17507 14694
rect 18162 14630 18226 14694
rect 18881 14630 18945 14694
rect 19600 14630 19664 14694
rect 20319 14630 20383 14694
rect 21038 14630 21102 14694
rect 21757 14630 21821 14694
rect 22476 14630 22540 14694
rect 23195 14630 23259 14694
rect 16724 14550 16788 14614
rect 17443 14550 17507 14614
rect 18162 14550 18226 14614
rect 18881 14550 18945 14614
rect 19600 14550 19664 14614
rect 20319 14550 20383 14614
rect 21038 14550 21102 14614
rect 21757 14550 21821 14614
rect 22476 14550 22540 14614
rect 23195 14550 23259 14614
rect 16724 14470 16788 14534
rect 17443 14470 17507 14534
rect 18162 14470 18226 14534
rect 18881 14470 18945 14534
rect 19600 14470 19664 14534
rect 20319 14470 20383 14534
rect 21038 14470 21102 14534
rect 21757 14470 21821 14534
rect 22476 14470 22540 14534
rect 23195 14470 23259 14534
rect 16724 14390 16788 14454
rect 17443 14390 17507 14454
rect 18162 14390 18226 14454
rect 18881 14390 18945 14454
rect 19600 14390 19664 14454
rect 20319 14390 20383 14454
rect 21038 14390 21102 14454
rect 21757 14390 21821 14454
rect 22476 14390 22540 14454
rect 23195 14390 23259 14454
rect 16724 14310 16788 14374
rect 17443 14310 17507 14374
rect 18162 14310 18226 14374
rect 18881 14310 18945 14374
rect 19600 14310 19664 14374
rect 20319 14310 20383 14374
rect 21038 14310 21102 14374
rect 21757 14310 21821 14374
rect 22476 14310 22540 14374
rect 23195 14310 23259 14374
rect 16724 14090 16788 14154
rect 17443 14090 17507 14154
rect 18162 14090 18226 14154
rect 18881 14090 18945 14154
rect 19600 14090 19664 14154
rect 20319 14090 20383 14154
rect 21038 14090 21102 14154
rect 21757 14090 21821 14154
rect 22476 14090 22540 14154
rect 23195 14090 23259 14154
rect 16724 14010 16788 14074
rect 17443 14010 17507 14074
rect 18162 14010 18226 14074
rect 18881 14010 18945 14074
rect 19600 14010 19664 14074
rect 20319 14010 20383 14074
rect 21038 14010 21102 14074
rect 21757 14010 21821 14074
rect 22476 14010 22540 14074
rect 23195 14010 23259 14074
rect 16724 13930 16788 13994
rect 17443 13930 17507 13994
rect 18162 13930 18226 13994
rect 18881 13930 18945 13994
rect 19600 13930 19664 13994
rect 20319 13930 20383 13994
rect 21038 13930 21102 13994
rect 21757 13930 21821 13994
rect 22476 13930 22540 13994
rect 23195 13930 23259 13994
rect 16724 13850 16788 13914
rect 17443 13850 17507 13914
rect 18162 13850 18226 13914
rect 18881 13850 18945 13914
rect 19600 13850 19664 13914
rect 20319 13850 20383 13914
rect 21038 13850 21102 13914
rect 21757 13850 21821 13914
rect 22476 13850 22540 13914
rect 23195 13850 23259 13914
rect 16724 13770 16788 13834
rect 17443 13770 17507 13834
rect 18162 13770 18226 13834
rect 18881 13770 18945 13834
rect 19600 13770 19664 13834
rect 20319 13770 20383 13834
rect 21038 13770 21102 13834
rect 21757 13770 21821 13834
rect 22476 13770 22540 13834
rect 23195 13770 23259 13834
rect 16724 13690 16788 13754
rect 17443 13690 17507 13754
rect 18162 13690 18226 13754
rect 18881 13690 18945 13754
rect 19600 13690 19664 13754
rect 20319 13690 20383 13754
rect 21038 13690 21102 13754
rect 21757 13690 21821 13754
rect 22476 13690 22540 13754
rect 23195 13690 23259 13754
rect 16724 13610 16788 13674
rect 17443 13610 17507 13674
rect 18162 13610 18226 13674
rect 18881 13610 18945 13674
rect 19600 13610 19664 13674
rect 20319 13610 20383 13674
rect 21038 13610 21102 13674
rect 21757 13610 21821 13674
rect 22476 13610 22540 13674
rect 23195 13610 23259 13674
rect 16138 13450 16202 13454
rect 16218 13450 16282 13454
rect 16138 13394 16182 13450
rect 16182 13394 16202 13450
rect 16218 13394 16238 13450
rect 16238 13394 16282 13450
rect 16138 13390 16202 13394
rect 16218 13390 16282 13394
rect 17264 13400 17328 13464
rect 924 13260 988 13264
rect 924 13204 928 13260
rect 928 13204 984 13260
rect 984 13204 988 13260
rect 924 13200 988 13204
rect 1004 13260 1068 13264
rect 1004 13204 1008 13260
rect 1008 13204 1064 13260
rect 1064 13204 1068 13260
rect 1004 13200 1068 13204
rect 1084 13260 1148 13264
rect 1084 13204 1088 13260
rect 1088 13204 1144 13260
rect 1144 13204 1148 13260
rect 1084 13200 1148 13204
rect 1164 13260 1228 13264
rect 1164 13204 1168 13260
rect 1168 13204 1224 13260
rect 1224 13204 1228 13260
rect 1164 13200 1228 13204
rect 1244 13260 1308 13264
rect 1244 13204 1248 13260
rect 1248 13204 1304 13260
rect 1304 13204 1308 13260
rect 1244 13200 1308 13204
rect 1324 13260 1388 13264
rect 1324 13204 1328 13260
rect 1328 13204 1384 13260
rect 1384 13204 1388 13260
rect 1324 13200 1388 13204
rect 1404 13260 1468 13264
rect 1404 13204 1408 13260
rect 1408 13204 1464 13260
rect 1464 13204 1468 13260
rect 1404 13200 1468 13204
rect 1484 13260 1548 13264
rect 1484 13204 1488 13260
rect 1488 13204 1544 13260
rect 1544 13204 1548 13260
rect 1484 13200 1548 13204
rect 1564 13260 1628 13264
rect 1564 13204 1568 13260
rect 1568 13204 1624 13260
rect 1624 13204 1628 13260
rect 1564 13200 1628 13204
rect 1644 13260 1708 13264
rect 1644 13204 1648 13260
rect 1648 13204 1704 13260
rect 1704 13204 1708 13260
rect 1644 13200 1708 13204
rect 1724 13260 1788 13264
rect 1724 13204 1728 13260
rect 1728 13204 1784 13260
rect 1784 13204 1788 13260
rect 1724 13200 1788 13204
rect 1804 13260 1868 13264
rect 1804 13204 1808 13260
rect 1808 13204 1864 13260
rect 1864 13204 1868 13260
rect 1804 13200 1868 13204
rect 1884 13260 1948 13264
rect 1884 13204 1888 13260
rect 1888 13204 1944 13260
rect 1944 13204 1948 13260
rect 1884 13200 1948 13204
rect 1964 13260 2028 13264
rect 1964 13204 1968 13260
rect 1968 13204 2024 13260
rect 2024 13204 2028 13260
rect 1964 13200 2028 13204
rect 2044 13260 2108 13264
rect 2044 13204 2048 13260
rect 2048 13204 2104 13260
rect 2104 13204 2108 13260
rect 2044 13200 2108 13204
rect 2124 13260 2188 13264
rect 2124 13204 2128 13260
rect 2128 13204 2184 13260
rect 2184 13204 2188 13260
rect 2124 13200 2188 13204
rect 2204 13260 2268 13264
rect 2204 13204 2208 13260
rect 2208 13204 2264 13260
rect 2264 13204 2268 13260
rect 2204 13200 2268 13204
rect 2284 13260 2348 13264
rect 2284 13204 2288 13260
rect 2288 13204 2344 13260
rect 2344 13204 2348 13260
rect 2284 13200 2348 13204
rect 2364 13260 2428 13264
rect 2364 13204 2368 13260
rect 2368 13204 2424 13260
rect 2424 13204 2428 13260
rect 2364 13200 2428 13204
rect 2444 13260 2508 13264
rect 2444 13204 2448 13260
rect 2448 13204 2504 13260
rect 2504 13204 2508 13260
rect 2444 13200 2508 13204
rect 46128 13260 46192 13264
rect 46128 13204 46132 13260
rect 46132 13204 46188 13260
rect 46188 13204 46192 13260
rect 46128 13200 46192 13204
rect 46208 13260 46272 13264
rect 46208 13204 46212 13260
rect 46212 13204 46268 13260
rect 46268 13204 46272 13260
rect 46208 13200 46272 13204
rect 46288 13260 46352 13264
rect 46288 13204 46292 13260
rect 46292 13204 46348 13260
rect 46348 13204 46352 13260
rect 46288 13200 46352 13204
rect 46368 13260 46432 13264
rect 46368 13204 46372 13260
rect 46372 13204 46428 13260
rect 46428 13204 46432 13260
rect 46368 13200 46432 13204
rect 46448 13260 46512 13264
rect 46448 13204 46452 13260
rect 46452 13204 46508 13260
rect 46508 13204 46512 13260
rect 46448 13200 46512 13204
rect 46528 13260 46592 13264
rect 46528 13204 46532 13260
rect 46532 13204 46588 13260
rect 46588 13204 46592 13260
rect 46528 13200 46592 13204
rect 46608 13260 46672 13264
rect 46608 13204 46612 13260
rect 46612 13204 46668 13260
rect 46668 13204 46672 13260
rect 46608 13200 46672 13204
rect 46688 13260 46752 13264
rect 46688 13204 46692 13260
rect 46692 13204 46748 13260
rect 46748 13204 46752 13260
rect 46688 13200 46752 13204
rect 46768 13260 46832 13264
rect 46768 13204 46772 13260
rect 46772 13204 46828 13260
rect 46828 13204 46832 13260
rect 46768 13200 46832 13204
rect 46848 13260 46912 13264
rect 46848 13204 46852 13260
rect 46852 13204 46908 13260
rect 46908 13204 46912 13260
rect 46848 13200 46912 13204
rect 46928 13260 46992 13264
rect 46928 13204 46932 13260
rect 46932 13204 46988 13260
rect 46988 13204 46992 13260
rect 46928 13200 46992 13204
rect 47008 13260 47072 13264
rect 47008 13204 47012 13260
rect 47012 13204 47068 13260
rect 47068 13204 47072 13260
rect 47008 13200 47072 13204
rect 47088 13260 47152 13264
rect 47088 13204 47092 13260
rect 47092 13204 47148 13260
rect 47148 13204 47152 13260
rect 47088 13200 47152 13204
rect 47168 13260 47232 13264
rect 47168 13204 47172 13260
rect 47172 13204 47228 13260
rect 47228 13204 47232 13260
rect 47168 13200 47232 13204
rect 47248 13260 47312 13264
rect 47248 13204 47252 13260
rect 47252 13204 47308 13260
rect 47308 13204 47312 13260
rect 47248 13200 47312 13204
rect 47328 13260 47392 13264
rect 47328 13204 47332 13260
rect 47332 13204 47388 13260
rect 47388 13204 47392 13260
rect 47328 13200 47392 13204
rect 47408 13260 47472 13264
rect 47408 13204 47412 13260
rect 47412 13204 47468 13260
rect 47468 13204 47472 13260
rect 47408 13200 47472 13204
rect 47488 13260 47552 13264
rect 47488 13204 47492 13260
rect 47492 13204 47548 13260
rect 47548 13204 47552 13260
rect 47488 13200 47552 13204
rect 47568 13260 47632 13264
rect 47568 13204 47572 13260
rect 47572 13204 47628 13260
rect 47628 13204 47632 13260
rect 47568 13200 47632 13204
rect 47648 13260 47712 13264
rect 47648 13204 47652 13260
rect 47652 13204 47708 13260
rect 47708 13204 47712 13260
rect 47648 13200 47712 13204
rect 3372 11380 3436 11384
rect 3372 11324 3376 11380
rect 3376 11324 3432 11380
rect 3432 11324 3436 11380
rect 3372 11320 3436 11324
rect 3452 11380 3516 11384
rect 3452 11324 3456 11380
rect 3456 11324 3512 11380
rect 3512 11324 3516 11380
rect 3452 11320 3516 11324
rect 3532 11380 3596 11384
rect 3532 11324 3536 11380
rect 3536 11324 3592 11380
rect 3592 11324 3596 11380
rect 3532 11320 3596 11324
rect 3612 11380 3676 11384
rect 3612 11324 3616 11380
rect 3616 11324 3672 11380
rect 3672 11324 3676 11380
rect 3612 11320 3676 11324
rect 3692 11380 3756 11384
rect 3692 11324 3696 11380
rect 3696 11324 3752 11380
rect 3752 11324 3756 11380
rect 3692 11320 3756 11324
rect 3772 11380 3836 11384
rect 3772 11324 3776 11380
rect 3776 11324 3832 11380
rect 3832 11324 3836 11380
rect 3772 11320 3836 11324
rect 3852 11380 3916 11384
rect 3852 11324 3856 11380
rect 3856 11324 3912 11380
rect 3912 11324 3916 11380
rect 3852 11320 3916 11324
rect 3932 11380 3996 11384
rect 3932 11324 3936 11380
rect 3936 11324 3992 11380
rect 3992 11324 3996 11380
rect 3932 11320 3996 11324
rect 4012 11380 4076 11384
rect 4012 11324 4016 11380
rect 4016 11324 4072 11380
rect 4072 11324 4076 11380
rect 4012 11320 4076 11324
rect 4092 11380 4156 11384
rect 4092 11324 4096 11380
rect 4096 11324 4152 11380
rect 4152 11324 4156 11380
rect 4092 11320 4156 11324
rect 4172 11380 4236 11384
rect 4172 11324 4176 11380
rect 4176 11324 4232 11380
rect 4232 11324 4236 11380
rect 4172 11320 4236 11324
rect 4252 11380 4316 11384
rect 4252 11324 4256 11380
rect 4256 11324 4312 11380
rect 4312 11324 4316 11380
rect 4252 11320 4316 11324
rect 4332 11380 4396 11384
rect 4332 11324 4336 11380
rect 4336 11324 4392 11380
rect 4392 11324 4396 11380
rect 4332 11320 4396 11324
rect 4412 11380 4476 11384
rect 4412 11324 4416 11380
rect 4416 11324 4472 11380
rect 4472 11324 4476 11380
rect 4412 11320 4476 11324
rect 4492 11380 4556 11384
rect 4492 11324 4496 11380
rect 4496 11324 4552 11380
rect 4552 11324 4556 11380
rect 4492 11320 4556 11324
rect 4572 11380 4636 11384
rect 4572 11324 4576 11380
rect 4576 11324 4632 11380
rect 4632 11324 4636 11380
rect 4572 11320 4636 11324
rect 4652 11380 4716 11384
rect 4652 11324 4656 11380
rect 4656 11324 4712 11380
rect 4712 11324 4716 11380
rect 4652 11320 4716 11324
rect 4732 11380 4796 11384
rect 4732 11324 4736 11380
rect 4736 11324 4792 11380
rect 4792 11324 4796 11380
rect 4732 11320 4796 11324
rect 4812 11380 4876 11384
rect 4812 11324 4816 11380
rect 4816 11324 4872 11380
rect 4872 11324 4876 11380
rect 4812 11320 4876 11324
rect 4892 11380 4956 11384
rect 4892 11324 4896 11380
rect 4896 11324 4952 11380
rect 4952 11324 4956 11380
rect 4892 11320 4956 11324
rect 43680 11380 43744 11384
rect 43680 11324 43684 11380
rect 43684 11324 43740 11380
rect 43740 11324 43744 11380
rect 43680 11320 43744 11324
rect 43760 11380 43824 11384
rect 43760 11324 43764 11380
rect 43764 11324 43820 11380
rect 43820 11324 43824 11380
rect 43760 11320 43824 11324
rect 43840 11380 43904 11384
rect 43840 11324 43844 11380
rect 43844 11324 43900 11380
rect 43900 11324 43904 11380
rect 43840 11320 43904 11324
rect 43920 11380 43984 11384
rect 43920 11324 43924 11380
rect 43924 11324 43980 11380
rect 43980 11324 43984 11380
rect 43920 11320 43984 11324
rect 44000 11380 44064 11384
rect 44000 11324 44004 11380
rect 44004 11324 44060 11380
rect 44060 11324 44064 11380
rect 44000 11320 44064 11324
rect 44080 11380 44144 11384
rect 44080 11324 44084 11380
rect 44084 11324 44140 11380
rect 44140 11324 44144 11380
rect 44080 11320 44144 11324
rect 44160 11380 44224 11384
rect 44160 11324 44164 11380
rect 44164 11324 44220 11380
rect 44220 11324 44224 11380
rect 44160 11320 44224 11324
rect 44240 11380 44304 11384
rect 44240 11324 44244 11380
rect 44244 11324 44300 11380
rect 44300 11324 44304 11380
rect 44240 11320 44304 11324
rect 44320 11380 44384 11384
rect 44320 11324 44324 11380
rect 44324 11324 44380 11380
rect 44380 11324 44384 11380
rect 44320 11320 44384 11324
rect 44400 11380 44464 11384
rect 44400 11324 44404 11380
rect 44404 11324 44460 11380
rect 44460 11324 44464 11380
rect 44400 11320 44464 11324
rect 44480 11380 44544 11384
rect 44480 11324 44484 11380
rect 44484 11324 44540 11380
rect 44540 11324 44544 11380
rect 44480 11320 44544 11324
rect 44560 11380 44624 11384
rect 44560 11324 44564 11380
rect 44564 11324 44620 11380
rect 44620 11324 44624 11380
rect 44560 11320 44624 11324
rect 44640 11380 44704 11384
rect 44640 11324 44644 11380
rect 44644 11324 44700 11380
rect 44700 11324 44704 11380
rect 44640 11320 44704 11324
rect 44720 11380 44784 11384
rect 44720 11324 44724 11380
rect 44724 11324 44780 11380
rect 44780 11324 44784 11380
rect 44720 11320 44784 11324
rect 44800 11380 44864 11384
rect 44800 11324 44804 11380
rect 44804 11324 44860 11380
rect 44860 11324 44864 11380
rect 44800 11320 44864 11324
rect 44880 11380 44944 11384
rect 44880 11324 44884 11380
rect 44884 11324 44940 11380
rect 44940 11324 44944 11380
rect 44880 11320 44944 11324
rect 44960 11380 45024 11384
rect 44960 11324 44964 11380
rect 44964 11324 45020 11380
rect 45020 11324 45024 11380
rect 44960 11320 45024 11324
rect 45040 11380 45104 11384
rect 45040 11324 45044 11380
rect 45044 11324 45100 11380
rect 45100 11324 45104 11380
rect 45040 11320 45104 11324
rect 45120 11380 45184 11384
rect 45120 11324 45124 11380
rect 45124 11324 45180 11380
rect 45180 11324 45184 11380
rect 45120 11320 45184 11324
rect 45200 11380 45264 11384
rect 45200 11324 45204 11380
rect 45204 11324 45260 11380
rect 45260 11324 45264 11380
rect 45200 11320 45264 11324
rect 16724 11030 16788 11094
rect 17443 11030 17507 11094
rect 18162 11030 18226 11094
rect 18881 11030 18945 11094
rect 19600 11030 19664 11094
rect 20319 11030 20383 11094
rect 21038 11030 21102 11094
rect 21757 11030 21821 11094
rect 22476 11030 22540 11094
rect 23195 11030 23259 11094
rect 23474 11082 23538 11146
rect 16724 10950 16788 11014
rect 17443 10950 17507 11014
rect 18162 10950 18226 11014
rect 18881 10950 18945 11014
rect 19600 10950 19664 11014
rect 20319 10950 20383 11014
rect 21038 10950 21102 11014
rect 21757 10950 21821 11014
rect 22476 10950 22540 11014
rect 23195 10950 23259 11014
rect 16724 10870 16788 10934
rect 17443 10870 17507 10934
rect 18162 10870 18226 10934
rect 18881 10870 18945 10934
rect 19600 10870 19664 10934
rect 20319 10870 20383 10934
rect 21038 10870 21102 10934
rect 21757 10870 21821 10934
rect 22476 10870 22540 10934
rect 23195 10870 23259 10934
rect 16724 10790 16788 10854
rect 17443 10790 17507 10854
rect 18162 10790 18226 10854
rect 18881 10790 18945 10854
rect 19600 10790 19664 10854
rect 20319 10790 20383 10854
rect 21038 10790 21102 10854
rect 21757 10790 21821 10854
rect 22476 10790 22540 10854
rect 23195 10790 23259 10854
rect 16724 10710 16788 10774
rect 17443 10710 17507 10774
rect 18162 10710 18226 10774
rect 18881 10710 18945 10774
rect 19600 10710 19664 10774
rect 20319 10710 20383 10774
rect 21038 10710 21102 10774
rect 21757 10710 21821 10774
rect 22476 10710 22540 10774
rect 23195 10710 23259 10774
rect 16724 10630 16788 10694
rect 17443 10630 17507 10694
rect 18162 10630 18226 10694
rect 18881 10630 18945 10694
rect 19600 10630 19664 10694
rect 20319 10630 20383 10694
rect 21038 10630 21102 10694
rect 21757 10630 21821 10694
rect 22476 10630 22540 10694
rect 23195 10630 23259 10694
rect 16724 10550 16788 10614
rect 17443 10550 17507 10614
rect 18162 10550 18226 10614
rect 18881 10550 18945 10614
rect 19600 10550 19664 10614
rect 20319 10550 20383 10614
rect 21038 10550 21102 10614
rect 21757 10550 21821 10614
rect 22476 10550 22540 10614
rect 23195 10550 23259 10614
rect 16724 10330 16788 10394
rect 17443 10330 17507 10394
rect 18162 10330 18226 10394
rect 18881 10330 18945 10394
rect 19600 10330 19664 10394
rect 20319 10330 20383 10394
rect 21038 10330 21102 10394
rect 21757 10330 21821 10394
rect 22476 10330 22540 10394
rect 23195 10330 23259 10394
rect 16724 10250 16788 10314
rect 17443 10250 17507 10314
rect 18162 10250 18226 10314
rect 18881 10250 18945 10314
rect 19600 10250 19664 10314
rect 20319 10250 20383 10314
rect 21038 10250 21102 10314
rect 21757 10250 21821 10314
rect 22476 10250 22540 10314
rect 23195 10250 23259 10314
rect 16724 10170 16788 10234
rect 17443 10170 17507 10234
rect 18162 10170 18226 10234
rect 18881 10170 18945 10234
rect 19600 10170 19664 10234
rect 20319 10170 20383 10234
rect 21038 10170 21102 10234
rect 21757 10170 21821 10234
rect 22476 10170 22540 10234
rect 23195 10170 23259 10234
rect 16724 10090 16788 10154
rect 17443 10090 17507 10154
rect 18162 10090 18226 10154
rect 18881 10090 18945 10154
rect 19600 10090 19664 10154
rect 20319 10090 20383 10154
rect 21038 10090 21102 10154
rect 21757 10090 21821 10154
rect 22476 10090 22540 10154
rect 23195 10090 23259 10154
rect 16724 10010 16788 10074
rect 17443 10010 17507 10074
rect 18162 10010 18226 10074
rect 18881 10010 18945 10074
rect 19600 10010 19664 10074
rect 20319 10010 20383 10074
rect 21038 10010 21102 10074
rect 21757 10010 21821 10074
rect 22476 10010 22540 10074
rect 23195 10010 23259 10074
rect 16724 9930 16788 9994
rect 17443 9930 17507 9994
rect 18162 9930 18226 9994
rect 18881 9930 18945 9994
rect 19600 9930 19664 9994
rect 20319 9930 20383 9994
rect 21038 9930 21102 9994
rect 21757 9930 21821 9994
rect 22476 9930 22540 9994
rect 23195 9930 23259 9994
rect 16724 9850 16788 9914
rect 17443 9850 17507 9914
rect 18162 9850 18226 9914
rect 18881 9850 18945 9914
rect 19600 9850 19664 9914
rect 20319 9850 20383 9914
rect 21038 9850 21102 9914
rect 21757 9850 21821 9914
rect 22476 9850 22540 9914
rect 23195 9850 23259 9914
rect 16138 9690 16202 9694
rect 16218 9690 16282 9694
rect 16138 9634 16182 9690
rect 16182 9634 16202 9690
rect 16218 9634 16238 9690
rect 16238 9634 16282 9690
rect 16138 9630 16202 9634
rect 16218 9630 16282 9634
rect 17264 9618 17328 9682
rect 924 9500 988 9504
rect 924 9444 928 9500
rect 928 9444 984 9500
rect 984 9444 988 9500
rect 924 9440 988 9444
rect 1004 9500 1068 9504
rect 1004 9444 1008 9500
rect 1008 9444 1064 9500
rect 1064 9444 1068 9500
rect 1004 9440 1068 9444
rect 1084 9500 1148 9504
rect 1084 9444 1088 9500
rect 1088 9444 1144 9500
rect 1144 9444 1148 9500
rect 1084 9440 1148 9444
rect 1164 9500 1228 9504
rect 1164 9444 1168 9500
rect 1168 9444 1224 9500
rect 1224 9444 1228 9500
rect 1164 9440 1228 9444
rect 1244 9500 1308 9504
rect 1244 9444 1248 9500
rect 1248 9444 1304 9500
rect 1304 9444 1308 9500
rect 1244 9440 1308 9444
rect 1324 9500 1388 9504
rect 1324 9444 1328 9500
rect 1328 9444 1384 9500
rect 1384 9444 1388 9500
rect 1324 9440 1388 9444
rect 1404 9500 1468 9504
rect 1404 9444 1408 9500
rect 1408 9444 1464 9500
rect 1464 9444 1468 9500
rect 1404 9440 1468 9444
rect 1484 9500 1548 9504
rect 1484 9444 1488 9500
rect 1488 9444 1544 9500
rect 1544 9444 1548 9500
rect 1484 9440 1548 9444
rect 1564 9500 1628 9504
rect 1564 9444 1568 9500
rect 1568 9444 1624 9500
rect 1624 9444 1628 9500
rect 1564 9440 1628 9444
rect 1644 9500 1708 9504
rect 1644 9444 1648 9500
rect 1648 9444 1704 9500
rect 1704 9444 1708 9500
rect 1644 9440 1708 9444
rect 1724 9500 1788 9504
rect 1724 9444 1728 9500
rect 1728 9444 1784 9500
rect 1784 9444 1788 9500
rect 1724 9440 1788 9444
rect 1804 9500 1868 9504
rect 1804 9444 1808 9500
rect 1808 9444 1864 9500
rect 1864 9444 1868 9500
rect 1804 9440 1868 9444
rect 1884 9500 1948 9504
rect 1884 9444 1888 9500
rect 1888 9444 1944 9500
rect 1944 9444 1948 9500
rect 1884 9440 1948 9444
rect 1964 9500 2028 9504
rect 1964 9444 1968 9500
rect 1968 9444 2024 9500
rect 2024 9444 2028 9500
rect 1964 9440 2028 9444
rect 2044 9500 2108 9504
rect 2044 9444 2048 9500
rect 2048 9444 2104 9500
rect 2104 9444 2108 9500
rect 2044 9440 2108 9444
rect 2124 9500 2188 9504
rect 2124 9444 2128 9500
rect 2128 9444 2184 9500
rect 2184 9444 2188 9500
rect 2124 9440 2188 9444
rect 2204 9500 2268 9504
rect 2204 9444 2208 9500
rect 2208 9444 2264 9500
rect 2264 9444 2268 9500
rect 2204 9440 2268 9444
rect 2284 9500 2348 9504
rect 2284 9444 2288 9500
rect 2288 9444 2344 9500
rect 2344 9444 2348 9500
rect 2284 9440 2348 9444
rect 2364 9500 2428 9504
rect 2364 9444 2368 9500
rect 2368 9444 2424 9500
rect 2424 9444 2428 9500
rect 2364 9440 2428 9444
rect 2444 9500 2508 9504
rect 2444 9444 2448 9500
rect 2448 9444 2504 9500
rect 2504 9444 2508 9500
rect 2444 9440 2508 9444
rect 46128 9500 46192 9504
rect 46128 9444 46132 9500
rect 46132 9444 46188 9500
rect 46188 9444 46192 9500
rect 46128 9440 46192 9444
rect 46208 9500 46272 9504
rect 46208 9444 46212 9500
rect 46212 9444 46268 9500
rect 46268 9444 46272 9500
rect 46208 9440 46272 9444
rect 46288 9500 46352 9504
rect 46288 9444 46292 9500
rect 46292 9444 46348 9500
rect 46348 9444 46352 9500
rect 46288 9440 46352 9444
rect 46368 9500 46432 9504
rect 46368 9444 46372 9500
rect 46372 9444 46428 9500
rect 46428 9444 46432 9500
rect 46368 9440 46432 9444
rect 46448 9500 46512 9504
rect 46448 9444 46452 9500
rect 46452 9444 46508 9500
rect 46508 9444 46512 9500
rect 46448 9440 46512 9444
rect 46528 9500 46592 9504
rect 46528 9444 46532 9500
rect 46532 9444 46588 9500
rect 46588 9444 46592 9500
rect 46528 9440 46592 9444
rect 46608 9500 46672 9504
rect 46608 9444 46612 9500
rect 46612 9444 46668 9500
rect 46668 9444 46672 9500
rect 46608 9440 46672 9444
rect 46688 9500 46752 9504
rect 46688 9444 46692 9500
rect 46692 9444 46748 9500
rect 46748 9444 46752 9500
rect 46688 9440 46752 9444
rect 46768 9500 46832 9504
rect 46768 9444 46772 9500
rect 46772 9444 46828 9500
rect 46828 9444 46832 9500
rect 46768 9440 46832 9444
rect 46848 9500 46912 9504
rect 46848 9444 46852 9500
rect 46852 9444 46908 9500
rect 46908 9444 46912 9500
rect 46848 9440 46912 9444
rect 46928 9500 46992 9504
rect 46928 9444 46932 9500
rect 46932 9444 46988 9500
rect 46988 9444 46992 9500
rect 46928 9440 46992 9444
rect 47008 9500 47072 9504
rect 47008 9444 47012 9500
rect 47012 9444 47068 9500
rect 47068 9444 47072 9500
rect 47008 9440 47072 9444
rect 47088 9500 47152 9504
rect 47088 9444 47092 9500
rect 47092 9444 47148 9500
rect 47148 9444 47152 9500
rect 47088 9440 47152 9444
rect 47168 9500 47232 9504
rect 47168 9444 47172 9500
rect 47172 9444 47228 9500
rect 47228 9444 47232 9500
rect 47168 9440 47232 9444
rect 47248 9500 47312 9504
rect 47248 9444 47252 9500
rect 47252 9444 47308 9500
rect 47308 9444 47312 9500
rect 47248 9440 47312 9444
rect 47328 9500 47392 9504
rect 47328 9444 47332 9500
rect 47332 9444 47388 9500
rect 47388 9444 47392 9500
rect 47328 9440 47392 9444
rect 47408 9500 47472 9504
rect 47408 9444 47412 9500
rect 47412 9444 47468 9500
rect 47468 9444 47472 9500
rect 47408 9440 47472 9444
rect 47488 9500 47552 9504
rect 47488 9444 47492 9500
rect 47492 9444 47548 9500
rect 47548 9444 47552 9500
rect 47488 9440 47552 9444
rect 47568 9500 47632 9504
rect 47568 9444 47572 9500
rect 47572 9444 47628 9500
rect 47628 9444 47632 9500
rect 47568 9440 47632 9444
rect 47648 9500 47712 9504
rect 47648 9444 47652 9500
rect 47652 9444 47708 9500
rect 47708 9444 47712 9500
rect 47648 9440 47712 9444
rect 3372 7620 3436 7624
rect 3372 7564 3376 7620
rect 3376 7564 3432 7620
rect 3432 7564 3436 7620
rect 3372 7560 3436 7564
rect 3452 7620 3516 7624
rect 3452 7564 3456 7620
rect 3456 7564 3512 7620
rect 3512 7564 3516 7620
rect 3452 7560 3516 7564
rect 3532 7620 3596 7624
rect 3532 7564 3536 7620
rect 3536 7564 3592 7620
rect 3592 7564 3596 7620
rect 3532 7560 3596 7564
rect 3612 7620 3676 7624
rect 3612 7564 3616 7620
rect 3616 7564 3672 7620
rect 3672 7564 3676 7620
rect 3612 7560 3676 7564
rect 3692 7620 3756 7624
rect 3692 7564 3696 7620
rect 3696 7564 3752 7620
rect 3752 7564 3756 7620
rect 3692 7560 3756 7564
rect 3772 7620 3836 7624
rect 3772 7564 3776 7620
rect 3776 7564 3832 7620
rect 3832 7564 3836 7620
rect 3772 7560 3836 7564
rect 3852 7620 3916 7624
rect 3852 7564 3856 7620
rect 3856 7564 3912 7620
rect 3912 7564 3916 7620
rect 3852 7560 3916 7564
rect 3932 7620 3996 7624
rect 3932 7564 3936 7620
rect 3936 7564 3992 7620
rect 3992 7564 3996 7620
rect 3932 7560 3996 7564
rect 4012 7620 4076 7624
rect 4012 7564 4016 7620
rect 4016 7564 4072 7620
rect 4072 7564 4076 7620
rect 4012 7560 4076 7564
rect 4092 7620 4156 7624
rect 4092 7564 4096 7620
rect 4096 7564 4152 7620
rect 4152 7564 4156 7620
rect 4092 7560 4156 7564
rect 4172 7620 4236 7624
rect 4172 7564 4176 7620
rect 4176 7564 4232 7620
rect 4232 7564 4236 7620
rect 4172 7560 4236 7564
rect 4252 7620 4316 7624
rect 4252 7564 4256 7620
rect 4256 7564 4312 7620
rect 4312 7564 4316 7620
rect 4252 7560 4316 7564
rect 4332 7620 4396 7624
rect 4332 7564 4336 7620
rect 4336 7564 4392 7620
rect 4392 7564 4396 7620
rect 4332 7560 4396 7564
rect 4412 7620 4476 7624
rect 4412 7564 4416 7620
rect 4416 7564 4472 7620
rect 4472 7564 4476 7620
rect 4412 7560 4476 7564
rect 4492 7620 4556 7624
rect 4492 7564 4496 7620
rect 4496 7564 4552 7620
rect 4552 7564 4556 7620
rect 4492 7560 4556 7564
rect 4572 7620 4636 7624
rect 4572 7564 4576 7620
rect 4576 7564 4632 7620
rect 4632 7564 4636 7620
rect 4572 7560 4636 7564
rect 4652 7620 4716 7624
rect 4652 7564 4656 7620
rect 4656 7564 4712 7620
rect 4712 7564 4716 7620
rect 4652 7560 4716 7564
rect 4732 7620 4796 7624
rect 4732 7564 4736 7620
rect 4736 7564 4792 7620
rect 4792 7564 4796 7620
rect 4732 7560 4796 7564
rect 4812 7620 4876 7624
rect 4812 7564 4816 7620
rect 4816 7564 4872 7620
rect 4872 7564 4876 7620
rect 4812 7560 4876 7564
rect 4892 7620 4956 7624
rect 4892 7564 4896 7620
rect 4896 7564 4952 7620
rect 4952 7564 4956 7620
rect 4892 7560 4956 7564
rect 43680 7620 43744 7624
rect 43680 7564 43684 7620
rect 43684 7564 43740 7620
rect 43740 7564 43744 7620
rect 43680 7560 43744 7564
rect 43760 7620 43824 7624
rect 43760 7564 43764 7620
rect 43764 7564 43820 7620
rect 43820 7564 43824 7620
rect 43760 7560 43824 7564
rect 43840 7620 43904 7624
rect 43840 7564 43844 7620
rect 43844 7564 43900 7620
rect 43900 7564 43904 7620
rect 43840 7560 43904 7564
rect 43920 7620 43984 7624
rect 43920 7564 43924 7620
rect 43924 7564 43980 7620
rect 43980 7564 43984 7620
rect 43920 7560 43984 7564
rect 44000 7620 44064 7624
rect 44000 7564 44004 7620
rect 44004 7564 44060 7620
rect 44060 7564 44064 7620
rect 44000 7560 44064 7564
rect 44080 7620 44144 7624
rect 44080 7564 44084 7620
rect 44084 7564 44140 7620
rect 44140 7564 44144 7620
rect 44080 7560 44144 7564
rect 44160 7620 44224 7624
rect 44160 7564 44164 7620
rect 44164 7564 44220 7620
rect 44220 7564 44224 7620
rect 44160 7560 44224 7564
rect 44240 7620 44304 7624
rect 44240 7564 44244 7620
rect 44244 7564 44300 7620
rect 44300 7564 44304 7620
rect 44240 7560 44304 7564
rect 44320 7620 44384 7624
rect 44320 7564 44324 7620
rect 44324 7564 44380 7620
rect 44380 7564 44384 7620
rect 44320 7560 44384 7564
rect 44400 7620 44464 7624
rect 44400 7564 44404 7620
rect 44404 7564 44460 7620
rect 44460 7564 44464 7620
rect 44400 7560 44464 7564
rect 44480 7620 44544 7624
rect 44480 7564 44484 7620
rect 44484 7564 44540 7620
rect 44540 7564 44544 7620
rect 44480 7560 44544 7564
rect 44560 7620 44624 7624
rect 44560 7564 44564 7620
rect 44564 7564 44620 7620
rect 44620 7564 44624 7620
rect 44560 7560 44624 7564
rect 44640 7620 44704 7624
rect 44640 7564 44644 7620
rect 44644 7564 44700 7620
rect 44700 7564 44704 7620
rect 44640 7560 44704 7564
rect 44720 7620 44784 7624
rect 44720 7564 44724 7620
rect 44724 7564 44780 7620
rect 44780 7564 44784 7620
rect 44720 7560 44784 7564
rect 44800 7620 44864 7624
rect 44800 7564 44804 7620
rect 44804 7564 44860 7620
rect 44860 7564 44864 7620
rect 44800 7560 44864 7564
rect 44880 7620 44944 7624
rect 44880 7564 44884 7620
rect 44884 7564 44940 7620
rect 44940 7564 44944 7620
rect 44880 7560 44944 7564
rect 44960 7620 45024 7624
rect 44960 7564 44964 7620
rect 44964 7564 45020 7620
rect 45020 7564 45024 7620
rect 44960 7560 45024 7564
rect 45040 7620 45104 7624
rect 45040 7564 45044 7620
rect 45044 7564 45100 7620
rect 45100 7564 45104 7620
rect 45040 7560 45104 7564
rect 45120 7620 45184 7624
rect 45120 7564 45124 7620
rect 45124 7564 45180 7620
rect 45180 7564 45184 7620
rect 45120 7560 45184 7564
rect 45200 7620 45264 7624
rect 45200 7564 45204 7620
rect 45204 7564 45260 7620
rect 45260 7564 45264 7620
rect 45200 7560 45264 7564
rect 924 5740 988 5744
rect 924 5684 928 5740
rect 928 5684 984 5740
rect 984 5684 988 5740
rect 924 5680 988 5684
rect 1004 5740 1068 5744
rect 1004 5684 1008 5740
rect 1008 5684 1064 5740
rect 1064 5684 1068 5740
rect 1004 5680 1068 5684
rect 1084 5740 1148 5744
rect 1084 5684 1088 5740
rect 1088 5684 1144 5740
rect 1144 5684 1148 5740
rect 1084 5680 1148 5684
rect 1164 5740 1228 5744
rect 1164 5684 1168 5740
rect 1168 5684 1224 5740
rect 1224 5684 1228 5740
rect 1164 5680 1228 5684
rect 1244 5740 1308 5744
rect 1244 5684 1248 5740
rect 1248 5684 1304 5740
rect 1304 5684 1308 5740
rect 1244 5680 1308 5684
rect 1324 5740 1388 5744
rect 1324 5684 1328 5740
rect 1328 5684 1384 5740
rect 1384 5684 1388 5740
rect 1324 5680 1388 5684
rect 1404 5740 1468 5744
rect 1404 5684 1408 5740
rect 1408 5684 1464 5740
rect 1464 5684 1468 5740
rect 1404 5680 1468 5684
rect 1484 5740 1548 5744
rect 1484 5684 1488 5740
rect 1488 5684 1544 5740
rect 1544 5684 1548 5740
rect 1484 5680 1548 5684
rect 1564 5740 1628 5744
rect 1564 5684 1568 5740
rect 1568 5684 1624 5740
rect 1624 5684 1628 5740
rect 1564 5680 1628 5684
rect 1644 5740 1708 5744
rect 1644 5684 1648 5740
rect 1648 5684 1704 5740
rect 1704 5684 1708 5740
rect 1644 5680 1708 5684
rect 1724 5740 1788 5744
rect 1724 5684 1728 5740
rect 1728 5684 1784 5740
rect 1784 5684 1788 5740
rect 1724 5680 1788 5684
rect 1804 5740 1868 5744
rect 1804 5684 1808 5740
rect 1808 5684 1864 5740
rect 1864 5684 1868 5740
rect 1804 5680 1868 5684
rect 1884 5740 1948 5744
rect 1884 5684 1888 5740
rect 1888 5684 1944 5740
rect 1944 5684 1948 5740
rect 1884 5680 1948 5684
rect 1964 5740 2028 5744
rect 1964 5684 1968 5740
rect 1968 5684 2024 5740
rect 2024 5684 2028 5740
rect 1964 5680 2028 5684
rect 2044 5740 2108 5744
rect 2044 5684 2048 5740
rect 2048 5684 2104 5740
rect 2104 5684 2108 5740
rect 2044 5680 2108 5684
rect 2124 5740 2188 5744
rect 2124 5684 2128 5740
rect 2128 5684 2184 5740
rect 2184 5684 2188 5740
rect 2124 5680 2188 5684
rect 2204 5740 2268 5744
rect 2204 5684 2208 5740
rect 2208 5684 2264 5740
rect 2264 5684 2268 5740
rect 2204 5680 2268 5684
rect 2284 5740 2348 5744
rect 2284 5684 2288 5740
rect 2288 5684 2344 5740
rect 2344 5684 2348 5740
rect 2284 5680 2348 5684
rect 2364 5740 2428 5744
rect 2364 5684 2368 5740
rect 2368 5684 2424 5740
rect 2424 5684 2428 5740
rect 2364 5680 2428 5684
rect 2444 5740 2508 5744
rect 2444 5684 2448 5740
rect 2448 5684 2504 5740
rect 2504 5684 2508 5740
rect 2444 5680 2508 5684
rect 46128 5740 46192 5744
rect 46128 5684 46132 5740
rect 46132 5684 46188 5740
rect 46188 5684 46192 5740
rect 46128 5680 46192 5684
rect 46208 5740 46272 5744
rect 46208 5684 46212 5740
rect 46212 5684 46268 5740
rect 46268 5684 46272 5740
rect 46208 5680 46272 5684
rect 46288 5740 46352 5744
rect 46288 5684 46292 5740
rect 46292 5684 46348 5740
rect 46348 5684 46352 5740
rect 46288 5680 46352 5684
rect 46368 5740 46432 5744
rect 46368 5684 46372 5740
rect 46372 5684 46428 5740
rect 46428 5684 46432 5740
rect 46368 5680 46432 5684
rect 46448 5740 46512 5744
rect 46448 5684 46452 5740
rect 46452 5684 46508 5740
rect 46508 5684 46512 5740
rect 46448 5680 46512 5684
rect 46528 5740 46592 5744
rect 46528 5684 46532 5740
rect 46532 5684 46588 5740
rect 46588 5684 46592 5740
rect 46528 5680 46592 5684
rect 46608 5740 46672 5744
rect 46608 5684 46612 5740
rect 46612 5684 46668 5740
rect 46668 5684 46672 5740
rect 46608 5680 46672 5684
rect 46688 5740 46752 5744
rect 46688 5684 46692 5740
rect 46692 5684 46748 5740
rect 46748 5684 46752 5740
rect 46688 5680 46752 5684
rect 46768 5740 46832 5744
rect 46768 5684 46772 5740
rect 46772 5684 46828 5740
rect 46828 5684 46832 5740
rect 46768 5680 46832 5684
rect 46848 5740 46912 5744
rect 46848 5684 46852 5740
rect 46852 5684 46908 5740
rect 46908 5684 46912 5740
rect 46848 5680 46912 5684
rect 46928 5740 46992 5744
rect 46928 5684 46932 5740
rect 46932 5684 46988 5740
rect 46988 5684 46992 5740
rect 46928 5680 46992 5684
rect 47008 5740 47072 5744
rect 47008 5684 47012 5740
rect 47012 5684 47068 5740
rect 47068 5684 47072 5740
rect 47008 5680 47072 5684
rect 47088 5740 47152 5744
rect 47088 5684 47092 5740
rect 47092 5684 47148 5740
rect 47148 5684 47152 5740
rect 47088 5680 47152 5684
rect 47168 5740 47232 5744
rect 47168 5684 47172 5740
rect 47172 5684 47228 5740
rect 47228 5684 47232 5740
rect 47168 5680 47232 5684
rect 47248 5740 47312 5744
rect 47248 5684 47252 5740
rect 47252 5684 47308 5740
rect 47308 5684 47312 5740
rect 47248 5680 47312 5684
rect 47328 5740 47392 5744
rect 47328 5684 47332 5740
rect 47332 5684 47388 5740
rect 47388 5684 47392 5740
rect 47328 5680 47392 5684
rect 47408 5740 47472 5744
rect 47408 5684 47412 5740
rect 47412 5684 47468 5740
rect 47468 5684 47472 5740
rect 47408 5680 47472 5684
rect 47488 5740 47552 5744
rect 47488 5684 47492 5740
rect 47492 5684 47548 5740
rect 47548 5684 47552 5740
rect 47488 5680 47552 5684
rect 47568 5740 47632 5744
rect 47568 5684 47572 5740
rect 47572 5684 47628 5740
rect 47628 5684 47632 5740
rect 47568 5680 47632 5684
rect 47648 5740 47712 5744
rect 47648 5684 47652 5740
rect 47652 5684 47708 5740
rect 47708 5684 47712 5740
rect 47648 5680 47712 5684
<< mimcap >>
rect 6899 41054 7299 41102
rect 6899 40750 6947 41054
rect 7251 40750 7299 41054
rect 6899 40702 7299 40750
rect 7618 41054 8018 41102
rect 7618 40750 7666 41054
rect 7970 40750 8018 41054
rect 7618 40702 8018 40750
rect 8337 41054 8737 41102
rect 8337 40750 8385 41054
rect 8689 40750 8737 41054
rect 8337 40702 8737 40750
rect 9056 41054 9456 41102
rect 9056 40750 9104 41054
rect 9408 40750 9456 41054
rect 9056 40702 9456 40750
rect 9775 41054 10175 41102
rect 9775 40750 9823 41054
rect 10127 40750 10175 41054
rect 9775 40702 10175 40750
rect 10494 41054 10894 41102
rect 10494 40750 10542 41054
rect 10846 40750 10894 41054
rect 10494 40702 10894 40750
rect 11213 41054 11613 41102
rect 11213 40750 11261 41054
rect 11565 40750 11613 41054
rect 11213 40702 11613 40750
rect 11932 41054 12332 41102
rect 11932 40750 11980 41054
rect 12284 40750 12332 41054
rect 11932 40702 12332 40750
rect 12651 41054 13051 41102
rect 12651 40750 12699 41054
rect 13003 40750 13051 41054
rect 12651 40702 13051 40750
rect 13370 41054 13770 41102
rect 13370 40750 13418 41054
rect 13722 40750 13770 41054
rect 13370 40702 13770 40750
rect 6899 40354 7299 40402
rect 6899 40050 6947 40354
rect 7251 40050 7299 40354
rect 6899 40002 7299 40050
rect 7618 40354 8018 40402
rect 7618 40050 7666 40354
rect 7970 40050 8018 40354
rect 7618 40002 8018 40050
rect 8337 40354 8737 40402
rect 8337 40050 8385 40354
rect 8689 40050 8737 40354
rect 8337 40002 8737 40050
rect 9056 40354 9456 40402
rect 9056 40050 9104 40354
rect 9408 40050 9456 40354
rect 9056 40002 9456 40050
rect 9775 40354 10175 40402
rect 9775 40050 9823 40354
rect 10127 40050 10175 40354
rect 9775 40002 10175 40050
rect 10494 40354 10894 40402
rect 10494 40050 10542 40354
rect 10846 40050 10894 40354
rect 10494 40002 10894 40050
rect 11213 40354 11613 40402
rect 11213 40050 11261 40354
rect 11565 40050 11613 40354
rect 11213 40002 11613 40050
rect 11932 40354 12332 40402
rect 11932 40050 11980 40354
rect 12284 40050 12332 40354
rect 11932 40002 12332 40050
rect 12651 40354 13051 40402
rect 12651 40050 12699 40354
rect 13003 40050 13051 40354
rect 12651 40002 13051 40050
rect 13370 40354 13770 40402
rect 13370 40050 13418 40354
rect 13722 40050 13770 40354
rect 13370 40002 13770 40050
rect 6017 37294 6417 37342
rect 6017 36990 6065 37294
rect 6369 36990 6417 37294
rect 6017 36942 6417 36990
rect 6736 37294 7136 37342
rect 6736 36990 6784 37294
rect 7088 36990 7136 37294
rect 6736 36942 7136 36990
rect 7455 37294 7855 37342
rect 7455 36990 7503 37294
rect 7807 36990 7855 37294
rect 7455 36942 7855 36990
rect 8174 37294 8574 37342
rect 8174 36990 8222 37294
rect 8526 36990 8574 37294
rect 8174 36942 8574 36990
rect 8893 37294 9293 37342
rect 8893 36990 8941 37294
rect 9245 36990 9293 37294
rect 8893 36942 9293 36990
rect 9612 37294 10012 37342
rect 9612 36990 9660 37294
rect 9964 36990 10012 37294
rect 9612 36942 10012 36990
rect 10331 37294 10731 37342
rect 10331 36990 10379 37294
rect 10683 36990 10731 37294
rect 10331 36942 10731 36990
rect 11050 37294 11450 37342
rect 11050 36990 11098 37294
rect 11402 36990 11450 37294
rect 11050 36942 11450 36990
rect 11769 37294 12169 37342
rect 11769 36990 11817 37294
rect 12121 36990 12169 37294
rect 11769 36942 12169 36990
rect 12488 37294 12888 37342
rect 12488 36990 12536 37294
rect 12840 36990 12888 37294
rect 12488 36942 12888 36990
rect 13465 37294 13865 37342
rect 13465 36990 13513 37294
rect 13817 36990 13865 37294
rect 13465 36942 13865 36990
rect 14184 37294 14584 37342
rect 14184 36990 14232 37294
rect 14536 36990 14584 37294
rect 14184 36942 14584 36990
rect 14903 37294 15303 37342
rect 14903 36990 14951 37294
rect 15255 36990 15303 37294
rect 14903 36942 15303 36990
rect 15622 37294 16022 37342
rect 15622 36990 15670 37294
rect 15974 36990 16022 37294
rect 15622 36942 16022 36990
rect 16341 37294 16741 37342
rect 16341 36990 16389 37294
rect 16693 36990 16741 37294
rect 16341 36942 16741 36990
rect 17060 37294 17460 37342
rect 17060 36990 17108 37294
rect 17412 36990 17460 37294
rect 17060 36942 17460 36990
rect 17779 37294 18179 37342
rect 17779 36990 17827 37294
rect 18131 36990 18179 37294
rect 17779 36942 18179 36990
rect 18498 37294 18898 37342
rect 18498 36990 18546 37294
rect 18850 36990 18898 37294
rect 18498 36942 18898 36990
rect 19217 37294 19617 37342
rect 19217 36990 19265 37294
rect 19569 36990 19617 37294
rect 19217 36942 19617 36990
rect 19936 37294 20336 37342
rect 19936 36990 19984 37294
rect 20288 36990 20336 37294
rect 19936 36942 20336 36990
rect 20913 37294 21313 37342
rect 20913 36990 20961 37294
rect 21265 36990 21313 37294
rect 20913 36942 21313 36990
rect 21632 37294 22032 37342
rect 21632 36990 21680 37294
rect 21984 36990 22032 37294
rect 21632 36942 22032 36990
rect 22351 37294 22751 37342
rect 22351 36990 22399 37294
rect 22703 36990 22751 37294
rect 22351 36942 22751 36990
rect 23070 37294 23470 37342
rect 23070 36990 23118 37294
rect 23422 36990 23470 37294
rect 23070 36942 23470 36990
rect 23789 37294 24189 37342
rect 23789 36990 23837 37294
rect 24141 36990 24189 37294
rect 23789 36942 24189 36990
rect 24508 37294 24908 37342
rect 24508 36990 24556 37294
rect 24860 36990 24908 37294
rect 24508 36942 24908 36990
rect 25227 37294 25627 37342
rect 25227 36990 25275 37294
rect 25579 36990 25627 37294
rect 25227 36942 25627 36990
rect 25946 37294 26346 37342
rect 25946 36990 25994 37294
rect 26298 36990 26346 37294
rect 25946 36942 26346 36990
rect 26665 37294 27065 37342
rect 26665 36990 26713 37294
rect 27017 36990 27065 37294
rect 26665 36942 27065 36990
rect 27384 37294 27784 37342
rect 27384 36990 27432 37294
rect 27736 36990 27784 37294
rect 27384 36942 27784 36990
rect 6017 36594 6417 36642
rect 6017 36290 6065 36594
rect 6369 36290 6417 36594
rect 6017 36242 6417 36290
rect 6736 36594 7136 36642
rect 6736 36290 6784 36594
rect 7088 36290 7136 36594
rect 6736 36242 7136 36290
rect 7455 36594 7855 36642
rect 7455 36290 7503 36594
rect 7807 36290 7855 36594
rect 7455 36242 7855 36290
rect 8174 36594 8574 36642
rect 8174 36290 8222 36594
rect 8526 36290 8574 36594
rect 8174 36242 8574 36290
rect 8893 36594 9293 36642
rect 8893 36290 8941 36594
rect 9245 36290 9293 36594
rect 8893 36242 9293 36290
rect 9612 36594 10012 36642
rect 9612 36290 9660 36594
rect 9964 36290 10012 36594
rect 9612 36242 10012 36290
rect 10331 36594 10731 36642
rect 10331 36290 10379 36594
rect 10683 36290 10731 36594
rect 10331 36242 10731 36290
rect 11050 36594 11450 36642
rect 11050 36290 11098 36594
rect 11402 36290 11450 36594
rect 11050 36242 11450 36290
rect 11769 36594 12169 36642
rect 11769 36290 11817 36594
rect 12121 36290 12169 36594
rect 11769 36242 12169 36290
rect 12488 36594 12888 36642
rect 12488 36290 12536 36594
rect 12840 36290 12888 36594
rect 12488 36242 12888 36290
rect 13465 36594 13865 36642
rect 13465 36290 13513 36594
rect 13817 36290 13865 36594
rect 13465 36242 13865 36290
rect 14184 36594 14584 36642
rect 14184 36290 14232 36594
rect 14536 36290 14584 36594
rect 14184 36242 14584 36290
rect 14903 36594 15303 36642
rect 14903 36290 14951 36594
rect 15255 36290 15303 36594
rect 14903 36242 15303 36290
rect 15622 36594 16022 36642
rect 15622 36290 15670 36594
rect 15974 36290 16022 36594
rect 15622 36242 16022 36290
rect 16341 36594 16741 36642
rect 16341 36290 16389 36594
rect 16693 36290 16741 36594
rect 16341 36242 16741 36290
rect 17060 36594 17460 36642
rect 17060 36290 17108 36594
rect 17412 36290 17460 36594
rect 17060 36242 17460 36290
rect 17779 36594 18179 36642
rect 17779 36290 17827 36594
rect 18131 36290 18179 36594
rect 17779 36242 18179 36290
rect 18498 36594 18898 36642
rect 18498 36290 18546 36594
rect 18850 36290 18898 36594
rect 18498 36242 18898 36290
rect 19217 36594 19617 36642
rect 19217 36290 19265 36594
rect 19569 36290 19617 36594
rect 19217 36242 19617 36290
rect 19936 36594 20336 36642
rect 19936 36290 19984 36594
rect 20288 36290 20336 36594
rect 19936 36242 20336 36290
rect 20913 36594 21313 36642
rect 20913 36290 20961 36594
rect 21265 36290 21313 36594
rect 20913 36242 21313 36290
rect 21632 36594 22032 36642
rect 21632 36290 21680 36594
rect 21984 36290 22032 36594
rect 21632 36242 22032 36290
rect 22351 36594 22751 36642
rect 22351 36290 22399 36594
rect 22703 36290 22751 36594
rect 22351 36242 22751 36290
rect 23070 36594 23470 36642
rect 23070 36290 23118 36594
rect 23422 36290 23470 36594
rect 23070 36242 23470 36290
rect 23789 36594 24189 36642
rect 23789 36290 23837 36594
rect 24141 36290 24189 36594
rect 23789 36242 24189 36290
rect 24508 36594 24908 36642
rect 24508 36290 24556 36594
rect 24860 36290 24908 36594
rect 24508 36242 24908 36290
rect 25227 36594 25627 36642
rect 25227 36290 25275 36594
rect 25579 36290 25627 36594
rect 25227 36242 25627 36290
rect 25946 36594 26346 36642
rect 25946 36290 25994 36594
rect 26298 36290 26346 36594
rect 25946 36242 26346 36290
rect 26665 36594 27065 36642
rect 26665 36290 26713 36594
rect 27017 36290 27065 36594
rect 26665 36242 27065 36290
rect 27384 36594 27784 36642
rect 27384 36290 27432 36594
rect 27736 36290 27784 36594
rect 27384 36242 27784 36290
rect 6703 33534 7103 33582
rect 6703 33230 6751 33534
rect 7055 33230 7103 33534
rect 6703 33182 7103 33230
rect 7422 33534 7822 33582
rect 7422 33230 7470 33534
rect 7774 33230 7822 33534
rect 7422 33182 7822 33230
rect 8141 33534 8541 33582
rect 8141 33230 8189 33534
rect 8493 33230 8541 33534
rect 8141 33182 8541 33230
rect 8860 33534 9260 33582
rect 8860 33230 8908 33534
rect 9212 33230 9260 33534
rect 8860 33182 9260 33230
rect 9579 33534 9979 33582
rect 9579 33230 9627 33534
rect 9931 33230 9979 33534
rect 9579 33182 9979 33230
rect 10298 33534 10698 33582
rect 10298 33230 10346 33534
rect 10650 33230 10698 33534
rect 10298 33182 10698 33230
rect 11017 33534 11417 33582
rect 11017 33230 11065 33534
rect 11369 33230 11417 33534
rect 11017 33182 11417 33230
rect 11736 33534 12136 33582
rect 11736 33230 11784 33534
rect 12088 33230 12136 33534
rect 11736 33182 12136 33230
rect 12455 33534 12855 33582
rect 12455 33230 12503 33534
rect 12807 33230 12855 33534
rect 12455 33182 12855 33230
rect 13174 33534 13574 33582
rect 13174 33230 13222 33534
rect 13526 33230 13574 33534
rect 13174 33182 13574 33230
rect 6703 32834 7103 32882
rect 6703 32530 6751 32834
rect 7055 32530 7103 32834
rect 6703 32482 7103 32530
rect 7422 32834 7822 32882
rect 7422 32530 7470 32834
rect 7774 32530 7822 32834
rect 7422 32482 7822 32530
rect 8141 32834 8541 32882
rect 8141 32530 8189 32834
rect 8493 32530 8541 32834
rect 8141 32482 8541 32530
rect 8860 32834 9260 32882
rect 8860 32530 8908 32834
rect 9212 32530 9260 32834
rect 8860 32482 9260 32530
rect 9579 32834 9979 32882
rect 9579 32530 9627 32834
rect 9931 32530 9979 32834
rect 9579 32482 9979 32530
rect 10298 32834 10698 32882
rect 10298 32530 10346 32834
rect 10650 32530 10698 32834
rect 10298 32482 10698 32530
rect 11017 32834 11417 32882
rect 11017 32530 11065 32834
rect 11369 32530 11417 32834
rect 11017 32482 11417 32530
rect 11736 32834 12136 32882
rect 11736 32530 11784 32834
rect 12088 32530 12136 32834
rect 11736 32482 12136 32530
rect 12455 32834 12855 32882
rect 12455 32530 12503 32834
rect 12807 32530 12855 32834
rect 12455 32482 12855 32530
rect 13174 32834 13574 32882
rect 13174 32530 13222 32834
rect 13526 32530 13574 32834
rect 13174 32482 13574 32530
rect 15523 26014 15923 26062
rect 15523 25710 15571 26014
rect 15875 25710 15923 26014
rect 15523 25662 15923 25710
rect 16242 26014 16642 26062
rect 16242 25710 16290 26014
rect 16594 25710 16642 26014
rect 16242 25662 16642 25710
rect 16961 26014 17361 26062
rect 16961 25710 17009 26014
rect 17313 25710 17361 26014
rect 16961 25662 17361 25710
rect 17680 26014 18080 26062
rect 17680 25710 17728 26014
rect 18032 25710 18080 26014
rect 17680 25662 18080 25710
rect 18399 26014 18799 26062
rect 18399 25710 18447 26014
rect 18751 25710 18799 26014
rect 18399 25662 18799 25710
rect 19118 26014 19518 26062
rect 19118 25710 19166 26014
rect 19470 25710 19518 26014
rect 19118 25662 19518 25710
rect 19837 26014 20237 26062
rect 19837 25710 19885 26014
rect 20189 25710 20237 26014
rect 19837 25662 20237 25710
rect 20556 26014 20956 26062
rect 20556 25710 20604 26014
rect 20908 25710 20956 26014
rect 20556 25662 20956 25710
rect 21275 26014 21675 26062
rect 21275 25710 21323 26014
rect 21627 25710 21675 26014
rect 21275 25662 21675 25710
rect 21994 26014 22394 26062
rect 21994 25710 22042 26014
rect 22346 25710 22394 26014
rect 21994 25662 22394 25710
rect 15523 25314 15923 25362
rect 15523 25010 15571 25314
rect 15875 25010 15923 25314
rect 15523 24962 15923 25010
rect 16242 25314 16642 25362
rect 16242 25010 16290 25314
rect 16594 25010 16642 25314
rect 16242 24962 16642 25010
rect 16961 25314 17361 25362
rect 16961 25010 17009 25314
rect 17313 25010 17361 25314
rect 16961 24962 17361 25010
rect 17680 25314 18080 25362
rect 17680 25010 17728 25314
rect 18032 25010 18080 25314
rect 17680 24962 18080 25010
rect 18399 25314 18799 25362
rect 18399 25010 18447 25314
rect 18751 25010 18799 25314
rect 18399 24962 18799 25010
rect 19118 25314 19518 25362
rect 19118 25010 19166 25314
rect 19470 25010 19518 25314
rect 19118 24962 19518 25010
rect 19837 25314 20237 25362
rect 19837 25010 19885 25314
rect 20189 25010 20237 25314
rect 19837 24962 20237 25010
rect 20556 25314 20956 25362
rect 20556 25010 20604 25314
rect 20908 25010 20956 25314
rect 20556 24962 20956 25010
rect 21275 25314 21675 25362
rect 21275 25010 21323 25314
rect 21627 25010 21675 25314
rect 21275 24962 21675 25010
rect 21994 25314 22394 25362
rect 21994 25010 22042 25314
rect 22346 25010 22394 25314
rect 21994 24962 22394 25010
rect 13661 22254 14061 22302
rect 13661 21950 13709 22254
rect 14013 21950 14061 22254
rect 13661 21902 14061 21950
rect 14380 22254 14780 22302
rect 14380 21950 14428 22254
rect 14732 21950 14780 22254
rect 14380 21902 14780 21950
rect 15099 22254 15499 22302
rect 15099 21950 15147 22254
rect 15451 21950 15499 22254
rect 15099 21902 15499 21950
rect 15818 22254 16218 22302
rect 15818 21950 15866 22254
rect 16170 21950 16218 22254
rect 15818 21902 16218 21950
rect 16537 22254 16937 22302
rect 16537 21950 16585 22254
rect 16889 21950 16937 22254
rect 16537 21902 16937 21950
rect 17256 22254 17656 22302
rect 17256 21950 17304 22254
rect 17608 21950 17656 22254
rect 17256 21902 17656 21950
rect 17975 22254 18375 22302
rect 17975 21950 18023 22254
rect 18327 21950 18375 22254
rect 17975 21902 18375 21950
rect 18694 22254 19094 22302
rect 18694 21950 18742 22254
rect 19046 21950 19094 22254
rect 18694 21902 19094 21950
rect 19413 22254 19813 22302
rect 19413 21950 19461 22254
rect 19765 21950 19813 22254
rect 19413 21902 19813 21950
rect 20132 22254 20532 22302
rect 20132 21950 20180 22254
rect 20484 21950 20532 22254
rect 20132 21902 20532 21950
rect 13661 21554 14061 21602
rect 13661 21250 13709 21554
rect 14013 21250 14061 21554
rect 13661 21202 14061 21250
rect 14380 21554 14780 21602
rect 14380 21250 14428 21554
rect 14732 21250 14780 21554
rect 14380 21202 14780 21250
rect 15099 21554 15499 21602
rect 15099 21250 15147 21554
rect 15451 21250 15499 21554
rect 15099 21202 15499 21250
rect 15818 21554 16218 21602
rect 15818 21250 15866 21554
rect 16170 21250 16218 21554
rect 15818 21202 16218 21250
rect 16537 21554 16937 21602
rect 16537 21250 16585 21554
rect 16889 21250 16937 21554
rect 16537 21202 16937 21250
rect 17256 21554 17656 21602
rect 17256 21250 17304 21554
rect 17608 21250 17656 21554
rect 17256 21202 17656 21250
rect 17975 21554 18375 21602
rect 17975 21250 18023 21554
rect 18327 21250 18375 21554
rect 17975 21202 18375 21250
rect 18694 21554 19094 21602
rect 18694 21250 18742 21554
rect 19046 21250 19094 21554
rect 18694 21202 19094 21250
rect 19413 21554 19813 21602
rect 19413 21250 19461 21554
rect 19765 21250 19813 21554
rect 19413 21202 19813 21250
rect 20132 21554 20532 21602
rect 20132 21250 20180 21554
rect 20484 21250 20532 21554
rect 20132 21202 20532 21250
rect 16209 18494 16609 18542
rect 16209 18190 16257 18494
rect 16561 18190 16609 18494
rect 16209 18142 16609 18190
rect 16928 18494 17328 18542
rect 16928 18190 16976 18494
rect 17280 18190 17328 18494
rect 16928 18142 17328 18190
rect 17647 18494 18047 18542
rect 17647 18190 17695 18494
rect 17999 18190 18047 18494
rect 17647 18142 18047 18190
rect 18366 18494 18766 18542
rect 18366 18190 18414 18494
rect 18718 18190 18766 18494
rect 18366 18142 18766 18190
rect 19085 18494 19485 18542
rect 19085 18190 19133 18494
rect 19437 18190 19485 18494
rect 19085 18142 19485 18190
rect 19804 18494 20204 18542
rect 19804 18190 19852 18494
rect 20156 18190 20204 18494
rect 19804 18142 20204 18190
rect 20523 18494 20923 18542
rect 20523 18190 20571 18494
rect 20875 18190 20923 18494
rect 20523 18142 20923 18190
rect 21242 18494 21642 18542
rect 21242 18190 21290 18494
rect 21594 18190 21642 18494
rect 21242 18142 21642 18190
rect 21961 18494 22361 18542
rect 21961 18190 22009 18494
rect 22313 18190 22361 18494
rect 21961 18142 22361 18190
rect 22680 18494 23080 18542
rect 22680 18190 22728 18494
rect 23032 18190 23080 18494
rect 22680 18142 23080 18190
rect 16209 17794 16609 17842
rect 16209 17490 16257 17794
rect 16561 17490 16609 17794
rect 16209 17442 16609 17490
rect 16928 17794 17328 17842
rect 16928 17490 16976 17794
rect 17280 17490 17328 17794
rect 16928 17442 17328 17490
rect 17647 17794 18047 17842
rect 17647 17490 17695 17794
rect 17999 17490 18047 17794
rect 17647 17442 18047 17490
rect 18366 17794 18766 17842
rect 18366 17490 18414 17794
rect 18718 17490 18766 17794
rect 18366 17442 18766 17490
rect 19085 17794 19485 17842
rect 19085 17490 19133 17794
rect 19437 17490 19485 17794
rect 19085 17442 19485 17490
rect 19804 17794 20204 17842
rect 19804 17490 19852 17794
rect 20156 17490 20204 17794
rect 19804 17442 20204 17490
rect 20523 17794 20923 17842
rect 20523 17490 20571 17794
rect 20875 17490 20923 17794
rect 20523 17442 20923 17490
rect 21242 17794 21642 17842
rect 21242 17490 21290 17794
rect 21594 17490 21642 17794
rect 21242 17442 21642 17490
rect 21961 17794 22361 17842
rect 21961 17490 22009 17794
rect 22313 17490 22361 17794
rect 21961 17442 22361 17490
rect 22680 17794 23080 17842
rect 22680 17490 22728 17794
rect 23032 17490 23080 17794
rect 22680 17442 23080 17490
rect 16209 14734 16609 14782
rect 16209 14430 16257 14734
rect 16561 14430 16609 14734
rect 16209 14382 16609 14430
rect 16928 14734 17328 14782
rect 16928 14430 16976 14734
rect 17280 14430 17328 14734
rect 16928 14382 17328 14430
rect 17647 14734 18047 14782
rect 17647 14430 17695 14734
rect 17999 14430 18047 14734
rect 17647 14382 18047 14430
rect 18366 14734 18766 14782
rect 18366 14430 18414 14734
rect 18718 14430 18766 14734
rect 18366 14382 18766 14430
rect 19085 14734 19485 14782
rect 19085 14430 19133 14734
rect 19437 14430 19485 14734
rect 19085 14382 19485 14430
rect 19804 14734 20204 14782
rect 19804 14430 19852 14734
rect 20156 14430 20204 14734
rect 19804 14382 20204 14430
rect 20523 14734 20923 14782
rect 20523 14430 20571 14734
rect 20875 14430 20923 14734
rect 20523 14382 20923 14430
rect 21242 14734 21642 14782
rect 21242 14430 21290 14734
rect 21594 14430 21642 14734
rect 21242 14382 21642 14430
rect 21961 14734 22361 14782
rect 21961 14430 22009 14734
rect 22313 14430 22361 14734
rect 21961 14382 22361 14430
rect 22680 14734 23080 14782
rect 22680 14430 22728 14734
rect 23032 14430 23080 14734
rect 22680 14382 23080 14430
rect 16209 14034 16609 14082
rect 16209 13730 16257 14034
rect 16561 13730 16609 14034
rect 16209 13682 16609 13730
rect 16928 14034 17328 14082
rect 16928 13730 16976 14034
rect 17280 13730 17328 14034
rect 16928 13682 17328 13730
rect 17647 14034 18047 14082
rect 17647 13730 17695 14034
rect 17999 13730 18047 14034
rect 17647 13682 18047 13730
rect 18366 14034 18766 14082
rect 18366 13730 18414 14034
rect 18718 13730 18766 14034
rect 18366 13682 18766 13730
rect 19085 14034 19485 14082
rect 19085 13730 19133 14034
rect 19437 13730 19485 14034
rect 19085 13682 19485 13730
rect 19804 14034 20204 14082
rect 19804 13730 19852 14034
rect 20156 13730 20204 14034
rect 19804 13682 20204 13730
rect 20523 14034 20923 14082
rect 20523 13730 20571 14034
rect 20875 13730 20923 14034
rect 20523 13682 20923 13730
rect 21242 14034 21642 14082
rect 21242 13730 21290 14034
rect 21594 13730 21642 14034
rect 21242 13682 21642 13730
rect 21961 14034 22361 14082
rect 21961 13730 22009 14034
rect 22313 13730 22361 14034
rect 21961 13682 22361 13730
rect 22680 14034 23080 14082
rect 22680 13730 22728 14034
rect 23032 13730 23080 14034
rect 22680 13682 23080 13730
rect 16209 10974 16609 11022
rect 16209 10670 16257 10974
rect 16561 10670 16609 10974
rect 16209 10622 16609 10670
rect 16928 10974 17328 11022
rect 16928 10670 16976 10974
rect 17280 10670 17328 10974
rect 16928 10622 17328 10670
rect 17647 10974 18047 11022
rect 17647 10670 17695 10974
rect 17999 10670 18047 10974
rect 17647 10622 18047 10670
rect 18366 10974 18766 11022
rect 18366 10670 18414 10974
rect 18718 10670 18766 10974
rect 18366 10622 18766 10670
rect 19085 10974 19485 11022
rect 19085 10670 19133 10974
rect 19437 10670 19485 10974
rect 19085 10622 19485 10670
rect 19804 10974 20204 11022
rect 19804 10670 19852 10974
rect 20156 10670 20204 10974
rect 19804 10622 20204 10670
rect 20523 10974 20923 11022
rect 20523 10670 20571 10974
rect 20875 10670 20923 10974
rect 20523 10622 20923 10670
rect 21242 10974 21642 11022
rect 21242 10670 21290 10974
rect 21594 10670 21642 10974
rect 21242 10622 21642 10670
rect 21961 10974 22361 11022
rect 21961 10670 22009 10974
rect 22313 10670 22361 10974
rect 21961 10622 22361 10670
rect 22680 10974 23080 11022
rect 22680 10670 22728 10974
rect 23032 10670 23080 10974
rect 22680 10622 23080 10670
rect 16209 10274 16609 10322
rect 16209 9970 16257 10274
rect 16561 9970 16609 10274
rect 16209 9922 16609 9970
rect 16928 10274 17328 10322
rect 16928 9970 16976 10274
rect 17280 9970 17328 10274
rect 16928 9922 17328 9970
rect 17647 10274 18047 10322
rect 17647 9970 17695 10274
rect 17999 9970 18047 10274
rect 17647 9922 18047 9970
rect 18366 10274 18766 10322
rect 18366 9970 18414 10274
rect 18718 9970 18766 10274
rect 18366 9922 18766 9970
rect 19085 10274 19485 10322
rect 19085 9970 19133 10274
rect 19437 9970 19485 10274
rect 19085 9922 19485 9970
rect 19804 10274 20204 10322
rect 19804 9970 19852 10274
rect 20156 9970 20204 10274
rect 19804 9922 20204 9970
rect 20523 10274 20923 10322
rect 20523 9970 20571 10274
rect 20875 9970 20923 10274
rect 20523 9922 20923 9970
rect 21242 10274 21642 10322
rect 21242 9970 21290 10274
rect 21594 9970 21642 10274
rect 21242 9922 21642 9970
rect 21961 10274 22361 10322
rect 21961 9970 22009 10274
rect 22313 9970 22361 10274
rect 21961 9922 22361 9970
rect 22680 10274 23080 10322
rect 22680 9970 22728 10274
rect 23032 9970 23080 10274
rect 22680 9922 23080 9970
<< mimcapcontact >>
rect 6947 40750 7251 41054
rect 7666 40750 7970 41054
rect 8385 40750 8689 41054
rect 9104 40750 9408 41054
rect 9823 40750 10127 41054
rect 10542 40750 10846 41054
rect 11261 40750 11565 41054
rect 11980 40750 12284 41054
rect 12699 40750 13003 41054
rect 13418 40750 13722 41054
rect 6947 40050 7251 40354
rect 7666 40050 7970 40354
rect 8385 40050 8689 40354
rect 9104 40050 9408 40354
rect 9823 40050 10127 40354
rect 10542 40050 10846 40354
rect 11261 40050 11565 40354
rect 11980 40050 12284 40354
rect 12699 40050 13003 40354
rect 13418 40050 13722 40354
rect 6065 36990 6369 37294
rect 6784 36990 7088 37294
rect 7503 36990 7807 37294
rect 8222 36990 8526 37294
rect 8941 36990 9245 37294
rect 9660 36990 9964 37294
rect 10379 36990 10683 37294
rect 11098 36990 11402 37294
rect 11817 36990 12121 37294
rect 12536 36990 12840 37294
rect 13513 36990 13817 37294
rect 14232 36990 14536 37294
rect 14951 36990 15255 37294
rect 15670 36990 15974 37294
rect 16389 36990 16693 37294
rect 17108 36990 17412 37294
rect 17827 36990 18131 37294
rect 18546 36990 18850 37294
rect 19265 36990 19569 37294
rect 19984 36990 20288 37294
rect 20961 36990 21265 37294
rect 21680 36990 21984 37294
rect 22399 36990 22703 37294
rect 23118 36990 23422 37294
rect 23837 36990 24141 37294
rect 24556 36990 24860 37294
rect 25275 36990 25579 37294
rect 25994 36990 26298 37294
rect 26713 36990 27017 37294
rect 27432 36990 27736 37294
rect 6065 36290 6369 36594
rect 6784 36290 7088 36594
rect 7503 36290 7807 36594
rect 8222 36290 8526 36594
rect 8941 36290 9245 36594
rect 9660 36290 9964 36594
rect 10379 36290 10683 36594
rect 11098 36290 11402 36594
rect 11817 36290 12121 36594
rect 12536 36290 12840 36594
rect 13513 36290 13817 36594
rect 14232 36290 14536 36594
rect 14951 36290 15255 36594
rect 15670 36290 15974 36594
rect 16389 36290 16693 36594
rect 17108 36290 17412 36594
rect 17827 36290 18131 36594
rect 18546 36290 18850 36594
rect 19265 36290 19569 36594
rect 19984 36290 20288 36594
rect 20961 36290 21265 36594
rect 21680 36290 21984 36594
rect 22399 36290 22703 36594
rect 23118 36290 23422 36594
rect 23837 36290 24141 36594
rect 24556 36290 24860 36594
rect 25275 36290 25579 36594
rect 25994 36290 26298 36594
rect 26713 36290 27017 36594
rect 27432 36290 27736 36594
rect 6751 33230 7055 33534
rect 7470 33230 7774 33534
rect 8189 33230 8493 33534
rect 8908 33230 9212 33534
rect 9627 33230 9931 33534
rect 10346 33230 10650 33534
rect 11065 33230 11369 33534
rect 11784 33230 12088 33534
rect 12503 33230 12807 33534
rect 13222 33230 13526 33534
rect 6751 32530 7055 32834
rect 7470 32530 7774 32834
rect 8189 32530 8493 32834
rect 8908 32530 9212 32834
rect 9627 32530 9931 32834
rect 10346 32530 10650 32834
rect 11065 32530 11369 32834
rect 11784 32530 12088 32834
rect 12503 32530 12807 32834
rect 13222 32530 13526 32834
rect 15571 25710 15875 26014
rect 16290 25710 16594 26014
rect 17009 25710 17313 26014
rect 17728 25710 18032 26014
rect 18447 25710 18751 26014
rect 19166 25710 19470 26014
rect 19885 25710 20189 26014
rect 20604 25710 20908 26014
rect 21323 25710 21627 26014
rect 22042 25710 22346 26014
rect 15571 25010 15875 25314
rect 16290 25010 16594 25314
rect 17009 25010 17313 25314
rect 17728 25010 18032 25314
rect 18447 25010 18751 25314
rect 19166 25010 19470 25314
rect 19885 25010 20189 25314
rect 20604 25010 20908 25314
rect 21323 25010 21627 25314
rect 22042 25010 22346 25314
rect 13709 21950 14013 22254
rect 14428 21950 14732 22254
rect 15147 21950 15451 22254
rect 15866 21950 16170 22254
rect 16585 21950 16889 22254
rect 17304 21950 17608 22254
rect 18023 21950 18327 22254
rect 18742 21950 19046 22254
rect 19461 21950 19765 22254
rect 20180 21950 20484 22254
rect 13709 21250 14013 21554
rect 14428 21250 14732 21554
rect 15147 21250 15451 21554
rect 15866 21250 16170 21554
rect 16585 21250 16889 21554
rect 17304 21250 17608 21554
rect 18023 21250 18327 21554
rect 18742 21250 19046 21554
rect 19461 21250 19765 21554
rect 20180 21250 20484 21554
rect 16257 18190 16561 18494
rect 16976 18190 17280 18494
rect 17695 18190 17999 18494
rect 18414 18190 18718 18494
rect 19133 18190 19437 18494
rect 19852 18190 20156 18494
rect 20571 18190 20875 18494
rect 21290 18190 21594 18494
rect 22009 18190 22313 18494
rect 22728 18190 23032 18494
rect 16257 17490 16561 17794
rect 16976 17490 17280 17794
rect 17695 17490 17999 17794
rect 18414 17490 18718 17794
rect 19133 17490 19437 17794
rect 19852 17490 20156 17794
rect 20571 17490 20875 17794
rect 21290 17490 21594 17794
rect 22009 17490 22313 17794
rect 22728 17490 23032 17794
rect 16257 14430 16561 14734
rect 16976 14430 17280 14734
rect 17695 14430 17999 14734
rect 18414 14430 18718 14734
rect 19133 14430 19437 14734
rect 19852 14430 20156 14734
rect 20571 14430 20875 14734
rect 21290 14430 21594 14734
rect 22009 14430 22313 14734
rect 22728 14430 23032 14734
rect 16257 13730 16561 14034
rect 16976 13730 17280 14034
rect 17695 13730 17999 14034
rect 18414 13730 18718 14034
rect 19133 13730 19437 14034
rect 19852 13730 20156 14034
rect 20571 13730 20875 14034
rect 21290 13730 21594 14034
rect 22009 13730 22313 14034
rect 22728 13730 23032 14034
rect 16257 10670 16561 10974
rect 16976 10670 17280 10974
rect 17695 10670 17999 10974
rect 18414 10670 18718 10974
rect 19133 10670 19437 10974
rect 19852 10670 20156 10974
rect 20571 10670 20875 10974
rect 21290 10670 21594 10974
rect 22009 10670 22313 10974
rect 22728 10670 23032 10974
rect 16257 9970 16561 10274
rect 16976 9970 17280 10274
rect 17695 9970 17999 10274
rect 18414 9970 18718 10274
rect 19133 9970 19437 10274
rect 19852 9970 20156 10274
rect 20571 9970 20875 10274
rect 21290 9970 21594 10274
rect 22009 9970 22313 10274
rect 22728 9970 23032 10274
<< metal4 >>
rect 900 46270 2532 47192
rect 900 44754 958 46270
rect 2474 44754 2532 46270
rect 900 39584 2532 44754
rect 900 39520 924 39584
rect 988 39520 1004 39584
rect 1068 39520 1084 39584
rect 1148 39520 1164 39584
rect 1228 39520 1244 39584
rect 1308 39520 1324 39584
rect 1388 39520 1404 39584
rect 1468 39520 1484 39584
rect 1548 39520 1564 39584
rect 1628 39520 1644 39584
rect 1708 39520 1724 39584
rect 1788 39520 1804 39584
rect 1868 39520 1884 39584
rect 1948 39520 1964 39584
rect 2028 39520 2044 39584
rect 2108 39520 2124 39584
rect 2188 39520 2204 39584
rect 2268 39520 2284 39584
rect 2348 39520 2364 39584
rect 2428 39520 2444 39584
rect 2508 39520 2532 39584
rect 900 35824 2532 39520
rect 900 35760 924 35824
rect 988 35760 1004 35824
rect 1068 35760 1084 35824
rect 1148 35760 1164 35824
rect 1228 35760 1244 35824
rect 1308 35760 1324 35824
rect 1388 35760 1404 35824
rect 1468 35760 1484 35824
rect 1548 35760 1564 35824
rect 1628 35760 1644 35824
rect 1708 35760 1724 35824
rect 1788 35760 1804 35824
rect 1868 35760 1884 35824
rect 1948 35760 1964 35824
rect 2028 35760 2044 35824
rect 2108 35760 2124 35824
rect 2188 35760 2204 35824
rect 2268 35760 2284 35824
rect 2348 35760 2364 35824
rect 2428 35760 2444 35824
rect 2508 35760 2532 35824
rect 900 32064 2532 35760
rect 900 32000 924 32064
rect 988 32000 1004 32064
rect 1068 32000 1084 32064
rect 1148 32000 1164 32064
rect 1228 32000 1244 32064
rect 1308 32000 1324 32064
rect 1388 32000 1404 32064
rect 1468 32000 1484 32064
rect 1548 32000 1564 32064
rect 1628 32000 1644 32064
rect 1708 32000 1724 32064
rect 1788 32000 1804 32064
rect 1868 32000 1884 32064
rect 1948 32000 1964 32064
rect 2028 32000 2044 32064
rect 2108 32000 2124 32064
rect 2188 32000 2204 32064
rect 2268 32000 2284 32064
rect 2348 32000 2364 32064
rect 2428 32000 2444 32064
rect 2508 32000 2532 32064
rect 900 28304 2532 32000
rect 900 28240 924 28304
rect 988 28240 1004 28304
rect 1068 28240 1084 28304
rect 1148 28240 1164 28304
rect 1228 28240 1244 28304
rect 1308 28240 1324 28304
rect 1388 28240 1404 28304
rect 1468 28240 1484 28304
rect 1548 28240 1564 28304
rect 1628 28240 1644 28304
rect 1708 28240 1724 28304
rect 1788 28240 1804 28304
rect 1868 28240 1884 28304
rect 1948 28240 1964 28304
rect 2028 28240 2044 28304
rect 2108 28240 2124 28304
rect 2188 28240 2204 28304
rect 2268 28240 2284 28304
rect 2348 28240 2364 28304
rect 2428 28240 2444 28304
rect 2508 28240 2532 28304
rect 900 24544 2532 28240
rect 900 24480 924 24544
rect 988 24480 1004 24544
rect 1068 24480 1084 24544
rect 1148 24480 1164 24544
rect 1228 24480 1244 24544
rect 1308 24480 1324 24544
rect 1388 24480 1404 24544
rect 1468 24480 1484 24544
rect 1548 24480 1564 24544
rect 1628 24480 1644 24544
rect 1708 24480 1724 24544
rect 1788 24480 1804 24544
rect 1868 24480 1884 24544
rect 1948 24480 1964 24544
rect 2028 24480 2044 24544
rect 2108 24480 2124 24544
rect 2188 24480 2204 24544
rect 2268 24480 2284 24544
rect 2348 24480 2364 24544
rect 2428 24480 2444 24544
rect 2508 24480 2532 24544
rect 900 20784 2532 24480
rect 900 20720 924 20784
rect 988 20720 1004 20784
rect 1068 20720 1084 20784
rect 1148 20720 1164 20784
rect 1228 20720 1244 20784
rect 1308 20720 1324 20784
rect 1388 20720 1404 20784
rect 1468 20720 1484 20784
rect 1548 20720 1564 20784
rect 1628 20720 1644 20784
rect 1708 20720 1724 20784
rect 1788 20720 1804 20784
rect 1868 20720 1884 20784
rect 1948 20720 1964 20784
rect 2028 20720 2044 20784
rect 2108 20720 2124 20784
rect 2188 20720 2204 20784
rect 2268 20720 2284 20784
rect 2348 20720 2364 20784
rect 2428 20720 2444 20784
rect 2508 20720 2532 20784
rect 900 17024 2532 20720
rect 900 16960 924 17024
rect 988 16960 1004 17024
rect 1068 16960 1084 17024
rect 1148 16960 1164 17024
rect 1228 16960 1244 17024
rect 1308 16960 1324 17024
rect 1388 16960 1404 17024
rect 1468 16960 1484 17024
rect 1548 16960 1564 17024
rect 1628 16960 1644 17024
rect 1708 16960 1724 17024
rect 1788 16960 1804 17024
rect 1868 16960 1884 17024
rect 1948 16960 1964 17024
rect 2028 16960 2044 17024
rect 2108 16960 2124 17024
rect 2188 16960 2204 17024
rect 2268 16960 2284 17024
rect 2348 16960 2364 17024
rect 2428 16960 2444 17024
rect 2508 16960 2532 17024
rect 900 13264 2532 16960
rect 900 13200 924 13264
rect 988 13200 1004 13264
rect 1068 13200 1084 13264
rect 1148 13200 1164 13264
rect 1228 13200 1244 13264
rect 1308 13200 1324 13264
rect 1388 13200 1404 13264
rect 1468 13200 1484 13264
rect 1548 13200 1564 13264
rect 1628 13200 1644 13264
rect 1708 13200 1724 13264
rect 1788 13200 1804 13264
rect 1868 13200 1884 13264
rect 1948 13200 1964 13264
rect 2028 13200 2044 13264
rect 2108 13200 2124 13264
rect 2188 13200 2204 13264
rect 2268 13200 2284 13264
rect 2348 13200 2364 13264
rect 2428 13200 2444 13264
rect 2508 13200 2532 13264
rect 900 9504 2532 13200
rect 900 9440 924 9504
rect 988 9440 1004 9504
rect 1068 9440 1084 9504
rect 1148 9440 1164 9504
rect 1228 9440 1244 9504
rect 1308 9440 1324 9504
rect 1388 9440 1404 9504
rect 1468 9440 1484 9504
rect 1548 9440 1564 9504
rect 1628 9440 1644 9504
rect 1708 9440 1724 9504
rect 1788 9440 1804 9504
rect 1868 9440 1884 9504
rect 1948 9440 1964 9504
rect 2028 9440 2044 9504
rect 2108 9440 2124 9504
rect 2188 9440 2204 9504
rect 2268 9440 2284 9504
rect 2348 9440 2364 9504
rect 2428 9440 2444 9504
rect 2508 9440 2532 9504
rect 900 5744 2532 9440
rect 900 5680 924 5744
rect 988 5680 1004 5744
rect 1068 5680 1084 5744
rect 1148 5680 1164 5744
rect 1228 5680 1244 5744
rect 1308 5680 1324 5744
rect 1388 5680 1404 5744
rect 1468 5680 1484 5744
rect 1548 5680 1564 5744
rect 1628 5680 1644 5744
rect 1708 5680 1724 5744
rect 1788 5680 1804 5744
rect 1868 5680 1884 5744
rect 1948 5680 1964 5744
rect 2028 5680 2044 5744
rect 2108 5680 2124 5744
rect 2188 5680 2204 5744
rect 2268 5680 2284 5744
rect 2348 5680 2364 5744
rect 2428 5680 2444 5744
rect 2508 5680 2532 5744
rect 900 2390 2532 5680
rect 900 874 958 2390
rect 2474 874 2532 2390
rect 900 0 2532 874
rect 3348 43822 4980 47192
rect 3348 42306 3406 43822
rect 4922 42306 4980 43822
rect 3348 41464 4980 42306
rect 3348 41400 3372 41464
rect 3436 41400 3452 41464
rect 3516 41400 3532 41464
rect 3596 41400 3612 41464
rect 3676 41400 3692 41464
rect 3756 41400 3772 41464
rect 3836 41400 3852 41464
rect 3916 41400 3932 41464
rect 3996 41400 4012 41464
rect 4076 41400 4092 41464
rect 4156 41400 4172 41464
rect 4236 41400 4252 41464
rect 4316 41400 4332 41464
rect 4396 41400 4412 41464
rect 4476 41400 4492 41464
rect 4556 41400 4572 41464
rect 4636 41400 4652 41464
rect 4716 41400 4732 41464
rect 4796 41400 4812 41464
rect 4876 41400 4892 41464
rect 4956 41400 4980 41464
rect 43656 43822 45288 47192
rect 43656 42306 43714 43822
rect 45230 42306 45288 43822
rect 43656 41464 45288 42306
rect 3348 37704 4980 41400
rect 12433 41402 12499 41403
rect 12433 41338 12434 41402
rect 12498 41338 12499 41402
rect 12433 41337 12499 41338
rect 43656 41400 43680 41464
rect 43744 41400 43760 41464
rect 43824 41400 43840 41464
rect 43904 41400 43920 41464
rect 43984 41400 44000 41464
rect 44064 41400 44080 41464
rect 44144 41400 44160 41464
rect 44224 41400 44240 41464
rect 44304 41400 44320 41464
rect 44384 41400 44400 41464
rect 44464 41400 44480 41464
rect 44544 41400 44560 41464
rect 44624 41400 44640 41464
rect 44704 41400 44720 41464
rect 44784 41400 44800 41464
rect 44864 41400 44880 41464
rect 44944 41400 44960 41464
rect 45024 41400 45040 41464
rect 45104 41400 45120 41464
rect 45184 41400 45200 41464
rect 45264 41400 45288 41464
rect 12436 41190 12496 41337
rect 7398 41174 7494 41190
rect 7398 41110 7414 41174
rect 7478 41110 7494 41174
rect 7398 41094 7494 41110
rect 6938 41063 7258 41082
rect 6938 41054 7260 41063
rect 6938 40750 6947 41054
rect 7251 40750 7260 41054
rect 6938 40741 7260 40750
rect 7398 41030 7414 41094
rect 7478 41030 7494 41094
rect 8117 41174 8213 41190
rect 8117 41110 8133 41174
rect 8197 41110 8213 41174
rect 8117 41094 8213 41110
rect 7658 41063 7978 41082
rect 7398 41014 7494 41030
rect 7398 40950 7414 41014
rect 7478 40950 7494 41014
rect 7398 40934 7494 40950
rect 7398 40870 7414 40934
rect 7478 40870 7494 40934
rect 7398 40854 7494 40870
rect 7398 40790 7414 40854
rect 7478 40790 7494 40854
rect 7398 40774 7494 40790
rect 6938 40363 7258 40741
rect 7398 40710 7414 40774
rect 7478 40710 7494 40774
rect 7657 41054 7979 41063
rect 7657 40750 7666 41054
rect 7970 40750 7979 41054
rect 7657 40741 7979 40750
rect 8117 41030 8133 41094
rect 8197 41030 8213 41094
rect 8836 41174 8932 41190
rect 8836 41110 8852 41174
rect 8916 41110 8932 41174
rect 8836 41094 8932 41110
rect 8378 41063 8698 41082
rect 8117 41014 8213 41030
rect 8117 40950 8133 41014
rect 8197 40950 8213 41014
rect 8117 40934 8213 40950
rect 8117 40870 8133 40934
rect 8197 40870 8213 40934
rect 8117 40854 8213 40870
rect 8117 40790 8133 40854
rect 8197 40790 8213 40854
rect 8117 40774 8213 40790
rect 7398 40694 7494 40710
rect 7398 40630 7414 40694
rect 7478 40630 7494 40694
rect 7398 40614 7494 40630
rect 7398 40474 7494 40490
rect 7398 40410 7414 40474
rect 7478 40410 7494 40474
rect 7398 40394 7494 40410
rect 6938 40354 7260 40363
rect 6938 40050 6947 40354
rect 7251 40050 7260 40354
rect 6938 40041 7260 40050
rect 7398 40330 7414 40394
rect 7478 40330 7494 40394
rect 7658 40363 7978 40741
rect 8117 40710 8133 40774
rect 8197 40710 8213 40774
rect 8376 41054 8698 41063
rect 8376 40750 8385 41054
rect 8689 40750 8698 41054
rect 8376 40741 8698 40750
rect 8117 40694 8213 40710
rect 8117 40630 8133 40694
rect 8197 40630 8213 40694
rect 8117 40614 8213 40630
rect 8117 40474 8213 40490
rect 8117 40410 8133 40474
rect 8197 40410 8213 40474
rect 8117 40394 8213 40410
rect 7398 40314 7494 40330
rect 7398 40250 7414 40314
rect 7478 40250 7494 40314
rect 7398 40234 7494 40250
rect 7398 40170 7414 40234
rect 7478 40170 7494 40234
rect 7398 40154 7494 40170
rect 7398 40090 7414 40154
rect 7478 40090 7494 40154
rect 7398 40074 7494 40090
rect 6938 39802 7258 40041
rect 7398 40010 7414 40074
rect 7478 40010 7494 40074
rect 7657 40354 7979 40363
rect 7657 40050 7666 40354
rect 7970 40050 7979 40354
rect 7657 40041 7979 40050
rect 8117 40330 8133 40394
rect 8197 40330 8213 40394
rect 8378 40363 8698 40741
rect 8836 41030 8852 41094
rect 8916 41030 8932 41094
rect 9555 41174 9651 41190
rect 9555 41110 9571 41174
rect 9635 41110 9651 41174
rect 9555 41094 9651 41110
rect 9098 41063 9418 41082
rect 8836 41014 8932 41030
rect 8836 40950 8852 41014
rect 8916 40950 8932 41014
rect 8836 40934 8932 40950
rect 8836 40870 8852 40934
rect 8916 40870 8932 40934
rect 8836 40854 8932 40870
rect 8836 40790 8852 40854
rect 8916 40790 8932 40854
rect 8836 40774 8932 40790
rect 8836 40710 8852 40774
rect 8916 40710 8932 40774
rect 9095 41054 9418 41063
rect 9095 40750 9104 41054
rect 9408 40750 9418 41054
rect 9095 40741 9418 40750
rect 8836 40694 8932 40710
rect 8836 40630 8852 40694
rect 8916 40630 8932 40694
rect 8836 40614 8932 40630
rect 8117 40314 8213 40330
rect 8117 40250 8133 40314
rect 8197 40250 8213 40314
rect 8117 40234 8213 40250
rect 8117 40170 8133 40234
rect 8197 40170 8213 40234
rect 8117 40154 8213 40170
rect 8117 40090 8133 40154
rect 8197 40090 8213 40154
rect 8117 40074 8213 40090
rect 7398 39994 7494 40010
rect 7398 39930 7414 39994
rect 7478 39930 7494 39994
rect 7398 39914 7494 39930
rect 7658 39802 7978 40041
rect 8117 40010 8133 40074
rect 8197 40010 8213 40074
rect 8376 40354 8698 40363
rect 8376 40050 8385 40354
rect 8689 40050 8698 40354
rect 8376 40041 8698 40050
rect 8117 39994 8213 40010
rect 8117 39930 8133 39994
rect 8197 39930 8213 39994
rect 8117 39914 8213 39930
rect 8378 39802 8698 40041
rect 8836 40474 8932 40490
rect 8836 40410 8852 40474
rect 8916 40410 8932 40474
rect 8836 40394 8932 40410
rect 8836 40330 8852 40394
rect 8916 40330 8932 40394
rect 9098 40363 9418 40741
rect 9555 41030 9571 41094
rect 9635 41030 9651 41094
rect 10274 41174 10370 41190
rect 10274 41110 10290 41174
rect 10354 41110 10370 41174
rect 10274 41094 10370 41110
rect 9818 41063 10138 41082
rect 9555 41014 9651 41030
rect 9555 40950 9571 41014
rect 9635 40950 9651 41014
rect 9555 40934 9651 40950
rect 9555 40870 9571 40934
rect 9635 40870 9651 40934
rect 9555 40854 9651 40870
rect 9555 40790 9571 40854
rect 9635 40790 9651 40854
rect 9555 40774 9651 40790
rect 9555 40710 9571 40774
rect 9635 40710 9651 40774
rect 9814 41054 10138 41063
rect 9814 40750 9823 41054
rect 10127 40750 10138 41054
rect 9814 40741 10138 40750
rect 9555 40694 9651 40710
rect 9555 40630 9571 40694
rect 9635 40630 9651 40694
rect 9555 40614 9651 40630
rect 8836 40314 8932 40330
rect 8836 40250 8852 40314
rect 8916 40250 8932 40314
rect 8836 40234 8932 40250
rect 8836 40170 8852 40234
rect 8916 40170 8932 40234
rect 8836 40154 8932 40170
rect 8836 40090 8852 40154
rect 8916 40090 8932 40154
rect 8836 40074 8932 40090
rect 8836 40010 8852 40074
rect 8916 40010 8932 40074
rect 9095 40354 9418 40363
rect 9095 40050 9104 40354
rect 9408 40050 9418 40354
rect 9095 40041 9418 40050
rect 8836 39994 8932 40010
rect 8836 39930 8852 39994
rect 8916 39930 8932 39994
rect 8836 39914 8932 39930
rect 9098 39802 9418 40041
rect 9555 40474 9651 40490
rect 9555 40410 9571 40474
rect 9635 40410 9651 40474
rect 9555 40394 9651 40410
rect 9555 40330 9571 40394
rect 9635 40330 9651 40394
rect 9818 40363 10138 40741
rect 10274 41030 10290 41094
rect 10354 41030 10370 41094
rect 10993 41174 11089 41190
rect 10993 41110 11009 41174
rect 11073 41110 11089 41174
rect 10993 41094 11089 41110
rect 10538 41063 10858 41082
rect 10274 41014 10370 41030
rect 10274 40950 10290 41014
rect 10354 40950 10370 41014
rect 10274 40934 10370 40950
rect 10274 40870 10290 40934
rect 10354 40870 10370 40934
rect 10274 40854 10370 40870
rect 10274 40790 10290 40854
rect 10354 40790 10370 40854
rect 10274 40774 10370 40790
rect 10274 40710 10290 40774
rect 10354 40710 10370 40774
rect 10533 41054 10858 41063
rect 10533 40750 10542 41054
rect 10846 40750 10858 41054
rect 10533 40741 10858 40750
rect 10274 40694 10370 40710
rect 10274 40630 10290 40694
rect 10354 40630 10370 40694
rect 10274 40614 10370 40630
rect 9555 40314 9651 40330
rect 9555 40250 9571 40314
rect 9635 40250 9651 40314
rect 9555 40234 9651 40250
rect 9555 40170 9571 40234
rect 9635 40170 9651 40234
rect 9555 40154 9651 40170
rect 9555 40090 9571 40154
rect 9635 40090 9651 40154
rect 9555 40074 9651 40090
rect 9555 40010 9571 40074
rect 9635 40010 9651 40074
rect 9814 40354 10138 40363
rect 9814 40050 9823 40354
rect 10127 40050 10138 40354
rect 9814 40041 10138 40050
rect 9555 39994 9651 40010
rect 9555 39930 9571 39994
rect 9635 39930 9651 39994
rect 9555 39914 9651 39930
rect 9818 39802 10138 40041
rect 10274 40474 10370 40490
rect 10274 40410 10290 40474
rect 10354 40410 10370 40474
rect 10274 40394 10370 40410
rect 10274 40330 10290 40394
rect 10354 40330 10370 40394
rect 10538 40363 10858 40741
rect 10993 41030 11009 41094
rect 11073 41030 11089 41094
rect 11712 41174 11808 41190
rect 11712 41110 11728 41174
rect 11792 41110 11808 41174
rect 11712 41094 11808 41110
rect 11258 41063 11578 41082
rect 10993 41014 11089 41030
rect 10993 40950 11009 41014
rect 11073 40950 11089 41014
rect 10993 40934 11089 40950
rect 10993 40870 11009 40934
rect 11073 40870 11089 40934
rect 10993 40854 11089 40870
rect 10993 40790 11009 40854
rect 11073 40790 11089 40854
rect 10993 40774 11089 40790
rect 10993 40710 11009 40774
rect 11073 40710 11089 40774
rect 11252 41054 11578 41063
rect 11252 40750 11261 41054
rect 11565 40750 11578 41054
rect 11252 40741 11578 40750
rect 10993 40694 11089 40710
rect 10993 40630 11009 40694
rect 11073 40630 11089 40694
rect 10993 40614 11089 40630
rect 10274 40314 10370 40330
rect 10274 40250 10290 40314
rect 10354 40250 10370 40314
rect 10274 40234 10370 40250
rect 10274 40170 10290 40234
rect 10354 40170 10370 40234
rect 10274 40154 10370 40170
rect 10274 40090 10290 40154
rect 10354 40090 10370 40154
rect 10274 40074 10370 40090
rect 10274 40010 10290 40074
rect 10354 40010 10370 40074
rect 10533 40354 10858 40363
rect 10533 40050 10542 40354
rect 10846 40050 10858 40354
rect 10533 40041 10858 40050
rect 10274 39994 10370 40010
rect 10274 39930 10290 39994
rect 10354 39930 10370 39994
rect 10274 39914 10370 39930
rect 10538 39802 10858 40041
rect 10993 40474 11089 40490
rect 10993 40410 11009 40474
rect 11073 40410 11089 40474
rect 10993 40394 11089 40410
rect 10993 40330 11009 40394
rect 11073 40330 11089 40394
rect 11258 40363 11578 40741
rect 11712 41030 11728 41094
rect 11792 41030 11808 41094
rect 12431 41174 12527 41190
rect 12431 41110 12447 41174
rect 12511 41110 12527 41174
rect 12431 41094 12527 41110
rect 11978 41063 12298 41082
rect 11712 41014 11808 41030
rect 11712 40950 11728 41014
rect 11792 40950 11808 41014
rect 11712 40934 11808 40950
rect 11712 40870 11728 40934
rect 11792 40870 11808 40934
rect 11712 40854 11808 40870
rect 11712 40790 11728 40854
rect 11792 40790 11808 40854
rect 11712 40774 11808 40790
rect 11712 40710 11728 40774
rect 11792 40710 11808 40774
rect 11971 41054 12298 41063
rect 11971 40750 11980 41054
rect 12284 40750 12298 41054
rect 11971 40741 12298 40750
rect 11712 40694 11808 40710
rect 11712 40630 11728 40694
rect 11792 40630 11808 40694
rect 11712 40614 11808 40630
rect 10993 40314 11089 40330
rect 10993 40250 11009 40314
rect 11073 40250 11089 40314
rect 10993 40234 11089 40250
rect 10993 40170 11009 40234
rect 11073 40170 11089 40234
rect 10993 40154 11089 40170
rect 10993 40090 11009 40154
rect 11073 40090 11089 40154
rect 10993 40074 11089 40090
rect 10993 40010 11009 40074
rect 11073 40010 11089 40074
rect 11252 40354 11578 40363
rect 11252 40050 11261 40354
rect 11565 40050 11578 40354
rect 11252 40041 11578 40050
rect 10993 39994 11089 40010
rect 10993 39930 11009 39994
rect 11073 39930 11089 39994
rect 10993 39914 11089 39930
rect 11258 39802 11578 40041
rect 11712 40474 11808 40490
rect 11712 40410 11728 40474
rect 11792 40410 11808 40474
rect 11712 40394 11808 40410
rect 11712 40330 11728 40394
rect 11792 40330 11808 40394
rect 11978 40363 12298 40741
rect 12431 41030 12447 41094
rect 12511 41030 12527 41094
rect 13150 41174 13246 41190
rect 13150 41110 13166 41174
rect 13230 41110 13246 41174
rect 13150 41094 13246 41110
rect 12698 41063 13018 41082
rect 12431 41014 12527 41030
rect 12431 40950 12447 41014
rect 12511 40950 12527 41014
rect 12431 40934 12527 40950
rect 12431 40870 12447 40934
rect 12511 40870 12527 40934
rect 12431 40854 12527 40870
rect 12431 40790 12447 40854
rect 12511 40790 12527 40854
rect 12431 40774 12527 40790
rect 12431 40710 12447 40774
rect 12511 40710 12527 40774
rect 12690 41054 13018 41063
rect 12690 40750 12699 41054
rect 13003 40750 13018 41054
rect 12690 40741 13018 40750
rect 12431 40694 12527 40710
rect 12431 40630 12447 40694
rect 12511 40630 12527 40694
rect 12431 40614 12527 40630
rect 11712 40314 11808 40330
rect 11712 40250 11728 40314
rect 11792 40250 11808 40314
rect 11712 40234 11808 40250
rect 11712 40170 11728 40234
rect 11792 40170 11808 40234
rect 11712 40154 11808 40170
rect 11712 40090 11728 40154
rect 11792 40090 11808 40154
rect 11712 40074 11808 40090
rect 11712 40010 11728 40074
rect 11792 40010 11808 40074
rect 11971 40354 12298 40363
rect 11971 40050 11980 40354
rect 12284 40050 12298 40354
rect 11971 40041 12298 40050
rect 11712 39994 11808 40010
rect 11712 39930 11728 39994
rect 11792 39930 11808 39994
rect 11712 39914 11808 39930
rect 11978 39802 12298 40041
rect 12431 40474 12527 40490
rect 12431 40410 12447 40474
rect 12511 40410 12527 40474
rect 12431 40394 12527 40410
rect 12431 40330 12447 40394
rect 12511 40330 12527 40394
rect 12698 40363 13018 40741
rect 13150 41030 13166 41094
rect 13230 41030 13246 41094
rect 13869 41174 13965 41190
rect 13869 41110 13885 41174
rect 13949 41110 13965 41174
rect 13869 41094 13965 41110
rect 13418 41063 13738 41082
rect 13150 41014 13246 41030
rect 13150 40950 13166 41014
rect 13230 40950 13246 41014
rect 13150 40934 13246 40950
rect 13150 40870 13166 40934
rect 13230 40870 13246 40934
rect 13150 40854 13246 40870
rect 13150 40790 13166 40854
rect 13230 40790 13246 40854
rect 13150 40774 13246 40790
rect 13150 40710 13166 40774
rect 13230 40710 13246 40774
rect 13409 41054 13738 41063
rect 13409 40750 13418 41054
rect 13722 40750 13738 41054
rect 13409 40741 13738 40750
rect 13150 40694 13246 40710
rect 13150 40630 13166 40694
rect 13230 40630 13246 40694
rect 13150 40614 13246 40630
rect 12431 40314 12527 40330
rect 12431 40250 12447 40314
rect 12511 40250 12527 40314
rect 12431 40234 12527 40250
rect 12431 40170 12447 40234
rect 12511 40170 12527 40234
rect 12431 40154 12527 40170
rect 12431 40090 12447 40154
rect 12511 40090 12527 40154
rect 12431 40074 12527 40090
rect 12431 40010 12447 40074
rect 12511 40010 12527 40074
rect 12690 40354 13018 40363
rect 12690 40050 12699 40354
rect 13003 40050 13018 40354
rect 12690 40041 13018 40050
rect 12431 39994 12527 40010
rect 12431 39930 12447 39994
rect 12511 39930 12527 39994
rect 12431 39914 12527 39930
rect 12698 39802 13018 40041
rect 13150 40474 13246 40490
rect 13150 40410 13166 40474
rect 13230 40410 13246 40474
rect 13150 40394 13246 40410
rect 13150 40330 13166 40394
rect 13230 40330 13246 40394
rect 13418 40363 13738 40741
rect 13869 41030 13885 41094
rect 13949 41030 13965 41094
rect 13869 41014 13965 41030
rect 13869 40950 13885 41014
rect 13949 40950 13965 41014
rect 13869 40934 13965 40950
rect 13869 40870 13885 40934
rect 13949 40870 13965 40934
rect 13869 40854 13965 40870
rect 13869 40790 13885 40854
rect 13949 40790 13965 40854
rect 13869 40774 13965 40790
rect 13869 40710 13885 40774
rect 13949 40710 13965 40774
rect 13869 40694 13965 40710
rect 13869 40630 13885 40694
rect 13949 40630 13965 40694
rect 13869 40614 13965 40630
rect 13150 40314 13246 40330
rect 13150 40250 13166 40314
rect 13230 40250 13246 40314
rect 13150 40234 13246 40250
rect 13150 40170 13166 40234
rect 13230 40170 13246 40234
rect 13150 40154 13246 40170
rect 13150 40090 13166 40154
rect 13230 40090 13246 40154
rect 13150 40074 13246 40090
rect 13150 40010 13166 40074
rect 13230 40010 13246 40074
rect 13409 40354 13738 40363
rect 13409 40050 13418 40354
rect 13722 40050 13738 40354
rect 13409 40041 13738 40050
rect 13150 39994 13246 40010
rect 13150 39930 13166 39994
rect 13230 39930 13246 39994
rect 13150 39914 13246 39930
rect 13418 39802 13738 40041
rect 13869 40474 13965 40490
rect 13869 40410 13885 40474
rect 13949 40410 13965 40474
rect 13869 40394 13965 40410
rect 13869 40330 13885 40394
rect 13949 40330 13965 40394
rect 13869 40314 13965 40330
rect 13869 40250 13885 40314
rect 13949 40250 13965 40314
rect 13869 40234 13965 40250
rect 13869 40170 13885 40234
rect 13949 40170 13965 40234
rect 13869 40154 13965 40170
rect 13869 40090 13885 40154
rect 13949 40090 13965 40154
rect 13869 40074 13965 40090
rect 13869 40010 13885 40074
rect 13949 40010 13965 40074
rect 13869 39994 13965 40010
rect 13869 39930 13885 39994
rect 13949 39930 13965 39994
rect 13869 39914 13965 39930
rect 6800 39774 13968 39802
rect 6800 39710 6828 39774
rect 6892 39710 6908 39774
rect 6972 39710 13968 39774
rect 6800 39694 13968 39710
rect 6800 39682 13676 39694
rect 13675 39630 13676 39682
rect 13740 39682 13968 39694
rect 27613 39694 27679 39695
rect 13740 39630 13741 39682
rect 13675 39629 13741 39630
rect 27613 39630 27614 39694
rect 27678 39630 27679 39694
rect 27613 39629 27679 39630
rect 3348 37640 3372 37704
rect 3436 37640 3452 37704
rect 3516 37640 3532 37704
rect 3596 37640 3612 37704
rect 3676 37640 3692 37704
rect 3756 37640 3772 37704
rect 3836 37640 3852 37704
rect 3916 37640 3932 37704
rect 3996 37640 4012 37704
rect 4076 37640 4092 37704
rect 4156 37640 4172 37704
rect 4236 37640 4252 37704
rect 4316 37640 4332 37704
rect 4396 37640 4412 37704
rect 4476 37640 4492 37704
rect 4556 37640 4572 37704
rect 4636 37640 4652 37704
rect 4716 37640 4732 37704
rect 4796 37640 4812 37704
rect 4876 37640 4892 37704
rect 4956 37640 4980 37704
rect 3348 33944 4980 37640
rect 12985 37620 13051 37621
rect 12985 37556 12986 37620
rect 13050 37556 13051 37620
rect 12985 37555 13051 37556
rect 12988 37430 13048 37555
rect 6516 37414 6612 37430
rect 6516 37350 6532 37414
rect 6596 37350 6612 37414
rect 6516 37334 6612 37350
rect 6056 37303 6376 37322
rect 6056 37294 6378 37303
rect 6056 36990 6065 37294
rect 6369 36990 6378 37294
rect 6056 36981 6378 36990
rect 6516 37270 6532 37334
rect 6596 37270 6612 37334
rect 7235 37414 7331 37430
rect 7235 37350 7251 37414
rect 7315 37350 7331 37414
rect 7235 37334 7331 37350
rect 6776 37303 7096 37322
rect 6516 37254 6612 37270
rect 6516 37190 6532 37254
rect 6596 37190 6612 37254
rect 6516 37174 6612 37190
rect 6516 37110 6532 37174
rect 6596 37110 6612 37174
rect 6516 37094 6612 37110
rect 6516 37030 6532 37094
rect 6596 37030 6612 37094
rect 6516 37014 6612 37030
rect 6056 36603 6376 36981
rect 6516 36950 6532 37014
rect 6596 36950 6612 37014
rect 6775 37294 7097 37303
rect 6775 36990 6784 37294
rect 7088 36990 7097 37294
rect 6775 36981 7097 36990
rect 7235 37270 7251 37334
rect 7315 37270 7331 37334
rect 7954 37414 8050 37430
rect 7954 37350 7970 37414
rect 8034 37350 8050 37414
rect 7954 37334 8050 37350
rect 7496 37303 7816 37322
rect 7235 37254 7331 37270
rect 7235 37190 7251 37254
rect 7315 37190 7331 37254
rect 7235 37174 7331 37190
rect 7235 37110 7251 37174
rect 7315 37110 7331 37174
rect 7235 37094 7331 37110
rect 7235 37030 7251 37094
rect 7315 37030 7331 37094
rect 7235 37014 7331 37030
rect 6516 36934 6612 36950
rect 6516 36870 6532 36934
rect 6596 36870 6612 36934
rect 6516 36854 6612 36870
rect 6516 36714 6612 36730
rect 6516 36650 6532 36714
rect 6596 36650 6612 36714
rect 6516 36634 6612 36650
rect 6056 36594 6378 36603
rect 6056 36290 6065 36594
rect 6369 36290 6378 36594
rect 6056 36281 6378 36290
rect 6516 36570 6532 36634
rect 6596 36570 6612 36634
rect 6776 36603 7096 36981
rect 7235 36950 7251 37014
rect 7315 36950 7331 37014
rect 7494 37294 7816 37303
rect 7494 36990 7503 37294
rect 7807 36990 7816 37294
rect 7494 36981 7816 36990
rect 7235 36934 7331 36950
rect 7235 36870 7251 36934
rect 7315 36870 7331 36934
rect 7235 36854 7331 36870
rect 7235 36714 7331 36730
rect 7235 36650 7251 36714
rect 7315 36650 7331 36714
rect 7235 36634 7331 36650
rect 6516 36554 6612 36570
rect 6516 36490 6532 36554
rect 6596 36490 6612 36554
rect 6516 36474 6612 36490
rect 6516 36410 6532 36474
rect 6596 36410 6612 36474
rect 6516 36394 6612 36410
rect 6516 36330 6532 36394
rect 6596 36330 6612 36394
rect 6516 36314 6612 36330
rect 6056 36042 6376 36281
rect 6516 36250 6532 36314
rect 6596 36250 6612 36314
rect 6775 36594 7097 36603
rect 6775 36290 6784 36594
rect 7088 36290 7097 36594
rect 6775 36281 7097 36290
rect 7235 36570 7251 36634
rect 7315 36570 7331 36634
rect 7496 36603 7816 36981
rect 7954 37270 7970 37334
rect 8034 37270 8050 37334
rect 8673 37414 8769 37430
rect 8673 37350 8689 37414
rect 8753 37350 8769 37414
rect 8673 37334 8769 37350
rect 8216 37303 8536 37322
rect 7954 37254 8050 37270
rect 7954 37190 7970 37254
rect 8034 37190 8050 37254
rect 7954 37174 8050 37190
rect 7954 37110 7970 37174
rect 8034 37110 8050 37174
rect 7954 37094 8050 37110
rect 7954 37030 7970 37094
rect 8034 37030 8050 37094
rect 7954 37014 8050 37030
rect 7954 36950 7970 37014
rect 8034 36950 8050 37014
rect 8213 37294 8536 37303
rect 8213 36990 8222 37294
rect 8526 36990 8536 37294
rect 8213 36981 8536 36990
rect 7954 36934 8050 36950
rect 7954 36870 7970 36934
rect 8034 36870 8050 36934
rect 7954 36854 8050 36870
rect 7235 36554 7331 36570
rect 7235 36490 7251 36554
rect 7315 36490 7331 36554
rect 7235 36474 7331 36490
rect 7235 36410 7251 36474
rect 7315 36410 7331 36474
rect 7235 36394 7331 36410
rect 7235 36330 7251 36394
rect 7315 36330 7331 36394
rect 7235 36314 7331 36330
rect 6516 36234 6612 36250
rect 6516 36170 6532 36234
rect 6596 36170 6612 36234
rect 6516 36154 6612 36170
rect 6776 36042 7096 36281
rect 7235 36250 7251 36314
rect 7315 36250 7331 36314
rect 7494 36594 7816 36603
rect 7494 36290 7503 36594
rect 7807 36290 7816 36594
rect 7494 36281 7816 36290
rect 7235 36234 7331 36250
rect 7235 36170 7251 36234
rect 7315 36170 7331 36234
rect 7235 36154 7331 36170
rect 7496 36042 7816 36281
rect 7954 36714 8050 36730
rect 7954 36650 7970 36714
rect 8034 36650 8050 36714
rect 7954 36634 8050 36650
rect 7954 36570 7970 36634
rect 8034 36570 8050 36634
rect 8216 36603 8536 36981
rect 8673 37270 8689 37334
rect 8753 37270 8769 37334
rect 9392 37414 9488 37430
rect 9392 37350 9408 37414
rect 9472 37350 9488 37414
rect 9392 37334 9488 37350
rect 8936 37303 9256 37322
rect 8673 37254 8769 37270
rect 8673 37190 8689 37254
rect 8753 37190 8769 37254
rect 8673 37174 8769 37190
rect 8673 37110 8689 37174
rect 8753 37110 8769 37174
rect 8673 37094 8769 37110
rect 8673 37030 8689 37094
rect 8753 37030 8769 37094
rect 8673 37014 8769 37030
rect 8673 36950 8689 37014
rect 8753 36950 8769 37014
rect 8932 37294 9256 37303
rect 8932 36990 8941 37294
rect 9245 36990 9256 37294
rect 8932 36981 9256 36990
rect 8673 36934 8769 36950
rect 8673 36870 8689 36934
rect 8753 36870 8769 36934
rect 8673 36854 8769 36870
rect 7954 36554 8050 36570
rect 7954 36490 7970 36554
rect 8034 36490 8050 36554
rect 7954 36474 8050 36490
rect 7954 36410 7970 36474
rect 8034 36410 8050 36474
rect 7954 36394 8050 36410
rect 7954 36330 7970 36394
rect 8034 36330 8050 36394
rect 7954 36314 8050 36330
rect 7954 36250 7970 36314
rect 8034 36250 8050 36314
rect 8213 36594 8536 36603
rect 8213 36290 8222 36594
rect 8526 36290 8536 36594
rect 8213 36281 8536 36290
rect 7954 36234 8050 36250
rect 7954 36170 7970 36234
rect 8034 36170 8050 36234
rect 7954 36154 8050 36170
rect 8216 36042 8536 36281
rect 8673 36714 8769 36730
rect 8673 36650 8689 36714
rect 8753 36650 8769 36714
rect 8673 36634 8769 36650
rect 8673 36570 8689 36634
rect 8753 36570 8769 36634
rect 8936 36603 9256 36981
rect 9392 37270 9408 37334
rect 9472 37270 9488 37334
rect 10111 37414 10207 37430
rect 10111 37350 10127 37414
rect 10191 37350 10207 37414
rect 10111 37334 10207 37350
rect 9656 37303 9976 37322
rect 9392 37254 9488 37270
rect 9392 37190 9408 37254
rect 9472 37190 9488 37254
rect 9392 37174 9488 37190
rect 9392 37110 9408 37174
rect 9472 37110 9488 37174
rect 9392 37094 9488 37110
rect 9392 37030 9408 37094
rect 9472 37030 9488 37094
rect 9392 37014 9488 37030
rect 9392 36950 9408 37014
rect 9472 36950 9488 37014
rect 9651 37294 9976 37303
rect 9651 36990 9660 37294
rect 9964 36990 9976 37294
rect 9651 36981 9976 36990
rect 9392 36934 9488 36950
rect 9392 36870 9408 36934
rect 9472 36870 9488 36934
rect 9392 36854 9488 36870
rect 8673 36554 8769 36570
rect 8673 36490 8689 36554
rect 8753 36490 8769 36554
rect 8673 36474 8769 36490
rect 8673 36410 8689 36474
rect 8753 36410 8769 36474
rect 8673 36394 8769 36410
rect 8673 36330 8689 36394
rect 8753 36330 8769 36394
rect 8673 36314 8769 36330
rect 8673 36250 8689 36314
rect 8753 36250 8769 36314
rect 8932 36594 9256 36603
rect 8932 36290 8941 36594
rect 9245 36290 9256 36594
rect 8932 36281 9256 36290
rect 8673 36234 8769 36250
rect 8673 36170 8689 36234
rect 8753 36170 8769 36234
rect 8673 36154 8769 36170
rect 8936 36042 9256 36281
rect 9392 36714 9488 36730
rect 9392 36650 9408 36714
rect 9472 36650 9488 36714
rect 9392 36634 9488 36650
rect 9392 36570 9408 36634
rect 9472 36570 9488 36634
rect 9656 36603 9976 36981
rect 10111 37270 10127 37334
rect 10191 37270 10207 37334
rect 10830 37414 10926 37430
rect 10830 37350 10846 37414
rect 10910 37350 10926 37414
rect 10830 37334 10926 37350
rect 10376 37303 10696 37322
rect 10111 37254 10207 37270
rect 10111 37190 10127 37254
rect 10191 37190 10207 37254
rect 10111 37174 10207 37190
rect 10111 37110 10127 37174
rect 10191 37110 10207 37174
rect 10111 37094 10207 37110
rect 10111 37030 10127 37094
rect 10191 37030 10207 37094
rect 10111 37014 10207 37030
rect 10111 36950 10127 37014
rect 10191 36950 10207 37014
rect 10370 37294 10696 37303
rect 10370 36990 10379 37294
rect 10683 36990 10696 37294
rect 10370 36981 10696 36990
rect 10111 36934 10207 36950
rect 10111 36870 10127 36934
rect 10191 36870 10207 36934
rect 10111 36854 10207 36870
rect 9392 36554 9488 36570
rect 9392 36490 9408 36554
rect 9472 36490 9488 36554
rect 9392 36474 9488 36490
rect 9392 36410 9408 36474
rect 9472 36410 9488 36474
rect 9392 36394 9488 36410
rect 9392 36330 9408 36394
rect 9472 36330 9488 36394
rect 9392 36314 9488 36330
rect 9392 36250 9408 36314
rect 9472 36250 9488 36314
rect 9651 36594 9976 36603
rect 9651 36290 9660 36594
rect 9964 36290 9976 36594
rect 9651 36281 9976 36290
rect 9392 36234 9488 36250
rect 9392 36170 9408 36234
rect 9472 36170 9488 36234
rect 9392 36154 9488 36170
rect 9656 36042 9976 36281
rect 10111 36714 10207 36730
rect 10111 36650 10127 36714
rect 10191 36650 10207 36714
rect 10111 36634 10207 36650
rect 10111 36570 10127 36634
rect 10191 36570 10207 36634
rect 10376 36603 10696 36981
rect 10830 37270 10846 37334
rect 10910 37270 10926 37334
rect 11549 37414 11645 37430
rect 11549 37350 11565 37414
rect 11629 37350 11645 37414
rect 11549 37334 11645 37350
rect 11096 37303 11416 37322
rect 10830 37254 10926 37270
rect 10830 37190 10846 37254
rect 10910 37190 10926 37254
rect 10830 37174 10926 37190
rect 10830 37110 10846 37174
rect 10910 37110 10926 37174
rect 10830 37094 10926 37110
rect 10830 37030 10846 37094
rect 10910 37030 10926 37094
rect 10830 37014 10926 37030
rect 10830 36950 10846 37014
rect 10910 36950 10926 37014
rect 11089 37294 11416 37303
rect 11089 36990 11098 37294
rect 11402 36990 11416 37294
rect 11089 36981 11416 36990
rect 10830 36934 10926 36950
rect 10830 36870 10846 36934
rect 10910 36870 10926 36934
rect 10830 36854 10926 36870
rect 10111 36554 10207 36570
rect 10111 36490 10127 36554
rect 10191 36490 10207 36554
rect 10111 36474 10207 36490
rect 10111 36410 10127 36474
rect 10191 36410 10207 36474
rect 10111 36394 10207 36410
rect 10111 36330 10127 36394
rect 10191 36330 10207 36394
rect 10111 36314 10207 36330
rect 10111 36250 10127 36314
rect 10191 36250 10207 36314
rect 10370 36594 10696 36603
rect 10370 36290 10379 36594
rect 10683 36290 10696 36594
rect 10370 36281 10696 36290
rect 10111 36234 10207 36250
rect 10111 36170 10127 36234
rect 10191 36170 10207 36234
rect 10111 36154 10207 36170
rect 10376 36042 10696 36281
rect 10830 36714 10926 36730
rect 10830 36650 10846 36714
rect 10910 36650 10926 36714
rect 10830 36634 10926 36650
rect 10830 36570 10846 36634
rect 10910 36570 10926 36634
rect 11096 36603 11416 36981
rect 11549 37270 11565 37334
rect 11629 37270 11645 37334
rect 12268 37414 12364 37430
rect 12268 37350 12284 37414
rect 12348 37350 12364 37414
rect 12268 37334 12364 37350
rect 11816 37303 12136 37322
rect 11549 37254 11645 37270
rect 11549 37190 11565 37254
rect 11629 37190 11645 37254
rect 11549 37174 11645 37190
rect 11549 37110 11565 37174
rect 11629 37110 11645 37174
rect 11549 37094 11645 37110
rect 11549 37030 11565 37094
rect 11629 37030 11645 37094
rect 11549 37014 11645 37030
rect 11549 36950 11565 37014
rect 11629 36950 11645 37014
rect 11808 37294 12136 37303
rect 11808 36990 11817 37294
rect 12121 36990 12136 37294
rect 11808 36981 12136 36990
rect 11549 36934 11645 36950
rect 11549 36870 11565 36934
rect 11629 36870 11645 36934
rect 11549 36854 11645 36870
rect 10830 36554 10926 36570
rect 10830 36490 10846 36554
rect 10910 36490 10926 36554
rect 10830 36474 10926 36490
rect 10830 36410 10846 36474
rect 10910 36410 10926 36474
rect 10830 36394 10926 36410
rect 10830 36330 10846 36394
rect 10910 36330 10926 36394
rect 10830 36314 10926 36330
rect 10830 36250 10846 36314
rect 10910 36250 10926 36314
rect 11089 36594 11416 36603
rect 11089 36290 11098 36594
rect 11402 36290 11416 36594
rect 11089 36281 11416 36290
rect 10830 36234 10926 36250
rect 10830 36170 10846 36234
rect 10910 36170 10926 36234
rect 10830 36154 10926 36170
rect 11096 36042 11416 36281
rect 11549 36714 11645 36730
rect 11549 36650 11565 36714
rect 11629 36650 11645 36714
rect 11549 36634 11645 36650
rect 11549 36570 11565 36634
rect 11629 36570 11645 36634
rect 11816 36603 12136 36981
rect 12268 37270 12284 37334
rect 12348 37270 12364 37334
rect 12987 37414 13083 37430
rect 12987 37350 13003 37414
rect 13067 37350 13083 37414
rect 12987 37334 13083 37350
rect 12536 37303 12856 37322
rect 12268 37254 12364 37270
rect 12268 37190 12284 37254
rect 12348 37190 12364 37254
rect 12268 37174 12364 37190
rect 12268 37110 12284 37174
rect 12348 37110 12364 37174
rect 12268 37094 12364 37110
rect 12268 37030 12284 37094
rect 12348 37030 12364 37094
rect 12268 37014 12364 37030
rect 12268 36950 12284 37014
rect 12348 36950 12364 37014
rect 12527 37294 12856 37303
rect 12527 36990 12536 37294
rect 12840 36990 12856 37294
rect 12527 36981 12856 36990
rect 12268 36934 12364 36950
rect 12268 36870 12284 36934
rect 12348 36870 12364 36934
rect 12268 36854 12364 36870
rect 11549 36554 11645 36570
rect 11549 36490 11565 36554
rect 11629 36490 11645 36554
rect 11549 36474 11645 36490
rect 11549 36410 11565 36474
rect 11629 36410 11645 36474
rect 11549 36394 11645 36410
rect 11549 36330 11565 36394
rect 11629 36330 11645 36394
rect 11549 36314 11645 36330
rect 11549 36250 11565 36314
rect 11629 36250 11645 36314
rect 11808 36594 12136 36603
rect 11808 36290 11817 36594
rect 12121 36290 12136 36594
rect 11808 36281 12136 36290
rect 11549 36234 11645 36250
rect 11549 36170 11565 36234
rect 11629 36170 11645 36234
rect 11549 36154 11645 36170
rect 11816 36042 12136 36281
rect 12268 36714 12364 36730
rect 12268 36650 12284 36714
rect 12348 36650 12364 36714
rect 12268 36634 12364 36650
rect 12268 36570 12284 36634
rect 12348 36570 12364 36634
rect 12536 36603 12856 36981
rect 12987 37270 13003 37334
rect 13067 37270 13083 37334
rect 13678 37322 13738 39629
rect 16849 37620 16915 37621
rect 16849 37556 16850 37620
rect 16914 37556 16915 37620
rect 16849 37555 16915 37556
rect 16852 37430 16912 37555
rect 13964 37414 14060 37430
rect 13964 37350 13980 37414
rect 14044 37350 14060 37414
rect 13964 37334 14060 37350
rect 12987 37254 13083 37270
rect 12987 37190 13003 37254
rect 13067 37190 13083 37254
rect 12987 37174 13083 37190
rect 12987 37110 13003 37174
rect 13067 37110 13083 37174
rect 12987 37094 13083 37110
rect 12987 37030 13003 37094
rect 13067 37030 13083 37094
rect 12987 37014 13083 37030
rect 12987 36950 13003 37014
rect 13067 36950 13083 37014
rect 12987 36934 13083 36950
rect 12987 36870 13003 36934
rect 13067 36870 13083 36934
rect 12987 36854 13083 36870
rect 13504 37303 13824 37322
rect 13504 37294 13826 37303
rect 13504 36990 13513 37294
rect 13817 36990 13826 37294
rect 13504 36981 13826 36990
rect 13964 37270 13980 37334
rect 14044 37270 14060 37334
rect 14683 37414 14779 37430
rect 14683 37350 14699 37414
rect 14763 37350 14779 37414
rect 14683 37334 14779 37350
rect 14224 37303 14544 37322
rect 13964 37254 14060 37270
rect 13964 37190 13980 37254
rect 14044 37190 14060 37254
rect 13964 37174 14060 37190
rect 13964 37110 13980 37174
rect 14044 37110 14060 37174
rect 13964 37094 14060 37110
rect 13964 37030 13980 37094
rect 14044 37030 14060 37094
rect 13964 37014 14060 37030
rect 12268 36554 12364 36570
rect 12268 36490 12284 36554
rect 12348 36490 12364 36554
rect 12268 36474 12364 36490
rect 12268 36410 12284 36474
rect 12348 36410 12364 36474
rect 12268 36394 12364 36410
rect 12268 36330 12284 36394
rect 12348 36330 12364 36394
rect 12268 36314 12364 36330
rect 12268 36250 12284 36314
rect 12348 36250 12364 36314
rect 12527 36594 12856 36603
rect 12527 36290 12536 36594
rect 12840 36290 12856 36594
rect 12527 36281 12856 36290
rect 12268 36234 12364 36250
rect 12268 36170 12284 36234
rect 12348 36170 12364 36234
rect 12268 36154 12364 36170
rect 12536 36042 12856 36281
rect 12987 36714 13083 36730
rect 12987 36650 13003 36714
rect 13067 36650 13083 36714
rect 12987 36634 13083 36650
rect 12987 36570 13003 36634
rect 13067 36570 13083 36634
rect 12987 36554 13083 36570
rect 12987 36490 13003 36554
rect 13067 36490 13083 36554
rect 12987 36474 13083 36490
rect 12987 36410 13003 36474
rect 13067 36410 13083 36474
rect 12987 36394 13083 36410
rect 12987 36330 13003 36394
rect 13067 36330 13083 36394
rect 12987 36314 13083 36330
rect 12987 36250 13003 36314
rect 13067 36250 13083 36314
rect 12987 36234 13083 36250
rect 12987 36170 13003 36234
rect 13067 36170 13083 36234
rect 12987 36154 13083 36170
rect 13504 36603 13824 36981
rect 13964 36950 13980 37014
rect 14044 36950 14060 37014
rect 14223 37294 14545 37303
rect 14223 36990 14232 37294
rect 14536 36990 14545 37294
rect 14223 36981 14545 36990
rect 14683 37270 14699 37334
rect 14763 37270 14779 37334
rect 15402 37414 15498 37430
rect 15402 37350 15418 37414
rect 15482 37350 15498 37414
rect 15402 37334 15498 37350
rect 14944 37303 15264 37322
rect 14683 37254 14779 37270
rect 14683 37190 14699 37254
rect 14763 37190 14779 37254
rect 14683 37174 14779 37190
rect 14683 37110 14699 37174
rect 14763 37110 14779 37174
rect 14683 37094 14779 37110
rect 14683 37030 14699 37094
rect 14763 37030 14779 37094
rect 14683 37014 14779 37030
rect 13964 36934 14060 36950
rect 13964 36870 13980 36934
rect 14044 36870 14060 36934
rect 13964 36854 14060 36870
rect 13964 36714 14060 36730
rect 13964 36650 13980 36714
rect 14044 36650 14060 36714
rect 13964 36634 14060 36650
rect 13504 36594 13826 36603
rect 13504 36290 13513 36594
rect 13817 36290 13826 36594
rect 13504 36281 13826 36290
rect 13964 36570 13980 36634
rect 14044 36570 14060 36634
rect 14224 36603 14544 36981
rect 14683 36950 14699 37014
rect 14763 36950 14779 37014
rect 14942 37294 15264 37303
rect 14942 36990 14951 37294
rect 15255 36990 15264 37294
rect 14942 36981 15264 36990
rect 14683 36934 14779 36950
rect 14683 36870 14699 36934
rect 14763 36870 14779 36934
rect 14683 36854 14779 36870
rect 14683 36714 14779 36730
rect 14683 36650 14699 36714
rect 14763 36650 14779 36714
rect 14683 36634 14779 36650
rect 13964 36554 14060 36570
rect 13964 36490 13980 36554
rect 14044 36490 14060 36554
rect 13964 36474 14060 36490
rect 13964 36410 13980 36474
rect 14044 36410 14060 36474
rect 13964 36394 14060 36410
rect 13964 36330 13980 36394
rect 14044 36330 14060 36394
rect 13964 36314 14060 36330
rect 13504 36042 13824 36281
rect 13964 36250 13980 36314
rect 14044 36250 14060 36314
rect 14223 36594 14545 36603
rect 14223 36290 14232 36594
rect 14536 36290 14545 36594
rect 14223 36281 14545 36290
rect 14683 36570 14699 36634
rect 14763 36570 14779 36634
rect 14944 36603 15264 36981
rect 15402 37270 15418 37334
rect 15482 37270 15498 37334
rect 16121 37414 16217 37430
rect 16121 37350 16137 37414
rect 16201 37350 16217 37414
rect 16121 37334 16217 37350
rect 15664 37303 15984 37322
rect 15402 37254 15498 37270
rect 15402 37190 15418 37254
rect 15482 37190 15498 37254
rect 15402 37174 15498 37190
rect 15402 37110 15418 37174
rect 15482 37110 15498 37174
rect 15402 37094 15498 37110
rect 15402 37030 15418 37094
rect 15482 37030 15498 37094
rect 15402 37014 15498 37030
rect 15402 36950 15418 37014
rect 15482 36950 15498 37014
rect 15661 37294 15984 37303
rect 15661 36990 15670 37294
rect 15974 36990 15984 37294
rect 15661 36981 15984 36990
rect 15402 36934 15498 36950
rect 15402 36870 15418 36934
rect 15482 36870 15498 36934
rect 15402 36854 15498 36870
rect 14683 36554 14779 36570
rect 14683 36490 14699 36554
rect 14763 36490 14779 36554
rect 14683 36474 14779 36490
rect 14683 36410 14699 36474
rect 14763 36410 14779 36474
rect 14683 36394 14779 36410
rect 14683 36330 14699 36394
rect 14763 36330 14779 36394
rect 14683 36314 14779 36330
rect 13964 36234 14060 36250
rect 13964 36170 13980 36234
rect 14044 36170 14060 36234
rect 13964 36154 14060 36170
rect 14224 36042 14544 36281
rect 14683 36250 14699 36314
rect 14763 36250 14779 36314
rect 14942 36594 15264 36603
rect 14942 36290 14951 36594
rect 15255 36290 15264 36594
rect 14942 36281 15264 36290
rect 14683 36234 14779 36250
rect 14683 36170 14699 36234
rect 14763 36170 14779 36234
rect 14683 36154 14779 36170
rect 14944 36042 15264 36281
rect 15402 36714 15498 36730
rect 15402 36650 15418 36714
rect 15482 36650 15498 36714
rect 15402 36634 15498 36650
rect 15402 36570 15418 36634
rect 15482 36570 15498 36634
rect 15664 36603 15984 36981
rect 16121 37270 16137 37334
rect 16201 37270 16217 37334
rect 16840 37414 16936 37430
rect 16840 37350 16856 37414
rect 16920 37350 16936 37414
rect 16840 37334 16936 37350
rect 16384 37303 16704 37322
rect 16121 37254 16217 37270
rect 16121 37190 16137 37254
rect 16201 37190 16217 37254
rect 16121 37174 16217 37190
rect 16121 37110 16137 37174
rect 16201 37110 16217 37174
rect 16121 37094 16217 37110
rect 16121 37030 16137 37094
rect 16201 37030 16217 37094
rect 16121 37014 16217 37030
rect 16121 36950 16137 37014
rect 16201 36950 16217 37014
rect 16380 37294 16704 37303
rect 16380 36990 16389 37294
rect 16693 36990 16704 37294
rect 16380 36981 16704 36990
rect 16121 36934 16217 36950
rect 16121 36870 16137 36934
rect 16201 36870 16217 36934
rect 16121 36854 16217 36870
rect 15402 36554 15498 36570
rect 15402 36490 15418 36554
rect 15482 36490 15498 36554
rect 15402 36474 15498 36490
rect 15402 36410 15418 36474
rect 15482 36410 15498 36474
rect 15402 36394 15498 36410
rect 15402 36330 15418 36394
rect 15482 36330 15498 36394
rect 15402 36314 15498 36330
rect 15402 36250 15418 36314
rect 15482 36250 15498 36314
rect 15661 36594 15984 36603
rect 15661 36290 15670 36594
rect 15974 36290 15984 36594
rect 15661 36281 15984 36290
rect 15402 36234 15498 36250
rect 15402 36170 15418 36234
rect 15482 36170 15498 36234
rect 15402 36154 15498 36170
rect 15664 36042 15984 36281
rect 16121 36714 16217 36730
rect 16121 36650 16137 36714
rect 16201 36650 16217 36714
rect 16121 36634 16217 36650
rect 16121 36570 16137 36634
rect 16201 36570 16217 36634
rect 16384 36603 16704 36981
rect 16840 37270 16856 37334
rect 16920 37270 16936 37334
rect 17559 37414 17655 37430
rect 17559 37350 17575 37414
rect 17639 37350 17655 37414
rect 17559 37334 17655 37350
rect 17104 37303 17424 37322
rect 16840 37254 16936 37270
rect 16840 37190 16856 37254
rect 16920 37190 16936 37254
rect 16840 37174 16936 37190
rect 16840 37110 16856 37174
rect 16920 37110 16936 37174
rect 16840 37094 16936 37110
rect 16840 37030 16856 37094
rect 16920 37030 16936 37094
rect 16840 37014 16936 37030
rect 16840 36950 16856 37014
rect 16920 36950 16936 37014
rect 17099 37294 17424 37303
rect 17099 36990 17108 37294
rect 17412 36990 17424 37294
rect 17099 36981 17424 36990
rect 16840 36934 16936 36950
rect 16840 36870 16856 36934
rect 16920 36870 16936 36934
rect 16840 36854 16936 36870
rect 16121 36554 16217 36570
rect 16121 36490 16137 36554
rect 16201 36490 16217 36554
rect 16121 36474 16217 36490
rect 16121 36410 16137 36474
rect 16201 36410 16217 36474
rect 16121 36394 16217 36410
rect 16121 36330 16137 36394
rect 16201 36330 16217 36394
rect 16121 36314 16217 36330
rect 16121 36250 16137 36314
rect 16201 36250 16217 36314
rect 16380 36594 16704 36603
rect 16380 36290 16389 36594
rect 16693 36290 16704 36594
rect 16380 36281 16704 36290
rect 16121 36234 16217 36250
rect 16121 36170 16137 36234
rect 16201 36170 16217 36234
rect 16121 36154 16217 36170
rect 16384 36042 16704 36281
rect 16840 36714 16936 36730
rect 16840 36650 16856 36714
rect 16920 36650 16936 36714
rect 16840 36634 16936 36650
rect 16840 36570 16856 36634
rect 16920 36570 16936 36634
rect 17104 36603 17424 36981
rect 17559 37270 17575 37334
rect 17639 37270 17655 37334
rect 18278 37414 18374 37430
rect 18278 37350 18294 37414
rect 18358 37350 18374 37414
rect 18278 37334 18374 37350
rect 17824 37303 18144 37322
rect 17559 37254 17655 37270
rect 17559 37190 17575 37254
rect 17639 37190 17655 37254
rect 17559 37174 17655 37190
rect 17559 37110 17575 37174
rect 17639 37110 17655 37174
rect 17559 37094 17655 37110
rect 17559 37030 17575 37094
rect 17639 37030 17655 37094
rect 17559 37014 17655 37030
rect 17559 36950 17575 37014
rect 17639 36950 17655 37014
rect 17818 37294 18144 37303
rect 17818 36990 17827 37294
rect 18131 36990 18144 37294
rect 17818 36981 18144 36990
rect 17559 36934 17655 36950
rect 17559 36870 17575 36934
rect 17639 36870 17655 36934
rect 17559 36854 17655 36870
rect 16840 36554 16936 36570
rect 16840 36490 16856 36554
rect 16920 36490 16936 36554
rect 16840 36474 16936 36490
rect 16840 36410 16856 36474
rect 16920 36410 16936 36474
rect 16840 36394 16936 36410
rect 16840 36330 16856 36394
rect 16920 36330 16936 36394
rect 16840 36314 16936 36330
rect 16840 36250 16856 36314
rect 16920 36250 16936 36314
rect 17099 36594 17424 36603
rect 17099 36290 17108 36594
rect 17412 36290 17424 36594
rect 17099 36281 17424 36290
rect 16840 36234 16936 36250
rect 16840 36170 16856 36234
rect 16920 36170 16936 36234
rect 16840 36154 16936 36170
rect 17104 36042 17424 36281
rect 17559 36714 17655 36730
rect 17559 36650 17575 36714
rect 17639 36650 17655 36714
rect 17559 36634 17655 36650
rect 17559 36570 17575 36634
rect 17639 36570 17655 36634
rect 17824 36603 18144 36981
rect 18278 37270 18294 37334
rect 18358 37270 18374 37334
rect 18997 37414 19093 37430
rect 18997 37350 19013 37414
rect 19077 37350 19093 37414
rect 18997 37334 19093 37350
rect 18544 37303 18864 37322
rect 18278 37254 18374 37270
rect 18278 37190 18294 37254
rect 18358 37190 18374 37254
rect 18278 37174 18374 37190
rect 18278 37110 18294 37174
rect 18358 37110 18374 37174
rect 18278 37094 18374 37110
rect 18278 37030 18294 37094
rect 18358 37030 18374 37094
rect 18278 37014 18374 37030
rect 18278 36950 18294 37014
rect 18358 36950 18374 37014
rect 18537 37294 18864 37303
rect 18537 36990 18546 37294
rect 18850 36990 18864 37294
rect 18537 36981 18864 36990
rect 18278 36934 18374 36950
rect 18278 36870 18294 36934
rect 18358 36870 18374 36934
rect 18278 36854 18374 36870
rect 17559 36554 17655 36570
rect 17559 36490 17575 36554
rect 17639 36490 17655 36554
rect 17559 36474 17655 36490
rect 17559 36410 17575 36474
rect 17639 36410 17655 36474
rect 17559 36394 17655 36410
rect 17559 36330 17575 36394
rect 17639 36330 17655 36394
rect 17559 36314 17655 36330
rect 17559 36250 17575 36314
rect 17639 36250 17655 36314
rect 17818 36594 18144 36603
rect 17818 36290 17827 36594
rect 18131 36290 18144 36594
rect 17818 36281 18144 36290
rect 17559 36234 17655 36250
rect 17559 36170 17575 36234
rect 17639 36170 17655 36234
rect 17559 36154 17655 36170
rect 17824 36042 18144 36281
rect 18278 36714 18374 36730
rect 18278 36650 18294 36714
rect 18358 36650 18374 36714
rect 18278 36634 18374 36650
rect 18278 36570 18294 36634
rect 18358 36570 18374 36634
rect 18544 36603 18864 36981
rect 18997 37270 19013 37334
rect 19077 37270 19093 37334
rect 19716 37414 19812 37430
rect 19716 37350 19732 37414
rect 19796 37350 19812 37414
rect 19716 37334 19812 37350
rect 19264 37303 19584 37322
rect 18997 37254 19093 37270
rect 18997 37190 19013 37254
rect 19077 37190 19093 37254
rect 18997 37174 19093 37190
rect 18997 37110 19013 37174
rect 19077 37110 19093 37174
rect 18997 37094 19093 37110
rect 18997 37030 19013 37094
rect 19077 37030 19093 37094
rect 18997 37014 19093 37030
rect 18997 36950 19013 37014
rect 19077 36950 19093 37014
rect 19256 37294 19584 37303
rect 19256 36990 19265 37294
rect 19569 36990 19584 37294
rect 19256 36981 19584 36990
rect 18997 36934 19093 36950
rect 18997 36870 19013 36934
rect 19077 36870 19093 36934
rect 18997 36854 19093 36870
rect 18278 36554 18374 36570
rect 18278 36490 18294 36554
rect 18358 36490 18374 36554
rect 18278 36474 18374 36490
rect 18278 36410 18294 36474
rect 18358 36410 18374 36474
rect 18278 36394 18374 36410
rect 18278 36330 18294 36394
rect 18358 36330 18374 36394
rect 18278 36314 18374 36330
rect 18278 36250 18294 36314
rect 18358 36250 18374 36314
rect 18537 36594 18864 36603
rect 18537 36290 18546 36594
rect 18850 36290 18864 36594
rect 18537 36281 18864 36290
rect 18278 36234 18374 36250
rect 18278 36170 18294 36234
rect 18358 36170 18374 36234
rect 18278 36154 18374 36170
rect 18544 36042 18864 36281
rect 18997 36714 19093 36730
rect 18997 36650 19013 36714
rect 19077 36650 19093 36714
rect 18997 36634 19093 36650
rect 18997 36570 19013 36634
rect 19077 36570 19093 36634
rect 19264 36603 19584 36981
rect 19716 37270 19732 37334
rect 19796 37270 19812 37334
rect 20435 37414 20531 37430
rect 20435 37350 20451 37414
rect 20515 37350 20531 37414
rect 20435 37334 20531 37350
rect 19984 37303 20304 37322
rect 19716 37254 19812 37270
rect 19716 37190 19732 37254
rect 19796 37190 19812 37254
rect 19716 37174 19812 37190
rect 19716 37110 19732 37174
rect 19796 37110 19812 37174
rect 19716 37094 19812 37110
rect 19716 37030 19732 37094
rect 19796 37030 19812 37094
rect 19716 37014 19812 37030
rect 19716 36950 19732 37014
rect 19796 36950 19812 37014
rect 19975 37294 20304 37303
rect 19975 36990 19984 37294
rect 20288 36990 20304 37294
rect 19975 36981 20304 36990
rect 19716 36934 19812 36950
rect 19716 36870 19732 36934
rect 19796 36870 19812 36934
rect 19716 36854 19812 36870
rect 18997 36554 19093 36570
rect 18997 36490 19013 36554
rect 19077 36490 19093 36554
rect 18997 36474 19093 36490
rect 18997 36410 19013 36474
rect 19077 36410 19093 36474
rect 18997 36394 19093 36410
rect 18997 36330 19013 36394
rect 19077 36330 19093 36394
rect 18997 36314 19093 36330
rect 18997 36250 19013 36314
rect 19077 36250 19093 36314
rect 19256 36594 19584 36603
rect 19256 36290 19265 36594
rect 19569 36290 19584 36594
rect 19256 36281 19584 36290
rect 18997 36234 19093 36250
rect 18997 36170 19013 36234
rect 19077 36170 19093 36234
rect 18997 36154 19093 36170
rect 19264 36042 19584 36281
rect 19716 36714 19812 36730
rect 19716 36650 19732 36714
rect 19796 36650 19812 36714
rect 19716 36634 19812 36650
rect 19716 36570 19732 36634
rect 19796 36570 19812 36634
rect 19984 36603 20304 36981
rect 20435 37270 20451 37334
rect 20515 37270 20531 37334
rect 21412 37414 21508 37430
rect 21412 37350 21428 37414
rect 21492 37350 21508 37414
rect 21412 37334 21508 37350
rect 20435 37254 20531 37270
rect 20435 37190 20451 37254
rect 20515 37190 20531 37254
rect 20435 37174 20531 37190
rect 20435 37110 20451 37174
rect 20515 37110 20531 37174
rect 20435 37094 20531 37110
rect 20435 37030 20451 37094
rect 20515 37030 20531 37094
rect 20435 37014 20531 37030
rect 20435 36950 20451 37014
rect 20515 36950 20531 37014
rect 20435 36934 20531 36950
rect 20435 36870 20451 36934
rect 20515 36870 20531 36934
rect 20435 36854 20531 36870
rect 20952 37303 21272 37322
rect 20952 37294 21274 37303
rect 20952 36990 20961 37294
rect 21265 36990 21274 37294
rect 20952 36981 21274 36990
rect 21412 37270 21428 37334
rect 21492 37270 21508 37334
rect 22131 37414 22227 37430
rect 22131 37350 22147 37414
rect 22211 37350 22227 37414
rect 22131 37334 22227 37350
rect 21672 37303 21992 37322
rect 21412 37254 21508 37270
rect 21412 37190 21428 37254
rect 21492 37190 21508 37254
rect 21412 37174 21508 37190
rect 21412 37110 21428 37174
rect 21492 37110 21508 37174
rect 21412 37094 21508 37110
rect 21412 37030 21428 37094
rect 21492 37030 21508 37094
rect 21412 37014 21508 37030
rect 19716 36554 19812 36570
rect 19716 36490 19732 36554
rect 19796 36490 19812 36554
rect 19716 36474 19812 36490
rect 19716 36410 19732 36474
rect 19796 36410 19812 36474
rect 19716 36394 19812 36410
rect 19716 36330 19732 36394
rect 19796 36330 19812 36394
rect 19716 36314 19812 36330
rect 19716 36250 19732 36314
rect 19796 36250 19812 36314
rect 19975 36594 20304 36603
rect 19975 36290 19984 36594
rect 20288 36290 20304 36594
rect 19975 36281 20304 36290
rect 19716 36234 19812 36250
rect 19716 36170 19732 36234
rect 19796 36170 19812 36234
rect 19716 36154 19812 36170
rect 19984 36042 20304 36281
rect 20435 36714 20531 36730
rect 20435 36650 20451 36714
rect 20515 36650 20531 36714
rect 20435 36634 20531 36650
rect 20435 36570 20451 36634
rect 20515 36570 20531 36634
rect 20435 36554 20531 36570
rect 20435 36490 20451 36554
rect 20515 36490 20531 36554
rect 20435 36474 20531 36490
rect 20435 36410 20451 36474
rect 20515 36410 20531 36474
rect 20435 36394 20531 36410
rect 20435 36330 20451 36394
rect 20515 36330 20531 36394
rect 20435 36314 20531 36330
rect 20435 36250 20451 36314
rect 20515 36250 20531 36314
rect 20435 36234 20531 36250
rect 20435 36170 20451 36234
rect 20515 36170 20531 36234
rect 20435 36154 20531 36170
rect 20952 36603 21272 36981
rect 21412 36950 21428 37014
rect 21492 36950 21508 37014
rect 21671 37294 21993 37303
rect 21671 36990 21680 37294
rect 21984 36990 21993 37294
rect 21671 36981 21993 36990
rect 22131 37270 22147 37334
rect 22211 37270 22227 37334
rect 22850 37414 22946 37430
rect 22850 37350 22866 37414
rect 22930 37350 22946 37414
rect 22850 37334 22946 37350
rect 22392 37303 22712 37322
rect 22131 37254 22227 37270
rect 22131 37190 22147 37254
rect 22211 37190 22227 37254
rect 22131 37174 22227 37190
rect 22131 37110 22147 37174
rect 22211 37110 22227 37174
rect 22131 37094 22227 37110
rect 22131 37030 22147 37094
rect 22211 37030 22227 37094
rect 22131 37014 22227 37030
rect 21412 36934 21508 36950
rect 21412 36870 21428 36934
rect 21492 36870 21508 36934
rect 21412 36854 21508 36870
rect 21412 36714 21508 36730
rect 21412 36650 21428 36714
rect 21492 36650 21508 36714
rect 21412 36634 21508 36650
rect 20952 36594 21274 36603
rect 20952 36290 20961 36594
rect 21265 36290 21274 36594
rect 20952 36281 21274 36290
rect 21412 36570 21428 36634
rect 21492 36570 21508 36634
rect 21672 36603 21992 36981
rect 22131 36950 22147 37014
rect 22211 36950 22227 37014
rect 22390 37294 22712 37303
rect 22390 36990 22399 37294
rect 22703 36990 22712 37294
rect 22390 36981 22712 36990
rect 22131 36934 22227 36950
rect 22131 36870 22147 36934
rect 22211 36870 22227 36934
rect 22131 36854 22227 36870
rect 22131 36714 22227 36730
rect 22131 36650 22147 36714
rect 22211 36650 22227 36714
rect 22131 36634 22227 36650
rect 21412 36554 21508 36570
rect 21412 36490 21428 36554
rect 21492 36490 21508 36554
rect 21412 36474 21508 36490
rect 21412 36410 21428 36474
rect 21492 36410 21508 36474
rect 21412 36394 21508 36410
rect 21412 36330 21428 36394
rect 21492 36330 21508 36394
rect 21412 36314 21508 36330
rect 20952 36042 21272 36281
rect 21412 36250 21428 36314
rect 21492 36250 21508 36314
rect 21671 36594 21993 36603
rect 21671 36290 21680 36594
rect 21984 36290 21993 36594
rect 21671 36281 21993 36290
rect 22131 36570 22147 36634
rect 22211 36570 22227 36634
rect 22392 36603 22712 36981
rect 22850 37270 22866 37334
rect 22930 37270 22946 37334
rect 23569 37414 23665 37430
rect 23569 37350 23585 37414
rect 23649 37350 23665 37414
rect 23569 37334 23665 37350
rect 23112 37303 23432 37322
rect 22850 37254 22946 37270
rect 22850 37190 22866 37254
rect 22930 37190 22946 37254
rect 22850 37174 22946 37190
rect 22850 37110 22866 37174
rect 22930 37110 22946 37174
rect 22850 37094 22946 37110
rect 22850 37030 22866 37094
rect 22930 37030 22946 37094
rect 22850 37014 22946 37030
rect 22850 36950 22866 37014
rect 22930 36950 22946 37014
rect 23109 37294 23432 37303
rect 23109 36990 23118 37294
rect 23422 36990 23432 37294
rect 23109 36981 23432 36990
rect 22850 36934 22946 36950
rect 22850 36870 22866 36934
rect 22930 36870 22946 36934
rect 22850 36854 22946 36870
rect 22131 36554 22227 36570
rect 22131 36490 22147 36554
rect 22211 36490 22227 36554
rect 22131 36474 22227 36490
rect 22131 36410 22147 36474
rect 22211 36410 22227 36474
rect 22131 36394 22227 36410
rect 22131 36330 22147 36394
rect 22211 36330 22227 36394
rect 22131 36314 22227 36330
rect 21412 36234 21508 36250
rect 21412 36170 21428 36234
rect 21492 36170 21508 36234
rect 21412 36154 21508 36170
rect 21672 36042 21992 36281
rect 22131 36250 22147 36314
rect 22211 36250 22227 36314
rect 22390 36594 22712 36603
rect 22390 36290 22399 36594
rect 22703 36290 22712 36594
rect 22390 36281 22712 36290
rect 22131 36234 22227 36250
rect 22131 36170 22147 36234
rect 22211 36170 22227 36234
rect 22131 36154 22227 36170
rect 22392 36042 22712 36281
rect 22850 36714 22946 36730
rect 22850 36650 22866 36714
rect 22930 36650 22946 36714
rect 22850 36634 22946 36650
rect 22850 36570 22866 36634
rect 22930 36570 22946 36634
rect 23112 36603 23432 36981
rect 23569 37270 23585 37334
rect 23649 37270 23665 37334
rect 24288 37414 24384 37430
rect 24288 37350 24304 37414
rect 24368 37350 24384 37414
rect 24288 37334 24384 37350
rect 23832 37303 24152 37322
rect 23569 37254 23665 37270
rect 23569 37190 23585 37254
rect 23649 37190 23665 37254
rect 23569 37174 23665 37190
rect 23569 37110 23585 37174
rect 23649 37110 23665 37174
rect 23569 37094 23665 37110
rect 23569 37030 23585 37094
rect 23649 37030 23665 37094
rect 23569 37014 23665 37030
rect 23569 36950 23585 37014
rect 23649 36950 23665 37014
rect 23828 37294 24152 37303
rect 23828 36990 23837 37294
rect 24141 36990 24152 37294
rect 23828 36981 24152 36990
rect 23569 36934 23665 36950
rect 23569 36870 23585 36934
rect 23649 36870 23665 36934
rect 23569 36854 23665 36870
rect 22850 36554 22946 36570
rect 22850 36490 22866 36554
rect 22930 36490 22946 36554
rect 22850 36474 22946 36490
rect 22850 36410 22866 36474
rect 22930 36410 22946 36474
rect 22850 36394 22946 36410
rect 22850 36330 22866 36394
rect 22930 36330 22946 36394
rect 22850 36314 22946 36330
rect 22850 36250 22866 36314
rect 22930 36250 22946 36314
rect 23109 36594 23432 36603
rect 23109 36290 23118 36594
rect 23422 36290 23432 36594
rect 23109 36281 23432 36290
rect 22850 36234 22946 36250
rect 22850 36170 22866 36234
rect 22930 36170 22946 36234
rect 22850 36154 22946 36170
rect 23112 36042 23432 36281
rect 23569 36714 23665 36730
rect 23569 36650 23585 36714
rect 23649 36650 23665 36714
rect 23569 36634 23665 36650
rect 23569 36570 23585 36634
rect 23649 36570 23665 36634
rect 23832 36603 24152 36981
rect 24288 37270 24304 37334
rect 24368 37270 24384 37334
rect 25007 37414 25103 37430
rect 25007 37350 25023 37414
rect 25087 37350 25103 37414
rect 25007 37334 25103 37350
rect 24552 37303 24872 37322
rect 24288 37254 24384 37270
rect 24288 37190 24304 37254
rect 24368 37190 24384 37254
rect 24288 37174 24384 37190
rect 24288 37110 24304 37174
rect 24368 37110 24384 37174
rect 24288 37094 24384 37110
rect 24288 37030 24304 37094
rect 24368 37030 24384 37094
rect 24288 37014 24384 37030
rect 24288 36950 24304 37014
rect 24368 36950 24384 37014
rect 24547 37294 24872 37303
rect 24547 36990 24556 37294
rect 24860 36990 24872 37294
rect 24547 36981 24872 36990
rect 24288 36934 24384 36950
rect 24288 36870 24304 36934
rect 24368 36870 24384 36934
rect 24288 36854 24384 36870
rect 23569 36554 23665 36570
rect 23569 36490 23585 36554
rect 23649 36490 23665 36554
rect 23569 36474 23665 36490
rect 23569 36410 23585 36474
rect 23649 36410 23665 36474
rect 23569 36394 23665 36410
rect 23569 36330 23585 36394
rect 23649 36330 23665 36394
rect 23569 36314 23665 36330
rect 23569 36250 23585 36314
rect 23649 36250 23665 36314
rect 23828 36594 24152 36603
rect 23828 36290 23837 36594
rect 24141 36290 24152 36594
rect 23828 36281 24152 36290
rect 23569 36234 23665 36250
rect 23569 36170 23585 36234
rect 23649 36170 23665 36234
rect 23569 36154 23665 36170
rect 23832 36042 24152 36281
rect 24288 36714 24384 36730
rect 24288 36650 24304 36714
rect 24368 36650 24384 36714
rect 24288 36634 24384 36650
rect 24288 36570 24304 36634
rect 24368 36570 24384 36634
rect 24552 36603 24872 36981
rect 25007 37270 25023 37334
rect 25087 37270 25103 37334
rect 25726 37414 25822 37430
rect 25726 37350 25742 37414
rect 25806 37350 25822 37414
rect 25726 37334 25822 37350
rect 25272 37303 25592 37322
rect 25007 37254 25103 37270
rect 25007 37190 25023 37254
rect 25087 37190 25103 37254
rect 25007 37174 25103 37190
rect 25007 37110 25023 37174
rect 25087 37110 25103 37174
rect 25007 37094 25103 37110
rect 25007 37030 25023 37094
rect 25087 37030 25103 37094
rect 25007 37014 25103 37030
rect 25007 36950 25023 37014
rect 25087 36950 25103 37014
rect 25266 37294 25592 37303
rect 25266 36990 25275 37294
rect 25579 36990 25592 37294
rect 25266 36981 25592 36990
rect 25007 36934 25103 36950
rect 25007 36870 25023 36934
rect 25087 36870 25103 36934
rect 25007 36854 25103 36870
rect 24288 36554 24384 36570
rect 24288 36490 24304 36554
rect 24368 36490 24384 36554
rect 24288 36474 24384 36490
rect 24288 36410 24304 36474
rect 24368 36410 24384 36474
rect 24288 36394 24384 36410
rect 24288 36330 24304 36394
rect 24368 36330 24384 36394
rect 24288 36314 24384 36330
rect 24288 36250 24304 36314
rect 24368 36250 24384 36314
rect 24547 36594 24872 36603
rect 24547 36290 24556 36594
rect 24860 36290 24872 36594
rect 24547 36281 24872 36290
rect 24288 36234 24384 36250
rect 24288 36170 24304 36234
rect 24368 36170 24384 36234
rect 24288 36154 24384 36170
rect 24552 36042 24872 36281
rect 25007 36714 25103 36730
rect 25007 36650 25023 36714
rect 25087 36650 25103 36714
rect 25007 36634 25103 36650
rect 25007 36570 25023 36634
rect 25087 36570 25103 36634
rect 25272 36603 25592 36981
rect 25726 37270 25742 37334
rect 25806 37270 25822 37334
rect 26445 37414 26541 37430
rect 26445 37350 26461 37414
rect 26525 37350 26541 37414
rect 26445 37334 26541 37350
rect 25992 37303 26312 37322
rect 25726 37254 25822 37270
rect 25726 37190 25742 37254
rect 25806 37190 25822 37254
rect 25726 37174 25822 37190
rect 25726 37110 25742 37174
rect 25806 37110 25822 37174
rect 25726 37094 25822 37110
rect 25726 37030 25742 37094
rect 25806 37030 25822 37094
rect 25726 37014 25822 37030
rect 25726 36950 25742 37014
rect 25806 36950 25822 37014
rect 25985 37294 26312 37303
rect 25985 36990 25994 37294
rect 26298 36990 26312 37294
rect 25985 36981 26312 36990
rect 25726 36934 25822 36950
rect 25726 36870 25742 36934
rect 25806 36870 25822 36934
rect 25726 36854 25822 36870
rect 25007 36554 25103 36570
rect 25007 36490 25023 36554
rect 25087 36490 25103 36554
rect 25007 36474 25103 36490
rect 25007 36410 25023 36474
rect 25087 36410 25103 36474
rect 25007 36394 25103 36410
rect 25007 36330 25023 36394
rect 25087 36330 25103 36394
rect 25007 36314 25103 36330
rect 25007 36250 25023 36314
rect 25087 36250 25103 36314
rect 25266 36594 25592 36603
rect 25266 36290 25275 36594
rect 25579 36290 25592 36594
rect 25266 36281 25592 36290
rect 25007 36234 25103 36250
rect 25007 36170 25023 36234
rect 25087 36170 25103 36234
rect 25007 36154 25103 36170
rect 25272 36042 25592 36281
rect 25726 36714 25822 36730
rect 25726 36650 25742 36714
rect 25806 36650 25822 36714
rect 25726 36634 25822 36650
rect 25726 36570 25742 36634
rect 25806 36570 25822 36634
rect 25992 36603 26312 36981
rect 26445 37270 26461 37334
rect 26525 37270 26541 37334
rect 27164 37414 27260 37430
rect 27164 37350 27180 37414
rect 27244 37350 27260 37414
rect 27164 37334 27260 37350
rect 26712 37303 27032 37322
rect 26445 37254 26541 37270
rect 26445 37190 26461 37254
rect 26525 37190 26541 37254
rect 26445 37174 26541 37190
rect 26445 37110 26461 37174
rect 26525 37110 26541 37174
rect 26445 37094 26541 37110
rect 26445 37030 26461 37094
rect 26525 37030 26541 37094
rect 26445 37014 26541 37030
rect 26445 36950 26461 37014
rect 26525 36950 26541 37014
rect 26704 37294 27032 37303
rect 26704 36990 26713 37294
rect 27017 36990 27032 37294
rect 26704 36981 27032 36990
rect 26445 36934 26541 36950
rect 26445 36870 26461 36934
rect 26525 36870 26541 36934
rect 26445 36854 26541 36870
rect 25726 36554 25822 36570
rect 25726 36490 25742 36554
rect 25806 36490 25822 36554
rect 25726 36474 25822 36490
rect 25726 36410 25742 36474
rect 25806 36410 25822 36474
rect 25726 36394 25822 36410
rect 25726 36330 25742 36394
rect 25806 36330 25822 36394
rect 25726 36314 25822 36330
rect 25726 36250 25742 36314
rect 25806 36250 25822 36314
rect 25985 36594 26312 36603
rect 25985 36290 25994 36594
rect 26298 36290 26312 36594
rect 25985 36281 26312 36290
rect 25726 36234 25822 36250
rect 25726 36170 25742 36234
rect 25806 36170 25822 36234
rect 25726 36154 25822 36170
rect 25992 36042 26312 36281
rect 26445 36714 26541 36730
rect 26445 36650 26461 36714
rect 26525 36650 26541 36714
rect 26445 36634 26541 36650
rect 26445 36570 26461 36634
rect 26525 36570 26541 36634
rect 26712 36603 27032 36981
rect 27164 37270 27180 37334
rect 27244 37270 27260 37334
rect 27616 37322 27676 39629
rect 43656 37704 45288 41400
rect 43656 37640 43680 37704
rect 43744 37640 43760 37704
rect 43824 37640 43840 37704
rect 43904 37640 43920 37704
rect 43984 37640 44000 37704
rect 44064 37640 44080 37704
rect 44144 37640 44160 37704
rect 44224 37640 44240 37704
rect 44304 37640 44320 37704
rect 44384 37640 44400 37704
rect 44464 37640 44480 37704
rect 44544 37640 44560 37704
rect 44624 37640 44640 37704
rect 44704 37640 44720 37704
rect 44784 37640 44800 37704
rect 44864 37640 44880 37704
rect 44944 37640 44960 37704
rect 45024 37640 45040 37704
rect 45104 37640 45120 37704
rect 45184 37640 45200 37704
rect 45264 37640 45288 37704
rect 27889 37620 27955 37621
rect 27889 37556 27890 37620
rect 27954 37556 27955 37620
rect 27889 37555 27955 37556
rect 27892 37430 27952 37555
rect 27883 37414 27979 37430
rect 27883 37350 27899 37414
rect 27963 37350 27979 37414
rect 27883 37334 27979 37350
rect 27432 37303 27752 37322
rect 27164 37254 27260 37270
rect 27164 37190 27180 37254
rect 27244 37190 27260 37254
rect 27164 37174 27260 37190
rect 27164 37110 27180 37174
rect 27244 37110 27260 37174
rect 27164 37094 27260 37110
rect 27164 37030 27180 37094
rect 27244 37030 27260 37094
rect 27164 37014 27260 37030
rect 27164 36950 27180 37014
rect 27244 36950 27260 37014
rect 27423 37294 27752 37303
rect 27423 36990 27432 37294
rect 27736 36990 27752 37294
rect 27423 36981 27752 36990
rect 27164 36934 27260 36950
rect 27164 36870 27180 36934
rect 27244 36870 27260 36934
rect 27164 36854 27260 36870
rect 26445 36554 26541 36570
rect 26445 36490 26461 36554
rect 26525 36490 26541 36554
rect 26445 36474 26541 36490
rect 26445 36410 26461 36474
rect 26525 36410 26541 36474
rect 26445 36394 26541 36410
rect 26445 36330 26461 36394
rect 26525 36330 26541 36394
rect 26445 36314 26541 36330
rect 26445 36250 26461 36314
rect 26525 36250 26541 36314
rect 26704 36594 27032 36603
rect 26704 36290 26713 36594
rect 27017 36290 27032 36594
rect 26704 36281 27032 36290
rect 26445 36234 26541 36250
rect 26445 36170 26461 36234
rect 26525 36170 26541 36234
rect 26445 36154 26541 36170
rect 26712 36042 27032 36281
rect 27164 36714 27260 36730
rect 27164 36650 27180 36714
rect 27244 36650 27260 36714
rect 27164 36634 27260 36650
rect 27164 36570 27180 36634
rect 27244 36570 27260 36634
rect 27432 36603 27752 36981
rect 27883 37270 27899 37334
rect 27963 37270 27979 37334
rect 27883 37254 27979 37270
rect 27883 37190 27899 37254
rect 27963 37190 27979 37254
rect 27883 37174 27979 37190
rect 27883 37110 27899 37174
rect 27963 37110 27979 37174
rect 27883 37094 27979 37110
rect 27883 37030 27899 37094
rect 27963 37030 27979 37094
rect 27883 37014 27979 37030
rect 27883 36950 27899 37014
rect 27963 36950 27979 37014
rect 27883 36934 27979 36950
rect 27883 36870 27899 36934
rect 27963 36870 27979 36934
rect 27883 36854 27979 36870
rect 27164 36554 27260 36570
rect 27164 36490 27180 36554
rect 27244 36490 27260 36554
rect 27164 36474 27260 36490
rect 27164 36410 27180 36474
rect 27244 36410 27260 36474
rect 27164 36394 27260 36410
rect 27164 36330 27180 36394
rect 27244 36330 27260 36394
rect 27164 36314 27260 36330
rect 27164 36250 27180 36314
rect 27244 36250 27260 36314
rect 27423 36594 27752 36603
rect 27423 36290 27432 36594
rect 27736 36290 27752 36594
rect 27423 36281 27752 36290
rect 27164 36234 27260 36250
rect 27164 36170 27180 36234
rect 27244 36170 27260 36234
rect 27164 36154 27260 36170
rect 27432 36042 27752 36281
rect 27883 36714 27979 36730
rect 27883 36650 27899 36714
rect 27963 36650 27979 36714
rect 27883 36634 27979 36650
rect 27883 36570 27899 36634
rect 27963 36570 27979 36634
rect 27883 36554 27979 36570
rect 27883 36490 27899 36554
rect 27963 36490 27979 36554
rect 27883 36474 27979 36490
rect 27883 36410 27899 36474
rect 27963 36410 27979 36474
rect 27883 36394 27979 36410
rect 27883 36330 27899 36394
rect 27963 36330 27979 36394
rect 27883 36314 27979 36330
rect 27883 36250 27899 36314
rect 27963 36250 27979 36314
rect 27883 36234 27979 36250
rect 27883 36170 27899 36234
rect 27963 36170 27979 36234
rect 27883 36154 27979 36170
rect 5918 36032 13086 36042
rect 13366 36032 20534 36042
rect 5918 36014 20534 36032
rect 5918 35950 5946 36014
rect 6010 35950 6026 36014
rect 6090 35972 13394 36014
rect 6090 35950 13086 35972
rect 5918 35922 13086 35950
rect 13366 35950 13394 35972
rect 13458 35950 13474 36014
rect 13538 35950 20534 36014
rect 13366 35922 20534 35950
rect 20814 36014 27982 36042
rect 20814 35950 20842 36014
rect 20906 35950 20922 36014
rect 20986 35950 27982 36014
rect 20814 35922 27982 35950
rect 3348 33880 3372 33944
rect 3436 33880 3452 33944
rect 3516 33880 3532 33944
rect 3596 33880 3612 33944
rect 3676 33880 3692 33944
rect 3756 33880 3772 33944
rect 3836 33880 3852 33944
rect 3916 33880 3932 33944
rect 3996 33880 4012 33944
rect 4076 33880 4092 33944
rect 4156 33880 4172 33944
rect 4236 33880 4252 33944
rect 4316 33880 4332 33944
rect 4396 33880 4412 33944
rect 4476 33880 4492 33944
rect 4556 33880 4572 33944
rect 4636 33880 4652 33944
rect 4716 33880 4732 33944
rect 4796 33880 4812 33944
rect 4876 33880 4892 33944
rect 4956 33880 4980 33944
rect 3348 30184 4980 33880
rect 10087 33838 10153 33839
rect 10087 33774 10088 33838
rect 10152 33774 10153 33838
rect 10087 33773 10153 33774
rect 10090 33670 10150 33773
rect 7202 33654 7298 33670
rect 7202 33590 7218 33654
rect 7282 33590 7298 33654
rect 7202 33574 7298 33590
rect 6742 33543 7062 33562
rect 6742 33534 7064 33543
rect 6742 33230 6751 33534
rect 7055 33230 7064 33534
rect 6742 33221 7064 33230
rect 7202 33510 7218 33574
rect 7282 33510 7298 33574
rect 7921 33654 8017 33670
rect 7921 33590 7937 33654
rect 8001 33590 8017 33654
rect 7921 33574 8017 33590
rect 7462 33543 7782 33562
rect 7202 33494 7298 33510
rect 7202 33430 7218 33494
rect 7282 33430 7298 33494
rect 7202 33414 7298 33430
rect 7202 33350 7218 33414
rect 7282 33350 7298 33414
rect 7202 33334 7298 33350
rect 7202 33270 7218 33334
rect 7282 33270 7298 33334
rect 7202 33254 7298 33270
rect 6742 32843 7062 33221
rect 7202 33190 7218 33254
rect 7282 33190 7298 33254
rect 7461 33534 7783 33543
rect 7461 33230 7470 33534
rect 7774 33230 7783 33534
rect 7461 33221 7783 33230
rect 7921 33510 7937 33574
rect 8001 33510 8017 33574
rect 8640 33654 8736 33670
rect 8640 33590 8656 33654
rect 8720 33590 8736 33654
rect 8640 33574 8736 33590
rect 8182 33543 8502 33562
rect 7921 33494 8017 33510
rect 7921 33430 7937 33494
rect 8001 33430 8017 33494
rect 7921 33414 8017 33430
rect 7921 33350 7937 33414
rect 8001 33350 8017 33414
rect 7921 33334 8017 33350
rect 7921 33270 7937 33334
rect 8001 33270 8017 33334
rect 7921 33254 8017 33270
rect 7202 33174 7298 33190
rect 7202 33110 7218 33174
rect 7282 33110 7298 33174
rect 7202 33094 7298 33110
rect 7202 32954 7298 32970
rect 7202 32890 7218 32954
rect 7282 32890 7298 32954
rect 7202 32874 7298 32890
rect 6742 32834 7064 32843
rect 6742 32530 6751 32834
rect 7055 32530 7064 32834
rect 6742 32521 7064 32530
rect 7202 32810 7218 32874
rect 7282 32810 7298 32874
rect 7462 32843 7782 33221
rect 7921 33190 7937 33254
rect 8001 33190 8017 33254
rect 8180 33534 8502 33543
rect 8180 33230 8189 33534
rect 8493 33230 8502 33534
rect 8180 33221 8502 33230
rect 7921 33174 8017 33190
rect 7921 33110 7937 33174
rect 8001 33110 8017 33174
rect 7921 33094 8017 33110
rect 7921 32954 8017 32970
rect 7921 32890 7937 32954
rect 8001 32890 8017 32954
rect 7921 32874 8017 32890
rect 7202 32794 7298 32810
rect 7202 32730 7218 32794
rect 7282 32730 7298 32794
rect 7202 32714 7298 32730
rect 7202 32650 7218 32714
rect 7282 32650 7298 32714
rect 7202 32634 7298 32650
rect 7202 32570 7218 32634
rect 7282 32570 7298 32634
rect 7202 32554 7298 32570
rect 6742 32282 7062 32521
rect 7202 32490 7218 32554
rect 7282 32490 7298 32554
rect 7461 32834 7783 32843
rect 7461 32530 7470 32834
rect 7774 32530 7783 32834
rect 7461 32521 7783 32530
rect 7921 32810 7937 32874
rect 8001 32810 8017 32874
rect 8182 32843 8502 33221
rect 8640 33510 8656 33574
rect 8720 33510 8736 33574
rect 9359 33654 9455 33670
rect 9359 33590 9375 33654
rect 9439 33590 9455 33654
rect 9359 33574 9455 33590
rect 8902 33543 9222 33562
rect 8640 33494 8736 33510
rect 8640 33430 8656 33494
rect 8720 33430 8736 33494
rect 8640 33414 8736 33430
rect 8640 33350 8656 33414
rect 8720 33350 8736 33414
rect 8640 33334 8736 33350
rect 8640 33270 8656 33334
rect 8720 33270 8736 33334
rect 8640 33254 8736 33270
rect 8640 33190 8656 33254
rect 8720 33190 8736 33254
rect 8899 33534 9222 33543
rect 8899 33230 8908 33534
rect 9212 33230 9222 33534
rect 8899 33221 9222 33230
rect 8640 33174 8736 33190
rect 8640 33110 8656 33174
rect 8720 33110 8736 33174
rect 8640 33094 8736 33110
rect 7921 32794 8017 32810
rect 7921 32730 7937 32794
rect 8001 32730 8017 32794
rect 7921 32714 8017 32730
rect 7921 32650 7937 32714
rect 8001 32650 8017 32714
rect 7921 32634 8017 32650
rect 7921 32570 7937 32634
rect 8001 32570 8017 32634
rect 7921 32554 8017 32570
rect 7202 32474 7298 32490
rect 7202 32410 7218 32474
rect 7282 32410 7298 32474
rect 7202 32394 7298 32410
rect 7462 32282 7782 32521
rect 7921 32490 7937 32554
rect 8001 32490 8017 32554
rect 8180 32834 8502 32843
rect 8180 32530 8189 32834
rect 8493 32530 8502 32834
rect 8180 32521 8502 32530
rect 7921 32474 8017 32490
rect 7921 32410 7937 32474
rect 8001 32410 8017 32474
rect 7921 32394 8017 32410
rect 8182 32282 8502 32521
rect 8640 32954 8736 32970
rect 8640 32890 8656 32954
rect 8720 32890 8736 32954
rect 8640 32874 8736 32890
rect 8640 32810 8656 32874
rect 8720 32810 8736 32874
rect 8902 32843 9222 33221
rect 9359 33510 9375 33574
rect 9439 33510 9455 33574
rect 10078 33654 10174 33670
rect 10078 33590 10094 33654
rect 10158 33590 10174 33654
rect 10078 33574 10174 33590
rect 9622 33543 9942 33562
rect 9359 33494 9455 33510
rect 9359 33430 9375 33494
rect 9439 33430 9455 33494
rect 9359 33414 9455 33430
rect 9359 33350 9375 33414
rect 9439 33350 9455 33414
rect 9359 33334 9455 33350
rect 9359 33270 9375 33334
rect 9439 33270 9455 33334
rect 9359 33254 9455 33270
rect 9359 33190 9375 33254
rect 9439 33190 9455 33254
rect 9618 33534 9942 33543
rect 9618 33230 9627 33534
rect 9931 33230 9942 33534
rect 9618 33221 9942 33230
rect 9359 33174 9455 33190
rect 9359 33110 9375 33174
rect 9439 33110 9455 33174
rect 9359 33094 9455 33110
rect 8640 32794 8736 32810
rect 8640 32730 8656 32794
rect 8720 32730 8736 32794
rect 8640 32714 8736 32730
rect 8640 32650 8656 32714
rect 8720 32650 8736 32714
rect 8640 32634 8736 32650
rect 8640 32570 8656 32634
rect 8720 32570 8736 32634
rect 8640 32554 8736 32570
rect 8640 32490 8656 32554
rect 8720 32490 8736 32554
rect 8899 32834 9222 32843
rect 8899 32530 8908 32834
rect 9212 32530 9222 32834
rect 8899 32521 9222 32530
rect 8640 32474 8736 32490
rect 8640 32410 8656 32474
rect 8720 32410 8736 32474
rect 8640 32394 8736 32410
rect 8902 32282 9222 32521
rect 9359 32954 9455 32970
rect 9359 32890 9375 32954
rect 9439 32890 9455 32954
rect 9359 32874 9455 32890
rect 9359 32810 9375 32874
rect 9439 32810 9455 32874
rect 9622 32843 9942 33221
rect 10078 33510 10094 33574
rect 10158 33510 10174 33574
rect 10797 33654 10893 33670
rect 10797 33590 10813 33654
rect 10877 33590 10893 33654
rect 10797 33574 10893 33590
rect 10342 33543 10662 33562
rect 10078 33494 10174 33510
rect 10078 33430 10094 33494
rect 10158 33430 10174 33494
rect 10078 33414 10174 33430
rect 10078 33350 10094 33414
rect 10158 33350 10174 33414
rect 10078 33334 10174 33350
rect 10078 33270 10094 33334
rect 10158 33270 10174 33334
rect 10078 33254 10174 33270
rect 10078 33190 10094 33254
rect 10158 33190 10174 33254
rect 10337 33534 10662 33543
rect 10337 33230 10346 33534
rect 10650 33230 10662 33534
rect 10337 33221 10662 33230
rect 10078 33174 10174 33190
rect 10078 33110 10094 33174
rect 10158 33110 10174 33174
rect 10078 33094 10174 33110
rect 9359 32794 9455 32810
rect 9359 32730 9375 32794
rect 9439 32730 9455 32794
rect 9359 32714 9455 32730
rect 9359 32650 9375 32714
rect 9439 32650 9455 32714
rect 9359 32634 9455 32650
rect 9359 32570 9375 32634
rect 9439 32570 9455 32634
rect 9359 32554 9455 32570
rect 9359 32490 9375 32554
rect 9439 32490 9455 32554
rect 9618 32834 9942 32843
rect 9618 32530 9627 32834
rect 9931 32530 9942 32834
rect 9618 32521 9942 32530
rect 9359 32474 9455 32490
rect 9359 32410 9375 32474
rect 9439 32410 9455 32474
rect 9359 32394 9455 32410
rect 9622 32282 9942 32521
rect 10078 32954 10174 32970
rect 10078 32890 10094 32954
rect 10158 32890 10174 32954
rect 10078 32874 10174 32890
rect 10078 32810 10094 32874
rect 10158 32810 10174 32874
rect 10342 32843 10662 33221
rect 10797 33510 10813 33574
rect 10877 33510 10893 33574
rect 11516 33654 11612 33670
rect 11516 33590 11532 33654
rect 11596 33590 11612 33654
rect 11516 33574 11612 33590
rect 11062 33543 11382 33562
rect 10797 33494 10893 33510
rect 10797 33430 10813 33494
rect 10877 33430 10893 33494
rect 10797 33414 10893 33430
rect 10797 33350 10813 33414
rect 10877 33350 10893 33414
rect 10797 33334 10893 33350
rect 10797 33270 10813 33334
rect 10877 33270 10893 33334
rect 10797 33254 10893 33270
rect 10797 33190 10813 33254
rect 10877 33190 10893 33254
rect 11056 33534 11382 33543
rect 11056 33230 11065 33534
rect 11369 33230 11382 33534
rect 11056 33221 11382 33230
rect 10797 33174 10893 33190
rect 10797 33110 10813 33174
rect 10877 33110 10893 33174
rect 10797 33094 10893 33110
rect 10078 32794 10174 32810
rect 10078 32730 10094 32794
rect 10158 32730 10174 32794
rect 10078 32714 10174 32730
rect 10078 32650 10094 32714
rect 10158 32650 10174 32714
rect 10078 32634 10174 32650
rect 10078 32570 10094 32634
rect 10158 32570 10174 32634
rect 10078 32554 10174 32570
rect 10078 32490 10094 32554
rect 10158 32490 10174 32554
rect 10337 32834 10662 32843
rect 10337 32530 10346 32834
rect 10650 32530 10662 32834
rect 10337 32521 10662 32530
rect 10078 32474 10174 32490
rect 10078 32410 10094 32474
rect 10158 32410 10174 32474
rect 10078 32394 10174 32410
rect 10342 32282 10662 32521
rect 10797 32954 10893 32970
rect 10797 32890 10813 32954
rect 10877 32890 10893 32954
rect 10797 32874 10893 32890
rect 10797 32810 10813 32874
rect 10877 32810 10893 32874
rect 11062 32843 11382 33221
rect 11516 33510 11532 33574
rect 11596 33510 11612 33574
rect 12235 33654 12331 33670
rect 12235 33590 12251 33654
rect 12315 33590 12331 33654
rect 12235 33574 12331 33590
rect 11782 33543 12102 33562
rect 11516 33494 11612 33510
rect 11516 33430 11532 33494
rect 11596 33430 11612 33494
rect 11516 33414 11612 33430
rect 11516 33350 11532 33414
rect 11596 33350 11612 33414
rect 11516 33334 11612 33350
rect 11516 33270 11532 33334
rect 11596 33270 11612 33334
rect 11516 33254 11612 33270
rect 11516 33190 11532 33254
rect 11596 33190 11612 33254
rect 11775 33534 12102 33543
rect 11775 33230 11784 33534
rect 12088 33230 12102 33534
rect 11775 33221 12102 33230
rect 11516 33174 11612 33190
rect 11516 33110 11532 33174
rect 11596 33110 11612 33174
rect 11516 33094 11612 33110
rect 10797 32794 10893 32810
rect 10797 32730 10813 32794
rect 10877 32730 10893 32794
rect 10797 32714 10893 32730
rect 10797 32650 10813 32714
rect 10877 32650 10893 32714
rect 10797 32634 10893 32650
rect 10797 32570 10813 32634
rect 10877 32570 10893 32634
rect 10797 32554 10893 32570
rect 10797 32490 10813 32554
rect 10877 32490 10893 32554
rect 11056 32834 11382 32843
rect 11056 32530 11065 32834
rect 11369 32530 11382 32834
rect 11056 32521 11382 32530
rect 10797 32474 10893 32490
rect 10797 32410 10813 32474
rect 10877 32410 10893 32474
rect 10797 32394 10893 32410
rect 11062 32282 11382 32521
rect 11516 32954 11612 32970
rect 11516 32890 11532 32954
rect 11596 32890 11612 32954
rect 11516 32874 11612 32890
rect 11516 32810 11532 32874
rect 11596 32810 11612 32874
rect 11782 32843 12102 33221
rect 12235 33510 12251 33574
rect 12315 33510 12331 33574
rect 12954 33654 13050 33670
rect 12954 33590 12970 33654
rect 13034 33590 13050 33654
rect 12954 33574 13050 33590
rect 12502 33543 12822 33562
rect 12235 33494 12331 33510
rect 12235 33430 12251 33494
rect 12315 33430 12331 33494
rect 12235 33414 12331 33430
rect 12235 33350 12251 33414
rect 12315 33350 12331 33414
rect 12235 33334 12331 33350
rect 12235 33270 12251 33334
rect 12315 33270 12331 33334
rect 12235 33254 12331 33270
rect 12235 33190 12251 33254
rect 12315 33190 12331 33254
rect 12494 33534 12822 33543
rect 12494 33230 12503 33534
rect 12807 33230 12822 33534
rect 12494 33221 12822 33230
rect 12235 33174 12331 33190
rect 12235 33110 12251 33174
rect 12315 33110 12331 33174
rect 12235 33094 12331 33110
rect 11516 32794 11612 32810
rect 11516 32730 11532 32794
rect 11596 32730 11612 32794
rect 11516 32714 11612 32730
rect 11516 32650 11532 32714
rect 11596 32650 11612 32714
rect 11516 32634 11612 32650
rect 11516 32570 11532 32634
rect 11596 32570 11612 32634
rect 11516 32554 11612 32570
rect 11516 32490 11532 32554
rect 11596 32490 11612 32554
rect 11775 32834 12102 32843
rect 11775 32530 11784 32834
rect 12088 32530 12102 32834
rect 11775 32521 12102 32530
rect 11516 32474 11612 32490
rect 11516 32410 11532 32474
rect 11596 32410 11612 32474
rect 11516 32394 11612 32410
rect 11782 32282 12102 32521
rect 12235 32954 12331 32970
rect 12235 32890 12251 32954
rect 12315 32890 12331 32954
rect 12235 32874 12331 32890
rect 12235 32810 12251 32874
rect 12315 32810 12331 32874
rect 12502 32843 12822 33221
rect 12954 33510 12970 33574
rect 13034 33510 13050 33574
rect 13402 33562 13462 35922
rect 43656 33944 45288 37640
rect 43656 33880 43680 33944
rect 43744 33880 43760 33944
rect 43824 33880 43840 33944
rect 43904 33880 43920 33944
rect 43984 33880 44000 33944
rect 44064 33880 44080 33944
rect 44144 33880 44160 33944
rect 44224 33880 44240 33944
rect 44304 33880 44320 33944
rect 44384 33880 44400 33944
rect 44464 33880 44480 33944
rect 44544 33880 44560 33944
rect 44624 33880 44640 33944
rect 44704 33880 44720 33944
rect 44784 33880 44800 33944
rect 44864 33880 44880 33944
rect 44944 33880 44960 33944
rect 45024 33880 45040 33944
rect 45104 33880 45120 33944
rect 45184 33880 45200 33944
rect 45264 33880 45288 33944
rect 13673 33654 13769 33670
rect 13673 33590 13689 33654
rect 13753 33590 13769 33654
rect 13673 33574 13769 33590
rect 13222 33543 13542 33562
rect 12954 33494 13050 33510
rect 12954 33430 12970 33494
rect 13034 33430 13050 33494
rect 12954 33414 13050 33430
rect 12954 33350 12970 33414
rect 13034 33350 13050 33414
rect 12954 33334 13050 33350
rect 12954 33270 12970 33334
rect 13034 33270 13050 33334
rect 12954 33254 13050 33270
rect 12954 33190 12970 33254
rect 13034 33190 13050 33254
rect 13213 33534 13542 33543
rect 13213 33230 13222 33534
rect 13526 33230 13542 33534
rect 13213 33221 13542 33230
rect 12954 33174 13050 33190
rect 12954 33110 12970 33174
rect 13034 33110 13050 33174
rect 12954 33094 13050 33110
rect 12235 32794 12331 32810
rect 12235 32730 12251 32794
rect 12315 32730 12331 32794
rect 12235 32714 12331 32730
rect 12235 32650 12251 32714
rect 12315 32650 12331 32714
rect 12235 32634 12331 32650
rect 12235 32570 12251 32634
rect 12315 32570 12331 32634
rect 12235 32554 12331 32570
rect 12235 32490 12251 32554
rect 12315 32490 12331 32554
rect 12494 32834 12822 32843
rect 12494 32530 12503 32834
rect 12807 32530 12822 32834
rect 12494 32521 12822 32530
rect 12235 32474 12331 32490
rect 12235 32410 12251 32474
rect 12315 32410 12331 32474
rect 12235 32394 12331 32410
rect 12502 32282 12822 32521
rect 12954 32954 13050 32970
rect 12954 32890 12970 32954
rect 13034 32890 13050 32954
rect 12954 32874 13050 32890
rect 12954 32810 12970 32874
rect 13034 32810 13050 32874
rect 13222 32843 13542 33221
rect 13673 33510 13689 33574
rect 13753 33510 13769 33574
rect 13673 33494 13769 33510
rect 13673 33430 13689 33494
rect 13753 33430 13769 33494
rect 13673 33414 13769 33430
rect 13673 33350 13689 33414
rect 13753 33350 13769 33414
rect 13673 33334 13769 33350
rect 13673 33270 13689 33334
rect 13753 33270 13769 33334
rect 13673 33254 13769 33270
rect 13673 33190 13689 33254
rect 13753 33190 13769 33254
rect 13673 33174 13769 33190
rect 13673 33110 13689 33174
rect 13753 33110 13769 33174
rect 13673 33094 13769 33110
rect 12954 32794 13050 32810
rect 12954 32730 12970 32794
rect 13034 32730 13050 32794
rect 12954 32714 13050 32730
rect 12954 32650 12970 32714
rect 13034 32650 13050 32714
rect 12954 32634 13050 32650
rect 12954 32570 12970 32634
rect 13034 32570 13050 32634
rect 12954 32554 13050 32570
rect 12954 32490 12970 32554
rect 13034 32490 13050 32554
rect 13213 32834 13542 32843
rect 13213 32530 13222 32834
rect 13526 32530 13542 32834
rect 13213 32521 13542 32530
rect 12954 32474 13050 32490
rect 12954 32410 12970 32474
rect 13034 32410 13050 32474
rect 12954 32394 13050 32410
rect 13222 32282 13542 32521
rect 13673 32954 13769 32970
rect 13673 32890 13689 32954
rect 13753 32890 13769 32954
rect 13673 32874 13769 32890
rect 13673 32810 13689 32874
rect 13753 32810 13769 32874
rect 13673 32794 13769 32810
rect 13673 32730 13689 32794
rect 13753 32730 13769 32794
rect 13673 32714 13769 32730
rect 13673 32650 13689 32714
rect 13753 32650 13769 32714
rect 13673 32634 13769 32650
rect 13673 32570 13689 32634
rect 13753 32570 13769 32634
rect 13673 32554 13769 32570
rect 13673 32490 13689 32554
rect 13753 32490 13769 32554
rect 13673 32474 13769 32490
rect 13673 32410 13689 32474
rect 13753 32410 13769 32474
rect 13673 32394 13769 32410
rect 6604 32254 13772 32282
rect 6604 32190 6632 32254
rect 6696 32190 6712 32254
rect 6776 32252 13772 32254
rect 6776 32190 13538 32252
rect 6604 32188 13538 32190
rect 13602 32188 13772 32252
rect 6604 32162 13772 32188
rect 3348 30120 3372 30184
rect 3436 30120 3452 30184
rect 3516 30120 3532 30184
rect 3596 30120 3612 30184
rect 3676 30120 3692 30184
rect 3756 30120 3772 30184
rect 3836 30120 3852 30184
rect 3916 30120 3932 30184
rect 3996 30120 4012 30184
rect 4076 30120 4092 30184
rect 4156 30120 4172 30184
rect 4236 30120 4252 30184
rect 4316 30120 4332 30184
rect 4396 30120 4412 30184
rect 4476 30120 4492 30184
rect 4556 30120 4572 30184
rect 4636 30120 4652 30184
rect 4716 30120 4732 30184
rect 4796 30120 4812 30184
rect 4876 30120 4892 30184
rect 4956 30120 4980 30184
rect 3348 26424 4980 30120
rect 43656 30184 45288 33880
rect 43656 30120 43680 30184
rect 43744 30120 43760 30184
rect 43824 30120 43840 30184
rect 43904 30120 43920 30184
rect 43984 30120 44000 30184
rect 44064 30120 44080 30184
rect 44144 30120 44160 30184
rect 44224 30120 44240 30184
rect 44304 30120 44320 30184
rect 44384 30120 44400 30184
rect 44464 30120 44480 30184
rect 44544 30120 44560 30184
rect 44624 30120 44640 30184
rect 44704 30120 44720 30184
rect 44784 30120 44800 30184
rect 44864 30120 44880 30184
rect 44944 30120 44960 30184
rect 45024 30120 45040 30184
rect 45104 30120 45120 30184
rect 45184 30120 45200 30184
rect 45264 30120 45288 30184
rect 18919 28592 18985 28593
rect 18919 28528 18920 28592
rect 18984 28528 18985 28592
rect 18919 28527 18985 28528
rect 3348 26360 3372 26424
rect 3436 26360 3452 26424
rect 3516 26360 3532 26424
rect 3596 26360 3612 26424
rect 3676 26360 3692 26424
rect 3756 26360 3772 26424
rect 3836 26360 3852 26424
rect 3916 26360 3932 26424
rect 3996 26360 4012 26424
rect 4076 26360 4092 26424
rect 4156 26360 4172 26424
rect 4236 26360 4252 26424
rect 4316 26360 4332 26424
rect 4396 26360 4412 26424
rect 4476 26360 4492 26424
rect 4556 26360 4572 26424
rect 4636 26360 4652 26424
rect 4716 26360 4732 26424
rect 4796 26360 4812 26424
rect 4876 26360 4892 26424
rect 4956 26360 4980 26424
rect 3348 22664 4980 26360
rect 18922 26150 18982 28527
rect 43656 26424 45288 30120
rect 43656 26360 43680 26424
rect 43744 26360 43760 26424
rect 43824 26360 43840 26424
rect 43904 26360 43920 26424
rect 43984 26360 44000 26424
rect 44064 26360 44080 26424
rect 44144 26360 44160 26424
rect 44224 26360 44240 26424
rect 44304 26360 44320 26424
rect 44384 26360 44400 26424
rect 44464 26360 44480 26424
rect 44544 26360 44560 26424
rect 44624 26360 44640 26424
rect 44704 26360 44720 26424
rect 44784 26360 44800 26424
rect 44864 26360 44880 26424
rect 44944 26360 44960 26424
rect 45024 26360 45040 26424
rect 45104 26360 45120 26424
rect 45184 26360 45200 26424
rect 45264 26360 45288 26424
rect 16022 26134 16118 26150
rect 16022 26070 16038 26134
rect 16102 26070 16118 26134
rect 16022 26054 16118 26070
rect 15562 26023 15882 26042
rect 15562 26014 15884 26023
rect 15562 25710 15571 26014
rect 15875 25710 15884 26014
rect 15562 25701 15884 25710
rect 16022 25990 16038 26054
rect 16102 25990 16118 26054
rect 16741 26134 16837 26150
rect 16741 26070 16757 26134
rect 16821 26070 16837 26134
rect 16741 26054 16837 26070
rect 16282 26023 16602 26042
rect 16022 25974 16118 25990
rect 16022 25910 16038 25974
rect 16102 25910 16118 25974
rect 16022 25894 16118 25910
rect 16022 25830 16038 25894
rect 16102 25830 16118 25894
rect 16022 25814 16118 25830
rect 16022 25750 16038 25814
rect 16102 25750 16118 25814
rect 16022 25734 16118 25750
rect 15562 25323 15882 25701
rect 16022 25670 16038 25734
rect 16102 25670 16118 25734
rect 16281 26014 16603 26023
rect 16281 25710 16290 26014
rect 16594 25710 16603 26014
rect 16281 25701 16603 25710
rect 16741 25990 16757 26054
rect 16821 25990 16837 26054
rect 17460 26134 17556 26150
rect 17460 26070 17476 26134
rect 17540 26070 17556 26134
rect 17460 26054 17556 26070
rect 17002 26023 17322 26042
rect 16741 25974 16837 25990
rect 16741 25910 16757 25974
rect 16821 25910 16837 25974
rect 16741 25894 16837 25910
rect 16741 25830 16757 25894
rect 16821 25830 16837 25894
rect 16741 25814 16837 25830
rect 16741 25750 16757 25814
rect 16821 25750 16837 25814
rect 16741 25734 16837 25750
rect 16022 25654 16118 25670
rect 16022 25590 16038 25654
rect 16102 25590 16118 25654
rect 16022 25574 16118 25590
rect 16022 25434 16118 25450
rect 16022 25370 16038 25434
rect 16102 25370 16118 25434
rect 16022 25354 16118 25370
rect 15562 25314 15884 25323
rect 15562 25010 15571 25314
rect 15875 25010 15884 25314
rect 15562 25001 15884 25010
rect 16022 25290 16038 25354
rect 16102 25290 16118 25354
rect 16282 25323 16602 25701
rect 16741 25670 16757 25734
rect 16821 25670 16837 25734
rect 17000 26014 17322 26023
rect 17000 25710 17009 26014
rect 17313 25710 17322 26014
rect 17000 25701 17322 25710
rect 16741 25654 16837 25670
rect 16741 25590 16757 25654
rect 16821 25590 16837 25654
rect 16741 25574 16837 25590
rect 16741 25434 16837 25450
rect 16741 25370 16757 25434
rect 16821 25370 16837 25434
rect 16741 25354 16837 25370
rect 16022 25274 16118 25290
rect 16022 25210 16038 25274
rect 16102 25210 16118 25274
rect 16022 25194 16118 25210
rect 16022 25130 16038 25194
rect 16102 25130 16118 25194
rect 16022 25114 16118 25130
rect 16022 25050 16038 25114
rect 16102 25050 16118 25114
rect 16022 25034 16118 25050
rect 15562 24762 15882 25001
rect 16022 24970 16038 25034
rect 16102 24970 16118 25034
rect 16281 25314 16603 25323
rect 16281 25010 16290 25314
rect 16594 25010 16603 25314
rect 16281 25001 16603 25010
rect 16741 25290 16757 25354
rect 16821 25290 16837 25354
rect 17002 25323 17322 25701
rect 17460 25990 17476 26054
rect 17540 25990 17556 26054
rect 18179 26134 18275 26150
rect 18179 26070 18195 26134
rect 18259 26070 18275 26134
rect 18179 26054 18275 26070
rect 17722 26023 18042 26042
rect 17460 25974 17556 25990
rect 17460 25910 17476 25974
rect 17540 25910 17556 25974
rect 17460 25894 17556 25910
rect 17460 25830 17476 25894
rect 17540 25830 17556 25894
rect 17460 25814 17556 25830
rect 17460 25750 17476 25814
rect 17540 25750 17556 25814
rect 17460 25734 17556 25750
rect 17460 25670 17476 25734
rect 17540 25670 17556 25734
rect 17719 26014 18042 26023
rect 17719 25710 17728 26014
rect 18032 25710 18042 26014
rect 17719 25701 18042 25710
rect 17460 25654 17556 25670
rect 17460 25590 17476 25654
rect 17540 25590 17556 25654
rect 17460 25574 17556 25590
rect 16741 25274 16837 25290
rect 16741 25210 16757 25274
rect 16821 25210 16837 25274
rect 16741 25194 16837 25210
rect 16741 25130 16757 25194
rect 16821 25130 16837 25194
rect 16741 25114 16837 25130
rect 16741 25050 16757 25114
rect 16821 25050 16837 25114
rect 16741 25034 16837 25050
rect 16022 24954 16118 24970
rect 16022 24890 16038 24954
rect 16102 24890 16118 24954
rect 16022 24874 16118 24890
rect 16282 24762 16602 25001
rect 16741 24970 16757 25034
rect 16821 24970 16837 25034
rect 17000 25314 17322 25323
rect 17000 25010 17009 25314
rect 17313 25010 17322 25314
rect 17000 25001 17322 25010
rect 16741 24954 16837 24970
rect 16741 24890 16757 24954
rect 16821 24890 16837 24954
rect 16741 24874 16837 24890
rect 17002 24762 17322 25001
rect 17460 25434 17556 25450
rect 17460 25370 17476 25434
rect 17540 25370 17556 25434
rect 17460 25354 17556 25370
rect 17460 25290 17476 25354
rect 17540 25290 17556 25354
rect 17722 25323 18042 25701
rect 18179 25990 18195 26054
rect 18259 25990 18275 26054
rect 18898 26134 18994 26150
rect 18898 26070 18914 26134
rect 18978 26070 18994 26134
rect 18898 26054 18994 26070
rect 18442 26023 18762 26042
rect 18179 25974 18275 25990
rect 18179 25910 18195 25974
rect 18259 25910 18275 25974
rect 18179 25894 18275 25910
rect 18179 25830 18195 25894
rect 18259 25830 18275 25894
rect 18179 25814 18275 25830
rect 18179 25750 18195 25814
rect 18259 25750 18275 25814
rect 18179 25734 18275 25750
rect 18179 25670 18195 25734
rect 18259 25670 18275 25734
rect 18438 26014 18762 26023
rect 18438 25710 18447 26014
rect 18751 25710 18762 26014
rect 18438 25701 18762 25710
rect 18179 25654 18275 25670
rect 18179 25590 18195 25654
rect 18259 25590 18275 25654
rect 18179 25574 18275 25590
rect 17460 25274 17556 25290
rect 17460 25210 17476 25274
rect 17540 25210 17556 25274
rect 17460 25194 17556 25210
rect 17460 25130 17476 25194
rect 17540 25130 17556 25194
rect 17460 25114 17556 25130
rect 17460 25050 17476 25114
rect 17540 25050 17556 25114
rect 17460 25034 17556 25050
rect 17460 24970 17476 25034
rect 17540 24970 17556 25034
rect 17719 25314 18042 25323
rect 17719 25010 17728 25314
rect 18032 25010 18042 25314
rect 17719 25001 18042 25010
rect 17460 24954 17556 24970
rect 17460 24890 17476 24954
rect 17540 24890 17556 24954
rect 17460 24874 17556 24890
rect 17722 24762 18042 25001
rect 18179 25434 18275 25450
rect 18179 25370 18195 25434
rect 18259 25370 18275 25434
rect 18179 25354 18275 25370
rect 18179 25290 18195 25354
rect 18259 25290 18275 25354
rect 18442 25323 18762 25701
rect 18898 25990 18914 26054
rect 18978 25990 18994 26054
rect 19617 26134 19713 26150
rect 19617 26070 19633 26134
rect 19697 26070 19713 26134
rect 19617 26054 19713 26070
rect 19162 26023 19482 26042
rect 18898 25974 18994 25990
rect 18898 25910 18914 25974
rect 18978 25910 18994 25974
rect 18898 25894 18994 25910
rect 18898 25830 18914 25894
rect 18978 25830 18994 25894
rect 18898 25814 18994 25830
rect 18898 25750 18914 25814
rect 18978 25750 18994 25814
rect 18898 25734 18994 25750
rect 18898 25670 18914 25734
rect 18978 25670 18994 25734
rect 19157 26014 19482 26023
rect 19157 25710 19166 26014
rect 19470 25710 19482 26014
rect 19157 25701 19482 25710
rect 18898 25654 18994 25670
rect 18898 25590 18914 25654
rect 18978 25590 18994 25654
rect 18898 25574 18994 25590
rect 18179 25274 18275 25290
rect 18179 25210 18195 25274
rect 18259 25210 18275 25274
rect 18179 25194 18275 25210
rect 18179 25130 18195 25194
rect 18259 25130 18275 25194
rect 18179 25114 18275 25130
rect 18179 25050 18195 25114
rect 18259 25050 18275 25114
rect 18179 25034 18275 25050
rect 18179 24970 18195 25034
rect 18259 24970 18275 25034
rect 18438 25314 18762 25323
rect 18438 25010 18447 25314
rect 18751 25010 18762 25314
rect 18438 25001 18762 25010
rect 18179 24954 18275 24970
rect 18179 24890 18195 24954
rect 18259 24890 18275 24954
rect 18179 24874 18275 24890
rect 18442 24762 18762 25001
rect 18898 25434 18994 25450
rect 18898 25370 18914 25434
rect 18978 25370 18994 25434
rect 18898 25354 18994 25370
rect 18898 25290 18914 25354
rect 18978 25290 18994 25354
rect 19162 25323 19482 25701
rect 19617 25990 19633 26054
rect 19697 25990 19713 26054
rect 20336 26134 20432 26150
rect 20336 26070 20352 26134
rect 20416 26070 20432 26134
rect 20336 26054 20432 26070
rect 19882 26023 20202 26042
rect 19617 25974 19713 25990
rect 19617 25910 19633 25974
rect 19697 25910 19713 25974
rect 19617 25894 19713 25910
rect 19617 25830 19633 25894
rect 19697 25830 19713 25894
rect 19617 25814 19713 25830
rect 19617 25750 19633 25814
rect 19697 25750 19713 25814
rect 19617 25734 19713 25750
rect 19617 25670 19633 25734
rect 19697 25670 19713 25734
rect 19876 26014 20202 26023
rect 19876 25710 19885 26014
rect 20189 25710 20202 26014
rect 19876 25701 20202 25710
rect 19617 25654 19713 25670
rect 19617 25590 19633 25654
rect 19697 25590 19713 25654
rect 19617 25574 19713 25590
rect 18898 25274 18994 25290
rect 18898 25210 18914 25274
rect 18978 25210 18994 25274
rect 18898 25194 18994 25210
rect 18898 25130 18914 25194
rect 18978 25130 18994 25194
rect 18898 25114 18994 25130
rect 18898 25050 18914 25114
rect 18978 25050 18994 25114
rect 18898 25034 18994 25050
rect 18898 24970 18914 25034
rect 18978 24970 18994 25034
rect 19157 25314 19482 25323
rect 19157 25010 19166 25314
rect 19470 25010 19482 25314
rect 19157 25001 19482 25010
rect 18898 24954 18994 24970
rect 18898 24890 18914 24954
rect 18978 24890 18994 24954
rect 18898 24874 18994 24890
rect 19162 24762 19482 25001
rect 19617 25434 19713 25450
rect 19617 25370 19633 25434
rect 19697 25370 19713 25434
rect 19617 25354 19713 25370
rect 19617 25290 19633 25354
rect 19697 25290 19713 25354
rect 19882 25323 20202 25701
rect 20336 25990 20352 26054
rect 20416 25990 20432 26054
rect 21055 26134 21151 26150
rect 21055 26070 21071 26134
rect 21135 26070 21151 26134
rect 21055 26054 21151 26070
rect 20602 26023 20922 26042
rect 20336 25974 20432 25990
rect 20336 25910 20352 25974
rect 20416 25910 20432 25974
rect 20336 25894 20432 25910
rect 20336 25830 20352 25894
rect 20416 25830 20432 25894
rect 20336 25814 20432 25830
rect 20336 25750 20352 25814
rect 20416 25750 20432 25814
rect 20336 25734 20432 25750
rect 20336 25670 20352 25734
rect 20416 25670 20432 25734
rect 20595 26014 20922 26023
rect 20595 25710 20604 26014
rect 20908 25710 20922 26014
rect 20595 25701 20922 25710
rect 20336 25654 20432 25670
rect 20336 25590 20352 25654
rect 20416 25590 20432 25654
rect 20336 25574 20432 25590
rect 19617 25274 19713 25290
rect 19617 25210 19633 25274
rect 19697 25210 19713 25274
rect 19617 25194 19713 25210
rect 19617 25130 19633 25194
rect 19697 25130 19713 25194
rect 19617 25114 19713 25130
rect 19617 25050 19633 25114
rect 19697 25050 19713 25114
rect 19617 25034 19713 25050
rect 19617 24970 19633 25034
rect 19697 24970 19713 25034
rect 19876 25314 20202 25323
rect 19876 25010 19885 25314
rect 20189 25010 20202 25314
rect 19876 25001 20202 25010
rect 19617 24954 19713 24970
rect 19617 24890 19633 24954
rect 19697 24890 19713 24954
rect 19617 24874 19713 24890
rect 19882 24762 20202 25001
rect 20336 25434 20432 25450
rect 20336 25370 20352 25434
rect 20416 25370 20432 25434
rect 20336 25354 20432 25370
rect 20336 25290 20352 25354
rect 20416 25290 20432 25354
rect 20602 25323 20922 25701
rect 21055 25990 21071 26054
rect 21135 25990 21151 26054
rect 21774 26134 21870 26150
rect 21774 26070 21790 26134
rect 21854 26070 21870 26134
rect 21774 26054 21870 26070
rect 21322 26023 21642 26042
rect 21055 25974 21151 25990
rect 21055 25910 21071 25974
rect 21135 25910 21151 25974
rect 21055 25894 21151 25910
rect 21055 25830 21071 25894
rect 21135 25830 21151 25894
rect 21055 25814 21151 25830
rect 21055 25750 21071 25814
rect 21135 25750 21151 25814
rect 21055 25734 21151 25750
rect 21055 25670 21071 25734
rect 21135 25670 21151 25734
rect 21314 26014 21642 26023
rect 21314 25710 21323 26014
rect 21627 25710 21642 26014
rect 21314 25701 21642 25710
rect 21055 25654 21151 25670
rect 21055 25590 21071 25654
rect 21135 25590 21151 25654
rect 21055 25574 21151 25590
rect 20336 25274 20432 25290
rect 20336 25210 20352 25274
rect 20416 25210 20432 25274
rect 20336 25194 20432 25210
rect 20336 25130 20352 25194
rect 20416 25130 20432 25194
rect 20336 25114 20432 25130
rect 20336 25050 20352 25114
rect 20416 25050 20432 25114
rect 20336 25034 20432 25050
rect 20336 24970 20352 25034
rect 20416 24970 20432 25034
rect 20595 25314 20922 25323
rect 20595 25010 20604 25314
rect 20908 25010 20922 25314
rect 20595 25001 20922 25010
rect 20336 24954 20432 24970
rect 20336 24890 20352 24954
rect 20416 24890 20432 24954
rect 20336 24874 20432 24890
rect 20602 24762 20922 25001
rect 21055 25434 21151 25450
rect 21055 25370 21071 25434
rect 21135 25370 21151 25434
rect 21055 25354 21151 25370
rect 21055 25290 21071 25354
rect 21135 25290 21151 25354
rect 21322 25323 21642 25701
rect 21774 25990 21790 26054
rect 21854 25990 21870 26054
rect 22493 26134 22589 26150
rect 22493 26070 22509 26134
rect 22573 26070 22589 26134
rect 22493 26054 22589 26070
rect 22042 26023 22362 26042
rect 21774 25974 21870 25990
rect 21774 25910 21790 25974
rect 21854 25910 21870 25974
rect 21774 25894 21870 25910
rect 21774 25830 21790 25894
rect 21854 25830 21870 25894
rect 21774 25814 21870 25830
rect 21774 25750 21790 25814
rect 21854 25750 21870 25814
rect 21774 25734 21870 25750
rect 21774 25670 21790 25734
rect 21854 25670 21870 25734
rect 22033 26014 22362 26023
rect 22033 25710 22042 26014
rect 22346 25710 22362 26014
rect 22033 25701 22362 25710
rect 21774 25654 21870 25670
rect 21774 25590 21790 25654
rect 21854 25590 21870 25654
rect 21774 25574 21870 25590
rect 21055 25274 21151 25290
rect 21055 25210 21071 25274
rect 21135 25210 21151 25274
rect 21055 25194 21151 25210
rect 21055 25130 21071 25194
rect 21135 25130 21151 25194
rect 21055 25114 21151 25130
rect 21055 25050 21071 25114
rect 21135 25050 21151 25114
rect 21055 25034 21151 25050
rect 21055 24970 21071 25034
rect 21135 24970 21151 25034
rect 21314 25314 21642 25323
rect 21314 25010 21323 25314
rect 21627 25010 21642 25314
rect 21314 25001 21642 25010
rect 21055 24954 21151 24970
rect 21055 24890 21071 24954
rect 21135 24890 21151 24954
rect 21055 24874 21151 24890
rect 21322 24762 21642 25001
rect 21774 25434 21870 25450
rect 21774 25370 21790 25434
rect 21854 25370 21870 25434
rect 21774 25354 21870 25370
rect 21774 25290 21790 25354
rect 21854 25290 21870 25354
rect 22042 25323 22362 25701
rect 22493 25990 22509 26054
rect 22573 25990 22589 26054
rect 22493 25974 22589 25990
rect 22493 25910 22509 25974
rect 22573 25910 22589 25974
rect 22493 25894 22589 25910
rect 22493 25830 22509 25894
rect 22573 25830 22589 25894
rect 22493 25814 22589 25830
rect 22493 25750 22509 25814
rect 22573 25750 22589 25814
rect 22493 25734 22589 25750
rect 22493 25670 22509 25734
rect 22573 25670 22589 25734
rect 22493 25654 22589 25670
rect 22493 25590 22509 25654
rect 22573 25590 22589 25654
rect 22493 25574 22589 25590
rect 21774 25274 21870 25290
rect 21774 25210 21790 25274
rect 21854 25210 21870 25274
rect 21774 25194 21870 25210
rect 21774 25130 21790 25194
rect 21854 25130 21870 25194
rect 21774 25114 21870 25130
rect 21774 25050 21790 25114
rect 21854 25050 21870 25114
rect 21774 25034 21870 25050
rect 21774 24970 21790 25034
rect 21854 24970 21870 25034
rect 22033 25314 22362 25323
rect 22033 25010 22042 25314
rect 22346 25010 22362 25314
rect 22033 25001 22362 25010
rect 21774 24954 21870 24970
rect 21774 24890 21790 24954
rect 21854 24890 21870 24954
rect 21774 24874 21870 24890
rect 22042 24762 22362 25001
rect 22493 25434 22589 25450
rect 22493 25370 22509 25434
rect 22573 25370 22589 25434
rect 22493 25354 22589 25370
rect 22493 25290 22509 25354
rect 22573 25290 22589 25354
rect 22493 25274 22589 25290
rect 22493 25210 22509 25274
rect 22573 25210 22589 25274
rect 22493 25194 22589 25210
rect 22493 25130 22509 25194
rect 22573 25130 22589 25194
rect 22493 25114 22589 25130
rect 22493 25050 22509 25114
rect 22573 25052 22589 25114
rect 22783 25054 22849 25055
rect 22783 25052 22784 25054
rect 22573 25050 22784 25052
rect 22493 25034 22784 25050
rect 22493 24970 22509 25034
rect 22573 24992 22784 25034
rect 22573 24970 22589 24992
rect 22783 24990 22784 24992
rect 22848 24990 22849 25054
rect 22783 24989 22849 24990
rect 22493 24954 22589 24970
rect 22493 24890 22509 24954
rect 22573 24890 22589 24954
rect 22493 24874 22589 24890
rect 15424 24734 22592 24762
rect 15424 24670 15452 24734
rect 15516 24670 15532 24734
rect 15596 24670 22592 24734
rect 15424 24642 22592 24670
rect 15472 24567 15532 24642
rect 15469 24566 15535 24567
rect 15469 24502 15470 24566
rect 15534 24502 15535 24566
rect 15469 24501 15535 24502
rect 3348 22600 3372 22664
rect 3436 22600 3452 22664
rect 3516 22600 3532 22664
rect 3596 22600 3612 22664
rect 3676 22600 3692 22664
rect 3756 22600 3772 22664
rect 3836 22600 3852 22664
rect 3916 22600 3932 22664
rect 3996 22600 4012 22664
rect 4076 22600 4092 22664
rect 4156 22600 4172 22664
rect 4236 22600 4252 22664
rect 4316 22600 4332 22664
rect 4396 22600 4412 22664
rect 4476 22600 4492 22664
rect 4556 22600 4572 22664
rect 4636 22600 4652 22664
rect 4716 22600 4732 22664
rect 4796 22600 4812 22664
rect 4876 22600 4892 22664
rect 4956 22600 4980 22664
rect 43656 22664 45288 26360
rect 3348 18904 4980 22600
rect 14227 22614 14293 22615
rect 14227 22550 14228 22614
rect 14292 22550 14293 22614
rect 14227 22549 14293 22550
rect 43656 22600 43680 22664
rect 43744 22600 43760 22664
rect 43824 22600 43840 22664
rect 43904 22600 43920 22664
rect 43984 22600 44000 22664
rect 44064 22600 44080 22664
rect 44144 22600 44160 22664
rect 44224 22600 44240 22664
rect 44304 22600 44320 22664
rect 44384 22600 44400 22664
rect 44464 22600 44480 22664
rect 44544 22600 44560 22664
rect 44624 22600 44640 22664
rect 44704 22600 44720 22664
rect 44784 22600 44800 22664
rect 44864 22600 44880 22664
rect 44944 22600 44960 22664
rect 45024 22600 45040 22664
rect 45104 22600 45120 22664
rect 45184 22600 45200 22664
rect 45264 22600 45288 22664
rect 14230 22390 14290 22549
rect 14160 22374 14290 22390
rect 14160 22310 14176 22374
rect 14240 22310 14290 22374
rect 14160 22308 14290 22310
rect 14879 22374 14975 22390
rect 14879 22310 14895 22374
rect 14959 22310 14975 22374
rect 14160 22294 14256 22308
rect 13700 22263 14020 22282
rect 13700 22254 14022 22263
rect 13700 21950 13709 22254
rect 14013 21950 14022 22254
rect 13700 21941 14022 21950
rect 14160 22230 14176 22294
rect 14240 22230 14256 22294
rect 14879 22294 14975 22310
rect 14420 22263 14740 22282
rect 14160 22214 14256 22230
rect 14160 22150 14176 22214
rect 14240 22150 14256 22214
rect 14160 22134 14256 22150
rect 14160 22070 14176 22134
rect 14240 22070 14256 22134
rect 14160 22054 14256 22070
rect 14160 21990 14176 22054
rect 14240 21990 14256 22054
rect 14160 21974 14256 21990
rect 13700 21563 14020 21941
rect 14160 21910 14176 21974
rect 14240 21910 14256 21974
rect 14419 22254 14741 22263
rect 14419 21950 14428 22254
rect 14732 21950 14741 22254
rect 14419 21941 14741 21950
rect 14879 22230 14895 22294
rect 14959 22230 14975 22294
rect 15598 22374 15694 22390
rect 15598 22310 15614 22374
rect 15678 22310 15694 22374
rect 15598 22294 15694 22310
rect 15140 22263 15460 22282
rect 14879 22214 14975 22230
rect 14879 22150 14895 22214
rect 14959 22150 14975 22214
rect 14879 22134 14975 22150
rect 14879 22070 14895 22134
rect 14959 22070 14975 22134
rect 14879 22054 14975 22070
rect 14879 21990 14895 22054
rect 14959 21990 14975 22054
rect 14879 21974 14975 21990
rect 14160 21894 14256 21910
rect 14160 21830 14176 21894
rect 14240 21830 14256 21894
rect 14160 21814 14256 21830
rect 14160 21674 14256 21690
rect 14160 21610 14176 21674
rect 14240 21610 14256 21674
rect 14160 21594 14256 21610
rect 13700 21554 14022 21563
rect 13700 21250 13709 21554
rect 14013 21250 14022 21554
rect 13700 21241 14022 21250
rect 14160 21530 14176 21594
rect 14240 21530 14256 21594
rect 14420 21563 14740 21941
rect 14879 21910 14895 21974
rect 14959 21910 14975 21974
rect 15138 22254 15460 22263
rect 15138 21950 15147 22254
rect 15451 21950 15460 22254
rect 15138 21941 15460 21950
rect 14879 21894 14975 21910
rect 14879 21830 14895 21894
rect 14959 21830 14975 21894
rect 14879 21814 14975 21830
rect 14879 21674 14975 21690
rect 14879 21610 14895 21674
rect 14959 21610 14975 21674
rect 14879 21594 14975 21610
rect 14160 21514 14256 21530
rect 14160 21450 14176 21514
rect 14240 21450 14256 21514
rect 14160 21434 14256 21450
rect 14160 21370 14176 21434
rect 14240 21370 14256 21434
rect 14160 21354 14256 21370
rect 14160 21290 14176 21354
rect 14240 21290 14256 21354
rect 14160 21274 14256 21290
rect 13700 21002 14020 21241
rect 14160 21210 14176 21274
rect 14240 21210 14256 21274
rect 14419 21554 14741 21563
rect 14419 21250 14428 21554
rect 14732 21250 14741 21554
rect 14419 21241 14741 21250
rect 14879 21530 14895 21594
rect 14959 21530 14975 21594
rect 15140 21563 15460 21941
rect 15598 22230 15614 22294
rect 15678 22230 15694 22294
rect 16317 22374 16413 22390
rect 16317 22310 16333 22374
rect 16397 22310 16413 22374
rect 16317 22294 16413 22310
rect 15860 22263 16180 22282
rect 15598 22214 15694 22230
rect 15598 22150 15614 22214
rect 15678 22150 15694 22214
rect 15598 22134 15694 22150
rect 15598 22070 15614 22134
rect 15678 22070 15694 22134
rect 15598 22054 15694 22070
rect 15598 21990 15614 22054
rect 15678 21990 15694 22054
rect 15598 21974 15694 21990
rect 15598 21910 15614 21974
rect 15678 21910 15694 21974
rect 15857 22254 16180 22263
rect 15857 21950 15866 22254
rect 16170 21950 16180 22254
rect 15857 21941 16180 21950
rect 15598 21894 15694 21910
rect 15598 21830 15614 21894
rect 15678 21830 15694 21894
rect 15598 21814 15694 21830
rect 14879 21514 14975 21530
rect 14879 21450 14895 21514
rect 14959 21450 14975 21514
rect 14879 21434 14975 21450
rect 14879 21370 14895 21434
rect 14959 21370 14975 21434
rect 14879 21354 14975 21370
rect 14879 21290 14895 21354
rect 14959 21290 14975 21354
rect 14879 21274 14975 21290
rect 14160 21194 14256 21210
rect 14160 21130 14176 21194
rect 14240 21130 14256 21194
rect 14160 21114 14256 21130
rect 14420 21002 14740 21241
rect 14879 21210 14895 21274
rect 14959 21210 14975 21274
rect 15138 21554 15460 21563
rect 15138 21250 15147 21554
rect 15451 21250 15460 21554
rect 15138 21241 15460 21250
rect 14879 21194 14975 21210
rect 14879 21130 14895 21194
rect 14959 21130 14975 21194
rect 14879 21114 14975 21130
rect 15140 21002 15460 21241
rect 15598 21674 15694 21690
rect 15598 21610 15614 21674
rect 15678 21610 15694 21674
rect 15598 21594 15694 21610
rect 15598 21530 15614 21594
rect 15678 21530 15694 21594
rect 15860 21563 16180 21941
rect 16317 22230 16333 22294
rect 16397 22230 16413 22294
rect 17036 22374 17132 22390
rect 17036 22310 17052 22374
rect 17116 22310 17132 22374
rect 17036 22294 17132 22310
rect 16580 22263 16900 22282
rect 16317 22214 16413 22230
rect 16317 22150 16333 22214
rect 16397 22150 16413 22214
rect 16317 22134 16413 22150
rect 16317 22070 16333 22134
rect 16397 22070 16413 22134
rect 16317 22054 16413 22070
rect 16317 21990 16333 22054
rect 16397 21990 16413 22054
rect 16317 21974 16413 21990
rect 16317 21910 16333 21974
rect 16397 21910 16413 21974
rect 16576 22254 16900 22263
rect 16576 21950 16585 22254
rect 16889 21950 16900 22254
rect 16576 21941 16900 21950
rect 16317 21894 16413 21910
rect 16317 21830 16333 21894
rect 16397 21830 16413 21894
rect 16317 21814 16413 21830
rect 15598 21514 15694 21530
rect 15598 21450 15614 21514
rect 15678 21450 15694 21514
rect 15598 21434 15694 21450
rect 15598 21370 15614 21434
rect 15678 21370 15694 21434
rect 15598 21354 15694 21370
rect 15598 21290 15614 21354
rect 15678 21290 15694 21354
rect 15598 21274 15694 21290
rect 15598 21210 15614 21274
rect 15678 21210 15694 21274
rect 15857 21554 16180 21563
rect 15857 21250 15866 21554
rect 16170 21250 16180 21554
rect 15857 21241 16180 21250
rect 15598 21194 15694 21210
rect 15598 21130 15614 21194
rect 15678 21130 15694 21194
rect 15598 21114 15694 21130
rect 15860 21002 16180 21241
rect 16317 21674 16413 21690
rect 16317 21610 16333 21674
rect 16397 21610 16413 21674
rect 16317 21594 16413 21610
rect 16317 21530 16333 21594
rect 16397 21530 16413 21594
rect 16580 21563 16900 21941
rect 17036 22230 17052 22294
rect 17116 22230 17132 22294
rect 17755 22374 17851 22390
rect 17755 22310 17771 22374
rect 17835 22310 17851 22374
rect 17755 22294 17851 22310
rect 17300 22263 17620 22282
rect 17036 22214 17132 22230
rect 17036 22150 17052 22214
rect 17116 22150 17132 22214
rect 17036 22134 17132 22150
rect 17036 22070 17052 22134
rect 17116 22070 17132 22134
rect 17036 22054 17132 22070
rect 17036 21990 17052 22054
rect 17116 21990 17132 22054
rect 17036 21974 17132 21990
rect 17036 21910 17052 21974
rect 17116 21910 17132 21974
rect 17295 22254 17620 22263
rect 17295 21950 17304 22254
rect 17608 21950 17620 22254
rect 17295 21941 17620 21950
rect 17036 21894 17132 21910
rect 17036 21830 17052 21894
rect 17116 21830 17132 21894
rect 17036 21814 17132 21830
rect 16317 21514 16413 21530
rect 16317 21450 16333 21514
rect 16397 21450 16413 21514
rect 16317 21434 16413 21450
rect 16317 21370 16333 21434
rect 16397 21370 16413 21434
rect 16317 21354 16413 21370
rect 16317 21290 16333 21354
rect 16397 21290 16413 21354
rect 16317 21274 16413 21290
rect 16317 21210 16333 21274
rect 16397 21210 16413 21274
rect 16576 21554 16900 21563
rect 16576 21250 16585 21554
rect 16889 21250 16900 21554
rect 16576 21241 16900 21250
rect 16317 21194 16413 21210
rect 16317 21130 16333 21194
rect 16397 21130 16413 21194
rect 16317 21114 16413 21130
rect 16580 21002 16900 21241
rect 17036 21674 17132 21690
rect 17036 21610 17052 21674
rect 17116 21610 17132 21674
rect 17036 21594 17132 21610
rect 17036 21530 17052 21594
rect 17116 21530 17132 21594
rect 17300 21563 17620 21941
rect 17755 22230 17771 22294
rect 17835 22230 17851 22294
rect 18474 22374 18570 22390
rect 18474 22310 18490 22374
rect 18554 22310 18570 22374
rect 18474 22294 18570 22310
rect 18020 22263 18340 22282
rect 17755 22214 17851 22230
rect 17755 22150 17771 22214
rect 17835 22150 17851 22214
rect 17755 22134 17851 22150
rect 17755 22070 17771 22134
rect 17835 22070 17851 22134
rect 17755 22054 17851 22070
rect 17755 21990 17771 22054
rect 17835 21990 17851 22054
rect 17755 21974 17851 21990
rect 17755 21910 17771 21974
rect 17835 21910 17851 21974
rect 18014 22254 18340 22263
rect 18014 21950 18023 22254
rect 18327 21950 18340 22254
rect 18014 21941 18340 21950
rect 17755 21894 17851 21910
rect 17755 21830 17771 21894
rect 17835 21830 17851 21894
rect 17755 21814 17851 21830
rect 17036 21514 17132 21530
rect 17036 21450 17052 21514
rect 17116 21450 17132 21514
rect 17036 21434 17132 21450
rect 17036 21370 17052 21434
rect 17116 21370 17132 21434
rect 17036 21354 17132 21370
rect 17036 21290 17052 21354
rect 17116 21290 17132 21354
rect 17036 21274 17132 21290
rect 17036 21210 17052 21274
rect 17116 21210 17132 21274
rect 17295 21554 17620 21563
rect 17295 21250 17304 21554
rect 17608 21250 17620 21554
rect 17295 21241 17620 21250
rect 17036 21194 17132 21210
rect 17036 21130 17052 21194
rect 17116 21130 17132 21194
rect 17036 21114 17132 21130
rect 17300 21002 17620 21241
rect 17755 21674 17851 21690
rect 17755 21610 17771 21674
rect 17835 21610 17851 21674
rect 17755 21594 17851 21610
rect 17755 21530 17771 21594
rect 17835 21530 17851 21594
rect 18020 21563 18340 21941
rect 18474 22230 18490 22294
rect 18554 22230 18570 22294
rect 19193 22374 19289 22390
rect 19193 22310 19209 22374
rect 19273 22310 19289 22374
rect 19193 22294 19289 22310
rect 18740 22263 19060 22282
rect 18474 22214 18570 22230
rect 18474 22150 18490 22214
rect 18554 22150 18570 22214
rect 18474 22134 18570 22150
rect 18474 22070 18490 22134
rect 18554 22070 18570 22134
rect 18474 22054 18570 22070
rect 18474 21990 18490 22054
rect 18554 21990 18570 22054
rect 18474 21974 18570 21990
rect 18474 21910 18490 21974
rect 18554 21910 18570 21974
rect 18733 22254 19060 22263
rect 18733 21950 18742 22254
rect 19046 21950 19060 22254
rect 18733 21941 19060 21950
rect 18474 21894 18570 21910
rect 18474 21830 18490 21894
rect 18554 21830 18570 21894
rect 18474 21814 18570 21830
rect 17755 21514 17851 21530
rect 17755 21450 17771 21514
rect 17835 21450 17851 21514
rect 17755 21434 17851 21450
rect 17755 21370 17771 21434
rect 17835 21370 17851 21434
rect 17755 21354 17851 21370
rect 17755 21290 17771 21354
rect 17835 21290 17851 21354
rect 17755 21274 17851 21290
rect 17755 21210 17771 21274
rect 17835 21210 17851 21274
rect 18014 21554 18340 21563
rect 18014 21250 18023 21554
rect 18327 21250 18340 21554
rect 18014 21241 18340 21250
rect 17755 21194 17851 21210
rect 17755 21130 17771 21194
rect 17835 21130 17851 21194
rect 17755 21114 17851 21130
rect 18020 21002 18340 21241
rect 18474 21674 18570 21690
rect 18474 21610 18490 21674
rect 18554 21610 18570 21674
rect 18474 21594 18570 21610
rect 18474 21530 18490 21594
rect 18554 21530 18570 21594
rect 18740 21563 19060 21941
rect 19193 22230 19209 22294
rect 19273 22230 19289 22294
rect 19912 22374 20008 22390
rect 19912 22310 19928 22374
rect 19992 22310 20008 22374
rect 19912 22294 20008 22310
rect 19460 22263 19780 22282
rect 19193 22214 19289 22230
rect 19193 22150 19209 22214
rect 19273 22150 19289 22214
rect 19193 22134 19289 22150
rect 19193 22070 19209 22134
rect 19273 22070 19289 22134
rect 19193 22054 19289 22070
rect 19193 21990 19209 22054
rect 19273 21990 19289 22054
rect 19193 21974 19289 21990
rect 19193 21910 19209 21974
rect 19273 21910 19289 21974
rect 19452 22254 19780 22263
rect 19452 21950 19461 22254
rect 19765 21950 19780 22254
rect 19452 21941 19780 21950
rect 19193 21894 19289 21910
rect 19193 21830 19209 21894
rect 19273 21830 19289 21894
rect 19193 21814 19289 21830
rect 18474 21514 18570 21530
rect 18474 21450 18490 21514
rect 18554 21450 18570 21514
rect 18474 21434 18570 21450
rect 18474 21370 18490 21434
rect 18554 21370 18570 21434
rect 18474 21354 18570 21370
rect 18474 21290 18490 21354
rect 18554 21290 18570 21354
rect 18474 21274 18570 21290
rect 18474 21210 18490 21274
rect 18554 21210 18570 21274
rect 18733 21554 19060 21563
rect 18733 21250 18742 21554
rect 19046 21250 19060 21554
rect 18733 21241 19060 21250
rect 18474 21194 18570 21210
rect 18474 21130 18490 21194
rect 18554 21130 18570 21194
rect 18474 21114 18570 21130
rect 18740 21002 19060 21241
rect 19193 21674 19289 21690
rect 19193 21610 19209 21674
rect 19273 21610 19289 21674
rect 19193 21594 19289 21610
rect 19193 21530 19209 21594
rect 19273 21530 19289 21594
rect 19460 21563 19780 21941
rect 19912 22230 19928 22294
rect 19992 22230 20008 22294
rect 20631 22374 20727 22390
rect 20631 22310 20647 22374
rect 20711 22310 20727 22374
rect 20631 22294 20727 22310
rect 20180 22263 20500 22282
rect 19912 22214 20008 22230
rect 19912 22150 19928 22214
rect 19992 22150 20008 22214
rect 19912 22134 20008 22150
rect 19912 22070 19928 22134
rect 19992 22070 20008 22134
rect 19912 22054 20008 22070
rect 19912 21990 19928 22054
rect 19992 21990 20008 22054
rect 19912 21974 20008 21990
rect 19912 21910 19928 21974
rect 19992 21910 20008 21974
rect 20171 22254 20500 22263
rect 20171 21950 20180 22254
rect 20484 21950 20500 22254
rect 20171 21941 20500 21950
rect 19912 21894 20008 21910
rect 19912 21830 19928 21894
rect 19992 21830 20008 21894
rect 19912 21814 20008 21830
rect 19193 21514 19289 21530
rect 19193 21450 19209 21514
rect 19273 21450 19289 21514
rect 19193 21434 19289 21450
rect 19193 21370 19209 21434
rect 19273 21370 19289 21434
rect 19193 21354 19289 21370
rect 19193 21290 19209 21354
rect 19273 21290 19289 21354
rect 19193 21274 19289 21290
rect 19193 21210 19209 21274
rect 19273 21210 19289 21274
rect 19452 21554 19780 21563
rect 19452 21250 19461 21554
rect 19765 21250 19780 21554
rect 19452 21241 19780 21250
rect 19193 21194 19289 21210
rect 19193 21130 19209 21194
rect 19273 21130 19289 21194
rect 19193 21114 19289 21130
rect 19460 21002 19780 21241
rect 19912 21674 20008 21690
rect 19912 21610 19928 21674
rect 19992 21610 20008 21674
rect 19912 21594 20008 21610
rect 19912 21530 19928 21594
rect 19992 21530 20008 21594
rect 20180 21563 20500 21941
rect 20631 22230 20647 22294
rect 20711 22230 20727 22294
rect 20631 22214 20727 22230
rect 20631 22150 20647 22214
rect 20711 22150 20727 22214
rect 20631 22134 20727 22150
rect 20631 22070 20647 22134
rect 20711 22070 20727 22134
rect 20631 22054 20727 22070
rect 20631 21990 20647 22054
rect 20711 21990 20727 22054
rect 20631 21974 20727 21990
rect 20631 21910 20647 21974
rect 20711 21910 20727 21974
rect 20631 21894 20727 21910
rect 20631 21830 20647 21894
rect 20711 21830 20727 21894
rect 20631 21814 20727 21830
rect 19912 21514 20008 21530
rect 19912 21450 19928 21514
rect 19992 21450 20008 21514
rect 19912 21434 20008 21450
rect 19912 21370 19928 21434
rect 19992 21370 20008 21434
rect 19912 21354 20008 21370
rect 19912 21290 19928 21354
rect 19992 21290 20008 21354
rect 19912 21274 20008 21290
rect 19912 21210 19928 21274
rect 19992 21210 20008 21274
rect 20171 21554 20500 21563
rect 20171 21250 20180 21554
rect 20484 21250 20500 21554
rect 20171 21241 20500 21250
rect 19912 21194 20008 21210
rect 19912 21130 19928 21194
rect 19992 21130 20008 21194
rect 19912 21114 20008 21130
rect 20180 21002 20500 21241
rect 20631 21674 20727 21690
rect 20631 21610 20647 21674
rect 20711 21636 20727 21674
rect 20851 21638 20917 21639
rect 20851 21636 20852 21638
rect 20711 21610 20852 21636
rect 20631 21594 20852 21610
rect 20631 21530 20647 21594
rect 20711 21576 20852 21594
rect 20711 21530 20727 21576
rect 20851 21574 20852 21576
rect 20916 21574 20917 21638
rect 20851 21573 20917 21574
rect 20631 21514 20727 21530
rect 20631 21450 20647 21514
rect 20711 21450 20727 21514
rect 20631 21434 20727 21450
rect 20631 21370 20647 21434
rect 20711 21370 20727 21434
rect 20631 21354 20727 21370
rect 20631 21290 20647 21354
rect 20711 21290 20727 21354
rect 20631 21274 20727 21290
rect 20631 21210 20647 21274
rect 20711 21210 20727 21274
rect 20631 21194 20727 21210
rect 20631 21130 20647 21194
rect 20711 21130 20727 21194
rect 20631 21114 20727 21130
rect 13562 20974 20730 21002
rect 13562 20910 13590 20974
rect 13654 20910 13670 20974
rect 13734 20910 20730 20974
rect 13562 20906 20730 20910
rect 13562 20882 14090 20906
rect 14089 20842 14090 20882
rect 14154 20882 20730 20906
rect 14154 20842 14155 20882
rect 14089 20841 14155 20842
rect 20854 19684 20914 21573
rect 20854 19624 21052 19684
rect 20992 18955 21052 19624
rect 3348 18840 3372 18904
rect 3436 18840 3452 18904
rect 3516 18840 3532 18904
rect 3596 18840 3612 18904
rect 3676 18840 3692 18904
rect 3756 18840 3772 18904
rect 3836 18840 3852 18904
rect 3916 18840 3932 18904
rect 3996 18840 4012 18904
rect 4076 18840 4092 18904
rect 4156 18840 4172 18904
rect 4236 18840 4252 18904
rect 4316 18840 4332 18904
rect 4396 18840 4412 18904
rect 4476 18840 4492 18904
rect 4556 18840 4572 18904
rect 4636 18840 4652 18904
rect 4716 18840 4732 18904
rect 4796 18840 4812 18904
rect 4876 18840 4892 18904
rect 4956 18840 4980 18904
rect 20989 18954 21055 18955
rect 20989 18890 20990 18954
rect 21054 18952 21055 18954
rect 21054 18890 21086 18952
rect 20989 18889 21086 18890
rect 3348 15144 4980 18840
rect 21026 18630 21086 18889
rect 43656 18904 45288 22600
rect 43656 18840 43680 18904
rect 43744 18840 43760 18904
rect 43824 18840 43840 18904
rect 43904 18840 43920 18904
rect 43984 18840 44000 18904
rect 44064 18840 44080 18904
rect 44144 18840 44160 18904
rect 44224 18840 44240 18904
rect 44304 18840 44320 18904
rect 44384 18840 44400 18904
rect 44464 18840 44480 18904
rect 44544 18840 44560 18904
rect 44624 18840 44640 18904
rect 44704 18840 44720 18904
rect 44784 18840 44800 18904
rect 44864 18840 44880 18904
rect 44944 18840 44960 18904
rect 45024 18840 45040 18904
rect 45104 18840 45120 18904
rect 45184 18840 45200 18904
rect 45264 18840 45288 18904
rect 16708 18614 16804 18630
rect 16708 18550 16724 18614
rect 16788 18550 16804 18614
rect 16708 18534 16804 18550
rect 16248 18503 16568 18522
rect 16248 18494 16570 18503
rect 16248 18190 16257 18494
rect 16561 18190 16570 18494
rect 16248 18181 16570 18190
rect 16708 18470 16724 18534
rect 16788 18470 16804 18534
rect 17427 18614 17523 18630
rect 17427 18550 17443 18614
rect 17507 18550 17523 18614
rect 17427 18534 17523 18550
rect 16968 18503 17288 18522
rect 16708 18454 16804 18470
rect 16708 18390 16724 18454
rect 16788 18390 16804 18454
rect 16708 18374 16804 18390
rect 16708 18310 16724 18374
rect 16788 18310 16804 18374
rect 16708 18294 16804 18310
rect 16708 18230 16724 18294
rect 16788 18230 16804 18294
rect 16708 18214 16804 18230
rect 16248 17803 16568 18181
rect 16708 18150 16724 18214
rect 16788 18150 16804 18214
rect 16967 18494 17289 18503
rect 16967 18190 16976 18494
rect 17280 18190 17289 18494
rect 16967 18181 17289 18190
rect 17427 18470 17443 18534
rect 17507 18470 17523 18534
rect 18146 18614 18242 18630
rect 18146 18550 18162 18614
rect 18226 18550 18242 18614
rect 18146 18534 18242 18550
rect 17688 18503 18008 18522
rect 17427 18454 17523 18470
rect 17427 18390 17443 18454
rect 17507 18390 17523 18454
rect 17427 18374 17523 18390
rect 17427 18310 17443 18374
rect 17507 18310 17523 18374
rect 17427 18294 17523 18310
rect 17427 18230 17443 18294
rect 17507 18230 17523 18294
rect 17427 18214 17523 18230
rect 16708 18134 16804 18150
rect 16708 18070 16724 18134
rect 16788 18070 16804 18134
rect 16708 18054 16804 18070
rect 16708 17914 16804 17930
rect 16708 17850 16724 17914
rect 16788 17850 16804 17914
rect 16708 17834 16804 17850
rect 16248 17794 16570 17803
rect 16248 17490 16257 17794
rect 16561 17490 16570 17794
rect 16248 17481 16570 17490
rect 16708 17770 16724 17834
rect 16788 17770 16804 17834
rect 16968 17803 17288 18181
rect 17427 18150 17443 18214
rect 17507 18150 17523 18214
rect 17686 18494 18008 18503
rect 17686 18190 17695 18494
rect 17999 18190 18008 18494
rect 17686 18181 18008 18190
rect 17427 18134 17523 18150
rect 17427 18070 17443 18134
rect 17507 18070 17523 18134
rect 17427 18054 17523 18070
rect 17427 17914 17523 17930
rect 17427 17850 17443 17914
rect 17507 17850 17523 17914
rect 17427 17834 17523 17850
rect 16708 17754 16804 17770
rect 16708 17690 16724 17754
rect 16788 17690 16804 17754
rect 16708 17674 16804 17690
rect 16708 17610 16724 17674
rect 16788 17610 16804 17674
rect 16708 17594 16804 17610
rect 16708 17530 16724 17594
rect 16788 17530 16804 17594
rect 16708 17514 16804 17530
rect 16248 17242 16568 17481
rect 16708 17450 16724 17514
rect 16788 17450 16804 17514
rect 16967 17794 17289 17803
rect 16967 17490 16976 17794
rect 17280 17490 17289 17794
rect 16967 17481 17289 17490
rect 17427 17770 17443 17834
rect 17507 17770 17523 17834
rect 17688 17803 18008 18181
rect 18146 18470 18162 18534
rect 18226 18470 18242 18534
rect 18865 18614 18961 18630
rect 18865 18550 18881 18614
rect 18945 18550 18961 18614
rect 18865 18534 18961 18550
rect 18408 18503 18728 18522
rect 18146 18454 18242 18470
rect 18146 18390 18162 18454
rect 18226 18390 18242 18454
rect 18146 18374 18242 18390
rect 18146 18310 18162 18374
rect 18226 18310 18242 18374
rect 18146 18294 18242 18310
rect 18146 18230 18162 18294
rect 18226 18230 18242 18294
rect 18146 18214 18242 18230
rect 18146 18150 18162 18214
rect 18226 18150 18242 18214
rect 18405 18494 18728 18503
rect 18405 18190 18414 18494
rect 18718 18190 18728 18494
rect 18405 18181 18728 18190
rect 18146 18134 18242 18150
rect 18146 18070 18162 18134
rect 18226 18070 18242 18134
rect 18146 18054 18242 18070
rect 17427 17754 17523 17770
rect 17427 17690 17443 17754
rect 17507 17690 17523 17754
rect 17427 17674 17523 17690
rect 17427 17610 17443 17674
rect 17507 17610 17523 17674
rect 17427 17594 17523 17610
rect 17427 17530 17443 17594
rect 17507 17530 17523 17594
rect 17427 17514 17523 17530
rect 16708 17434 16804 17450
rect 16708 17370 16724 17434
rect 16788 17370 16804 17434
rect 16708 17354 16804 17370
rect 16968 17242 17288 17481
rect 17427 17450 17443 17514
rect 17507 17450 17523 17514
rect 17686 17794 18008 17803
rect 17686 17490 17695 17794
rect 17999 17490 18008 17794
rect 17686 17481 18008 17490
rect 17427 17434 17523 17450
rect 17427 17370 17443 17434
rect 17507 17370 17523 17434
rect 17427 17354 17523 17370
rect 17688 17242 18008 17481
rect 18146 17914 18242 17930
rect 18146 17850 18162 17914
rect 18226 17850 18242 17914
rect 18146 17834 18242 17850
rect 18146 17770 18162 17834
rect 18226 17770 18242 17834
rect 18408 17803 18728 18181
rect 18865 18470 18881 18534
rect 18945 18470 18961 18534
rect 19584 18614 19680 18630
rect 19584 18550 19600 18614
rect 19664 18550 19680 18614
rect 19584 18534 19680 18550
rect 19128 18503 19448 18522
rect 18865 18454 18961 18470
rect 18865 18390 18881 18454
rect 18945 18390 18961 18454
rect 18865 18374 18961 18390
rect 18865 18310 18881 18374
rect 18945 18310 18961 18374
rect 18865 18294 18961 18310
rect 18865 18230 18881 18294
rect 18945 18230 18961 18294
rect 18865 18214 18961 18230
rect 18865 18150 18881 18214
rect 18945 18150 18961 18214
rect 19124 18494 19448 18503
rect 19124 18190 19133 18494
rect 19437 18190 19448 18494
rect 19124 18181 19448 18190
rect 18865 18134 18961 18150
rect 18865 18070 18881 18134
rect 18945 18070 18961 18134
rect 18865 18054 18961 18070
rect 18146 17754 18242 17770
rect 18146 17690 18162 17754
rect 18226 17690 18242 17754
rect 18146 17674 18242 17690
rect 18146 17610 18162 17674
rect 18226 17610 18242 17674
rect 18146 17594 18242 17610
rect 18146 17530 18162 17594
rect 18226 17530 18242 17594
rect 18146 17514 18242 17530
rect 18146 17450 18162 17514
rect 18226 17450 18242 17514
rect 18405 17794 18728 17803
rect 18405 17490 18414 17794
rect 18718 17490 18728 17794
rect 18405 17481 18728 17490
rect 18146 17434 18242 17450
rect 18146 17370 18162 17434
rect 18226 17370 18242 17434
rect 18146 17354 18242 17370
rect 18408 17242 18728 17481
rect 18865 17914 18961 17930
rect 18865 17850 18881 17914
rect 18945 17850 18961 17914
rect 18865 17834 18961 17850
rect 18865 17770 18881 17834
rect 18945 17770 18961 17834
rect 19128 17803 19448 18181
rect 19584 18470 19600 18534
rect 19664 18470 19680 18534
rect 20303 18614 20399 18630
rect 20303 18550 20319 18614
rect 20383 18550 20399 18614
rect 20303 18534 20399 18550
rect 19848 18503 20168 18522
rect 19584 18454 19680 18470
rect 19584 18390 19600 18454
rect 19664 18390 19680 18454
rect 19584 18374 19680 18390
rect 19584 18310 19600 18374
rect 19664 18310 19680 18374
rect 19584 18294 19680 18310
rect 19584 18230 19600 18294
rect 19664 18230 19680 18294
rect 19584 18214 19680 18230
rect 19584 18150 19600 18214
rect 19664 18150 19680 18214
rect 19843 18494 20168 18503
rect 19843 18190 19852 18494
rect 20156 18190 20168 18494
rect 19843 18181 20168 18190
rect 19584 18134 19680 18150
rect 19584 18070 19600 18134
rect 19664 18070 19680 18134
rect 19584 18054 19680 18070
rect 18865 17754 18961 17770
rect 18865 17690 18881 17754
rect 18945 17690 18961 17754
rect 18865 17674 18961 17690
rect 18865 17610 18881 17674
rect 18945 17610 18961 17674
rect 18865 17594 18961 17610
rect 18865 17530 18881 17594
rect 18945 17530 18961 17594
rect 18865 17514 18961 17530
rect 18865 17450 18881 17514
rect 18945 17450 18961 17514
rect 19124 17794 19448 17803
rect 19124 17490 19133 17794
rect 19437 17490 19448 17794
rect 19124 17481 19448 17490
rect 18865 17434 18961 17450
rect 18865 17370 18881 17434
rect 18945 17370 18961 17434
rect 18865 17354 18961 17370
rect 19128 17242 19448 17481
rect 19584 17914 19680 17930
rect 19584 17850 19600 17914
rect 19664 17850 19680 17914
rect 19584 17834 19680 17850
rect 19584 17770 19600 17834
rect 19664 17770 19680 17834
rect 19848 17803 20168 18181
rect 20303 18470 20319 18534
rect 20383 18470 20399 18534
rect 21022 18614 21118 18630
rect 21022 18550 21038 18614
rect 21102 18550 21118 18614
rect 21022 18534 21118 18550
rect 20568 18503 20888 18522
rect 20303 18454 20399 18470
rect 20303 18390 20319 18454
rect 20383 18390 20399 18454
rect 20303 18374 20399 18390
rect 20303 18310 20319 18374
rect 20383 18310 20399 18374
rect 20303 18294 20399 18310
rect 20303 18230 20319 18294
rect 20383 18230 20399 18294
rect 20303 18214 20399 18230
rect 20303 18150 20319 18214
rect 20383 18150 20399 18214
rect 20562 18494 20888 18503
rect 20562 18190 20571 18494
rect 20875 18190 20888 18494
rect 20562 18181 20888 18190
rect 20303 18134 20399 18150
rect 20303 18070 20319 18134
rect 20383 18070 20399 18134
rect 20303 18054 20399 18070
rect 19584 17754 19680 17770
rect 19584 17690 19600 17754
rect 19664 17690 19680 17754
rect 19584 17674 19680 17690
rect 19584 17610 19600 17674
rect 19664 17610 19680 17674
rect 19584 17594 19680 17610
rect 19584 17530 19600 17594
rect 19664 17530 19680 17594
rect 19584 17514 19680 17530
rect 19584 17450 19600 17514
rect 19664 17450 19680 17514
rect 19843 17794 20168 17803
rect 19843 17490 19852 17794
rect 20156 17490 20168 17794
rect 19843 17481 20168 17490
rect 19584 17434 19680 17450
rect 19584 17370 19600 17434
rect 19664 17370 19680 17434
rect 19584 17354 19680 17370
rect 19848 17242 20168 17481
rect 20303 17914 20399 17930
rect 20303 17850 20319 17914
rect 20383 17850 20399 17914
rect 20303 17834 20399 17850
rect 20303 17770 20319 17834
rect 20383 17770 20399 17834
rect 20568 17803 20888 18181
rect 21022 18470 21038 18534
rect 21102 18470 21118 18534
rect 21741 18614 21837 18630
rect 21741 18550 21757 18614
rect 21821 18550 21837 18614
rect 21741 18534 21837 18550
rect 21288 18503 21608 18522
rect 21022 18454 21118 18470
rect 21022 18390 21038 18454
rect 21102 18390 21118 18454
rect 21022 18374 21118 18390
rect 21022 18310 21038 18374
rect 21102 18310 21118 18374
rect 21022 18294 21118 18310
rect 21022 18230 21038 18294
rect 21102 18230 21118 18294
rect 21022 18214 21118 18230
rect 21022 18150 21038 18214
rect 21102 18150 21118 18214
rect 21281 18494 21608 18503
rect 21281 18190 21290 18494
rect 21594 18190 21608 18494
rect 21281 18181 21608 18190
rect 21022 18134 21118 18150
rect 21022 18070 21038 18134
rect 21102 18070 21118 18134
rect 21022 18054 21118 18070
rect 20303 17754 20399 17770
rect 20303 17690 20319 17754
rect 20383 17690 20399 17754
rect 20303 17674 20399 17690
rect 20303 17610 20319 17674
rect 20383 17610 20399 17674
rect 20303 17594 20399 17610
rect 20303 17530 20319 17594
rect 20383 17530 20399 17594
rect 20303 17514 20399 17530
rect 20303 17450 20319 17514
rect 20383 17450 20399 17514
rect 20562 17794 20888 17803
rect 20562 17490 20571 17794
rect 20875 17490 20888 17794
rect 20562 17481 20888 17490
rect 20303 17434 20399 17450
rect 20303 17370 20319 17434
rect 20383 17370 20399 17434
rect 20303 17354 20399 17370
rect 20568 17242 20888 17481
rect 21022 17914 21118 17930
rect 21022 17850 21038 17914
rect 21102 17850 21118 17914
rect 21022 17834 21118 17850
rect 21022 17770 21038 17834
rect 21102 17770 21118 17834
rect 21288 17803 21608 18181
rect 21741 18470 21757 18534
rect 21821 18470 21837 18534
rect 22460 18614 22556 18630
rect 22460 18550 22476 18614
rect 22540 18550 22556 18614
rect 22460 18534 22556 18550
rect 22008 18503 22328 18522
rect 21741 18454 21837 18470
rect 21741 18390 21757 18454
rect 21821 18390 21837 18454
rect 21741 18374 21837 18390
rect 21741 18310 21757 18374
rect 21821 18310 21837 18374
rect 21741 18294 21837 18310
rect 21741 18230 21757 18294
rect 21821 18230 21837 18294
rect 21741 18214 21837 18230
rect 21741 18150 21757 18214
rect 21821 18150 21837 18214
rect 22000 18494 22328 18503
rect 22000 18190 22009 18494
rect 22313 18190 22328 18494
rect 22000 18181 22328 18190
rect 21741 18134 21837 18150
rect 21741 18070 21757 18134
rect 21821 18070 21837 18134
rect 21741 18054 21837 18070
rect 21022 17754 21118 17770
rect 21022 17690 21038 17754
rect 21102 17690 21118 17754
rect 21022 17674 21118 17690
rect 21022 17610 21038 17674
rect 21102 17610 21118 17674
rect 21022 17594 21118 17610
rect 21022 17530 21038 17594
rect 21102 17530 21118 17594
rect 21022 17514 21118 17530
rect 21022 17450 21038 17514
rect 21102 17450 21118 17514
rect 21281 17794 21608 17803
rect 21281 17490 21290 17794
rect 21594 17490 21608 17794
rect 21281 17481 21608 17490
rect 21022 17434 21118 17450
rect 21022 17370 21038 17434
rect 21102 17370 21118 17434
rect 21022 17354 21118 17370
rect 21288 17242 21608 17481
rect 21741 17914 21837 17930
rect 21741 17850 21757 17914
rect 21821 17850 21837 17914
rect 21741 17834 21837 17850
rect 21741 17770 21757 17834
rect 21821 17770 21837 17834
rect 22008 17803 22328 18181
rect 22460 18470 22476 18534
rect 22540 18470 22556 18534
rect 23179 18614 23275 18630
rect 23179 18550 23195 18614
rect 23259 18550 23275 18614
rect 23179 18534 23275 18550
rect 22728 18503 23048 18522
rect 22460 18454 22556 18470
rect 22460 18390 22476 18454
rect 22540 18390 22556 18454
rect 22460 18374 22556 18390
rect 22460 18310 22476 18374
rect 22540 18310 22556 18374
rect 22460 18294 22556 18310
rect 22460 18230 22476 18294
rect 22540 18230 22556 18294
rect 22460 18214 22556 18230
rect 22460 18150 22476 18214
rect 22540 18150 22556 18214
rect 22719 18494 23048 18503
rect 22719 18190 22728 18494
rect 23032 18190 23048 18494
rect 22719 18181 23048 18190
rect 22460 18134 22556 18150
rect 22460 18070 22476 18134
rect 22540 18070 22556 18134
rect 22460 18054 22556 18070
rect 21741 17754 21837 17770
rect 21741 17690 21757 17754
rect 21821 17690 21837 17754
rect 21741 17674 21837 17690
rect 21741 17610 21757 17674
rect 21821 17610 21837 17674
rect 21741 17594 21837 17610
rect 21741 17530 21757 17594
rect 21821 17530 21837 17594
rect 21741 17514 21837 17530
rect 21741 17450 21757 17514
rect 21821 17450 21837 17514
rect 22000 17794 22328 17803
rect 22000 17490 22009 17794
rect 22313 17490 22328 17794
rect 22000 17481 22328 17490
rect 21741 17434 21837 17450
rect 21741 17370 21757 17434
rect 21821 17370 21837 17434
rect 21741 17354 21837 17370
rect 22008 17242 22328 17481
rect 22460 17914 22556 17930
rect 22460 17850 22476 17914
rect 22540 17850 22556 17914
rect 22460 17834 22556 17850
rect 22460 17770 22476 17834
rect 22540 17770 22556 17834
rect 22728 17803 23048 18181
rect 23179 18470 23195 18534
rect 23259 18470 23275 18534
rect 23179 18454 23275 18470
rect 23179 18390 23195 18454
rect 23259 18390 23275 18454
rect 23179 18374 23275 18390
rect 23179 18310 23195 18374
rect 23259 18310 23275 18374
rect 23179 18294 23275 18310
rect 23179 18230 23195 18294
rect 23259 18230 23275 18294
rect 23179 18214 23275 18230
rect 23179 18150 23195 18214
rect 23259 18150 23275 18214
rect 23179 18134 23275 18150
rect 23179 18070 23195 18134
rect 23259 18070 23275 18134
rect 23179 18054 23275 18070
rect 22460 17754 22556 17770
rect 22460 17690 22476 17754
rect 22540 17690 22556 17754
rect 22460 17674 22556 17690
rect 22460 17610 22476 17674
rect 22540 17610 22556 17674
rect 22460 17594 22556 17610
rect 22460 17530 22476 17594
rect 22540 17530 22556 17594
rect 22460 17514 22556 17530
rect 22460 17450 22476 17514
rect 22540 17450 22556 17514
rect 22719 17794 23048 17803
rect 22719 17490 22728 17794
rect 23032 17490 23048 17794
rect 22719 17481 23048 17490
rect 22460 17434 22556 17450
rect 22460 17370 22476 17434
rect 22540 17370 22556 17434
rect 22460 17354 22556 17370
rect 22728 17242 23048 17481
rect 23179 17914 23275 17930
rect 23179 17850 23195 17914
rect 23259 17850 23275 17914
rect 23179 17834 23275 17850
rect 23179 17770 23195 17834
rect 23259 17770 23275 17834
rect 23179 17754 23275 17770
rect 23179 17690 23195 17754
rect 23259 17690 23275 17754
rect 23179 17674 23275 17690
rect 23179 17610 23195 17674
rect 23259 17610 23275 17674
rect 23179 17594 23275 17610
rect 23179 17530 23195 17594
rect 23259 17530 23275 17594
rect 23179 17514 23275 17530
rect 23179 17450 23195 17514
rect 23259 17450 23275 17514
rect 23179 17434 23275 17450
rect 23179 17370 23195 17434
rect 23259 17370 23275 17434
rect 23179 17354 23275 17370
rect 16110 17214 23278 17242
rect 16110 17150 16138 17214
rect 16202 17150 16218 17214
rect 16282 17150 23278 17214
rect 16110 17122 23278 17150
rect 17404 17003 17464 17122
rect 17401 17002 17467 17003
rect 17401 16938 17402 17002
rect 17466 16938 17467 17002
rect 17401 16937 17467 16938
rect 19609 16392 19675 16393
rect 19609 16328 19610 16392
rect 19674 16328 19675 16392
rect 19609 16327 19675 16328
rect 3348 15080 3372 15144
rect 3436 15080 3452 15144
rect 3516 15080 3532 15144
rect 3596 15080 3612 15144
rect 3676 15080 3692 15144
rect 3756 15080 3772 15144
rect 3836 15080 3852 15144
rect 3916 15080 3932 15144
rect 3996 15080 4012 15144
rect 4076 15080 4092 15144
rect 4156 15080 4172 15144
rect 4236 15080 4252 15144
rect 4316 15080 4332 15144
rect 4396 15080 4412 15144
rect 4476 15080 4492 15144
rect 4556 15080 4572 15144
rect 4636 15080 4652 15144
rect 4716 15080 4732 15144
rect 4796 15080 4812 15144
rect 4876 15080 4892 15144
rect 4956 15080 4980 15144
rect 3348 11384 4980 15080
rect 19612 14870 19672 16327
rect 43656 15144 45288 18840
rect 43656 15080 43680 15144
rect 43744 15080 43760 15144
rect 43824 15080 43840 15144
rect 43904 15080 43920 15144
rect 43984 15080 44000 15144
rect 44064 15080 44080 15144
rect 44144 15080 44160 15144
rect 44224 15080 44240 15144
rect 44304 15080 44320 15144
rect 44384 15080 44400 15144
rect 44464 15080 44480 15144
rect 44544 15080 44560 15144
rect 44624 15080 44640 15144
rect 44704 15080 44720 15144
rect 44784 15080 44800 15144
rect 44864 15080 44880 15144
rect 44944 15080 44960 15144
rect 45024 15080 45040 15144
rect 45104 15080 45120 15144
rect 45184 15080 45200 15144
rect 45264 15080 45288 15144
rect 16708 14854 16804 14870
rect 16708 14790 16724 14854
rect 16788 14790 16804 14854
rect 16708 14774 16804 14790
rect 16248 14743 16568 14762
rect 16248 14734 16570 14743
rect 16248 14430 16257 14734
rect 16561 14430 16570 14734
rect 16248 14421 16570 14430
rect 16708 14710 16724 14774
rect 16788 14710 16804 14774
rect 17427 14854 17523 14870
rect 17427 14790 17443 14854
rect 17507 14790 17523 14854
rect 17427 14774 17523 14790
rect 16968 14743 17288 14762
rect 16708 14694 16804 14710
rect 16708 14630 16724 14694
rect 16788 14630 16804 14694
rect 16708 14614 16804 14630
rect 16708 14550 16724 14614
rect 16788 14550 16804 14614
rect 16708 14534 16804 14550
rect 16708 14470 16724 14534
rect 16788 14470 16804 14534
rect 16708 14454 16804 14470
rect 16248 14043 16568 14421
rect 16708 14390 16724 14454
rect 16788 14390 16804 14454
rect 16967 14734 17289 14743
rect 16967 14430 16976 14734
rect 17280 14430 17289 14734
rect 16967 14421 17289 14430
rect 17427 14710 17443 14774
rect 17507 14710 17523 14774
rect 18146 14854 18242 14870
rect 18146 14790 18162 14854
rect 18226 14790 18242 14854
rect 18146 14774 18242 14790
rect 17688 14743 18008 14762
rect 17427 14694 17523 14710
rect 17427 14630 17443 14694
rect 17507 14630 17523 14694
rect 17427 14614 17523 14630
rect 17427 14550 17443 14614
rect 17507 14550 17523 14614
rect 17427 14534 17523 14550
rect 17427 14470 17443 14534
rect 17507 14470 17523 14534
rect 17427 14454 17523 14470
rect 16708 14374 16804 14390
rect 16708 14310 16724 14374
rect 16788 14310 16804 14374
rect 16708 14294 16804 14310
rect 16708 14154 16804 14170
rect 16708 14090 16724 14154
rect 16788 14090 16804 14154
rect 16708 14074 16804 14090
rect 16248 14034 16570 14043
rect 16248 13730 16257 14034
rect 16561 13730 16570 14034
rect 16248 13721 16570 13730
rect 16708 14010 16724 14074
rect 16788 14010 16804 14074
rect 16968 14043 17288 14421
rect 17427 14390 17443 14454
rect 17507 14390 17523 14454
rect 17686 14734 18008 14743
rect 17686 14430 17695 14734
rect 17999 14430 18008 14734
rect 17686 14421 18008 14430
rect 17427 14374 17523 14390
rect 17427 14310 17443 14374
rect 17507 14310 17523 14374
rect 17427 14294 17523 14310
rect 17427 14154 17523 14170
rect 17427 14090 17443 14154
rect 17507 14090 17523 14154
rect 17427 14074 17523 14090
rect 16708 13994 16804 14010
rect 16708 13930 16724 13994
rect 16788 13930 16804 13994
rect 16708 13914 16804 13930
rect 16708 13850 16724 13914
rect 16788 13850 16804 13914
rect 16708 13834 16804 13850
rect 16708 13770 16724 13834
rect 16788 13770 16804 13834
rect 16708 13754 16804 13770
rect 16248 13482 16568 13721
rect 16708 13690 16724 13754
rect 16788 13690 16804 13754
rect 16967 14034 17289 14043
rect 16967 13730 16976 14034
rect 17280 13730 17289 14034
rect 16967 13721 17289 13730
rect 17427 14010 17443 14074
rect 17507 14010 17523 14074
rect 17688 14043 18008 14421
rect 18146 14710 18162 14774
rect 18226 14710 18242 14774
rect 18865 14854 18961 14870
rect 18865 14790 18881 14854
rect 18945 14790 18961 14854
rect 18865 14774 18961 14790
rect 18408 14743 18728 14762
rect 18146 14694 18242 14710
rect 18146 14630 18162 14694
rect 18226 14630 18242 14694
rect 18146 14614 18242 14630
rect 18146 14550 18162 14614
rect 18226 14550 18242 14614
rect 18146 14534 18242 14550
rect 18146 14470 18162 14534
rect 18226 14470 18242 14534
rect 18146 14454 18242 14470
rect 18146 14390 18162 14454
rect 18226 14390 18242 14454
rect 18405 14734 18728 14743
rect 18405 14430 18414 14734
rect 18718 14430 18728 14734
rect 18405 14421 18728 14430
rect 18146 14374 18242 14390
rect 18146 14310 18162 14374
rect 18226 14310 18242 14374
rect 18146 14294 18242 14310
rect 17427 13994 17523 14010
rect 17427 13930 17443 13994
rect 17507 13930 17523 13994
rect 17427 13914 17523 13930
rect 17427 13850 17443 13914
rect 17507 13850 17523 13914
rect 17427 13834 17523 13850
rect 17427 13770 17443 13834
rect 17507 13770 17523 13834
rect 17427 13754 17523 13770
rect 16708 13674 16804 13690
rect 16708 13610 16724 13674
rect 16788 13610 16804 13674
rect 16708 13594 16804 13610
rect 16968 13482 17288 13721
rect 17427 13690 17443 13754
rect 17507 13690 17523 13754
rect 17686 14034 18008 14043
rect 17686 13730 17695 14034
rect 17999 13730 18008 14034
rect 17686 13721 18008 13730
rect 17427 13674 17523 13690
rect 17427 13610 17443 13674
rect 17507 13610 17523 13674
rect 17427 13594 17523 13610
rect 17688 13482 18008 13721
rect 18146 14154 18242 14170
rect 18146 14090 18162 14154
rect 18226 14090 18242 14154
rect 18146 14074 18242 14090
rect 18146 14010 18162 14074
rect 18226 14010 18242 14074
rect 18408 14043 18728 14421
rect 18865 14710 18881 14774
rect 18945 14710 18961 14774
rect 19584 14854 19680 14870
rect 19584 14790 19600 14854
rect 19664 14790 19680 14854
rect 19584 14774 19680 14790
rect 19128 14743 19448 14762
rect 18865 14694 18961 14710
rect 18865 14630 18881 14694
rect 18945 14630 18961 14694
rect 18865 14614 18961 14630
rect 18865 14550 18881 14614
rect 18945 14550 18961 14614
rect 18865 14534 18961 14550
rect 18865 14470 18881 14534
rect 18945 14470 18961 14534
rect 18865 14454 18961 14470
rect 18865 14390 18881 14454
rect 18945 14390 18961 14454
rect 19124 14734 19448 14743
rect 19124 14430 19133 14734
rect 19437 14430 19448 14734
rect 19124 14421 19448 14430
rect 18865 14374 18961 14390
rect 18865 14310 18881 14374
rect 18945 14310 18961 14374
rect 18865 14294 18961 14310
rect 18146 13994 18242 14010
rect 18146 13930 18162 13994
rect 18226 13930 18242 13994
rect 18146 13914 18242 13930
rect 18146 13850 18162 13914
rect 18226 13850 18242 13914
rect 18146 13834 18242 13850
rect 18146 13770 18162 13834
rect 18226 13770 18242 13834
rect 18146 13754 18242 13770
rect 18146 13690 18162 13754
rect 18226 13690 18242 13754
rect 18405 14034 18728 14043
rect 18405 13730 18414 14034
rect 18718 13730 18728 14034
rect 18405 13721 18728 13730
rect 18146 13674 18242 13690
rect 18146 13610 18162 13674
rect 18226 13610 18242 13674
rect 18146 13594 18242 13610
rect 18408 13482 18728 13721
rect 18865 14154 18961 14170
rect 18865 14090 18881 14154
rect 18945 14090 18961 14154
rect 18865 14074 18961 14090
rect 18865 14010 18881 14074
rect 18945 14010 18961 14074
rect 19128 14043 19448 14421
rect 19584 14710 19600 14774
rect 19664 14710 19680 14774
rect 20303 14854 20399 14870
rect 20303 14790 20319 14854
rect 20383 14790 20399 14854
rect 20303 14774 20399 14790
rect 19848 14743 20168 14762
rect 19584 14694 19680 14710
rect 19584 14630 19600 14694
rect 19664 14630 19680 14694
rect 19584 14614 19680 14630
rect 19584 14550 19600 14614
rect 19664 14550 19680 14614
rect 19584 14534 19680 14550
rect 19584 14470 19600 14534
rect 19664 14470 19680 14534
rect 19584 14454 19680 14470
rect 19584 14390 19600 14454
rect 19664 14390 19680 14454
rect 19843 14734 20168 14743
rect 19843 14430 19852 14734
rect 20156 14430 20168 14734
rect 19843 14421 20168 14430
rect 19584 14374 19680 14390
rect 19584 14310 19600 14374
rect 19664 14310 19680 14374
rect 19584 14294 19680 14310
rect 18865 13994 18961 14010
rect 18865 13930 18881 13994
rect 18945 13930 18961 13994
rect 18865 13914 18961 13930
rect 18865 13850 18881 13914
rect 18945 13850 18961 13914
rect 18865 13834 18961 13850
rect 18865 13770 18881 13834
rect 18945 13770 18961 13834
rect 18865 13754 18961 13770
rect 18865 13690 18881 13754
rect 18945 13690 18961 13754
rect 19124 14034 19448 14043
rect 19124 13730 19133 14034
rect 19437 13730 19448 14034
rect 19124 13721 19448 13730
rect 18865 13674 18961 13690
rect 18865 13610 18881 13674
rect 18945 13610 18961 13674
rect 18865 13594 18961 13610
rect 19128 13482 19448 13721
rect 19584 14154 19680 14170
rect 19584 14090 19600 14154
rect 19664 14090 19680 14154
rect 19584 14074 19680 14090
rect 19584 14010 19600 14074
rect 19664 14010 19680 14074
rect 19848 14043 20168 14421
rect 20303 14710 20319 14774
rect 20383 14710 20399 14774
rect 21022 14854 21118 14870
rect 21022 14790 21038 14854
rect 21102 14790 21118 14854
rect 21022 14774 21118 14790
rect 20568 14743 20888 14762
rect 20303 14694 20399 14710
rect 20303 14630 20319 14694
rect 20383 14630 20399 14694
rect 20303 14614 20399 14630
rect 20303 14550 20319 14614
rect 20383 14550 20399 14614
rect 20303 14534 20399 14550
rect 20303 14470 20319 14534
rect 20383 14470 20399 14534
rect 20303 14454 20399 14470
rect 20303 14390 20319 14454
rect 20383 14390 20399 14454
rect 20562 14734 20888 14743
rect 20562 14430 20571 14734
rect 20875 14430 20888 14734
rect 20562 14421 20888 14430
rect 20303 14374 20399 14390
rect 20303 14310 20319 14374
rect 20383 14310 20399 14374
rect 20303 14294 20399 14310
rect 19584 13994 19680 14010
rect 19584 13930 19600 13994
rect 19664 13930 19680 13994
rect 19584 13914 19680 13930
rect 19584 13850 19600 13914
rect 19664 13850 19680 13914
rect 19584 13834 19680 13850
rect 19584 13770 19600 13834
rect 19664 13770 19680 13834
rect 19584 13754 19680 13770
rect 19584 13690 19600 13754
rect 19664 13690 19680 13754
rect 19843 14034 20168 14043
rect 19843 13730 19852 14034
rect 20156 13730 20168 14034
rect 19843 13721 20168 13730
rect 19584 13674 19680 13690
rect 19584 13610 19600 13674
rect 19664 13610 19680 13674
rect 19584 13594 19680 13610
rect 19848 13482 20168 13721
rect 20303 14154 20399 14170
rect 20303 14090 20319 14154
rect 20383 14090 20399 14154
rect 20303 14074 20399 14090
rect 20303 14010 20319 14074
rect 20383 14010 20399 14074
rect 20568 14043 20888 14421
rect 21022 14710 21038 14774
rect 21102 14710 21118 14774
rect 21741 14854 21837 14870
rect 21741 14790 21757 14854
rect 21821 14790 21837 14854
rect 21741 14774 21837 14790
rect 21288 14743 21608 14762
rect 21022 14694 21118 14710
rect 21022 14630 21038 14694
rect 21102 14630 21118 14694
rect 21022 14614 21118 14630
rect 21022 14550 21038 14614
rect 21102 14550 21118 14614
rect 21022 14534 21118 14550
rect 21022 14470 21038 14534
rect 21102 14470 21118 14534
rect 21022 14454 21118 14470
rect 21022 14390 21038 14454
rect 21102 14390 21118 14454
rect 21281 14734 21608 14743
rect 21281 14430 21290 14734
rect 21594 14430 21608 14734
rect 21281 14421 21608 14430
rect 21022 14374 21118 14390
rect 21022 14310 21038 14374
rect 21102 14310 21118 14374
rect 21022 14294 21118 14310
rect 20303 13994 20399 14010
rect 20303 13930 20319 13994
rect 20383 13930 20399 13994
rect 20303 13914 20399 13930
rect 20303 13850 20319 13914
rect 20383 13850 20399 13914
rect 20303 13834 20399 13850
rect 20303 13770 20319 13834
rect 20383 13770 20399 13834
rect 20303 13754 20399 13770
rect 20303 13690 20319 13754
rect 20383 13690 20399 13754
rect 20562 14034 20888 14043
rect 20562 13730 20571 14034
rect 20875 13730 20888 14034
rect 20562 13721 20888 13730
rect 20303 13674 20399 13690
rect 20303 13610 20319 13674
rect 20383 13610 20399 13674
rect 20303 13594 20399 13610
rect 20568 13482 20888 13721
rect 21022 14154 21118 14170
rect 21022 14090 21038 14154
rect 21102 14090 21118 14154
rect 21022 14074 21118 14090
rect 21022 14010 21038 14074
rect 21102 14010 21118 14074
rect 21288 14043 21608 14421
rect 21741 14710 21757 14774
rect 21821 14710 21837 14774
rect 22460 14854 22556 14870
rect 22460 14790 22476 14854
rect 22540 14790 22556 14854
rect 22460 14774 22556 14790
rect 22008 14743 22328 14762
rect 21741 14694 21837 14710
rect 21741 14630 21757 14694
rect 21821 14630 21837 14694
rect 21741 14614 21837 14630
rect 21741 14550 21757 14614
rect 21821 14550 21837 14614
rect 21741 14534 21837 14550
rect 21741 14470 21757 14534
rect 21821 14470 21837 14534
rect 21741 14454 21837 14470
rect 21741 14390 21757 14454
rect 21821 14390 21837 14454
rect 22000 14734 22328 14743
rect 22000 14430 22009 14734
rect 22313 14430 22328 14734
rect 22000 14421 22328 14430
rect 21741 14374 21837 14390
rect 21741 14310 21757 14374
rect 21821 14310 21837 14374
rect 21741 14294 21837 14310
rect 21022 13994 21118 14010
rect 21022 13930 21038 13994
rect 21102 13930 21118 13994
rect 21022 13914 21118 13930
rect 21022 13850 21038 13914
rect 21102 13850 21118 13914
rect 21022 13834 21118 13850
rect 21022 13770 21038 13834
rect 21102 13770 21118 13834
rect 21022 13754 21118 13770
rect 21022 13690 21038 13754
rect 21102 13690 21118 13754
rect 21281 14034 21608 14043
rect 21281 13730 21290 14034
rect 21594 13730 21608 14034
rect 21281 13721 21608 13730
rect 21022 13674 21118 13690
rect 21022 13610 21038 13674
rect 21102 13610 21118 13674
rect 21022 13594 21118 13610
rect 21288 13482 21608 13721
rect 21741 14154 21837 14170
rect 21741 14090 21757 14154
rect 21821 14090 21837 14154
rect 21741 14074 21837 14090
rect 21741 14010 21757 14074
rect 21821 14010 21837 14074
rect 22008 14043 22328 14421
rect 22460 14710 22476 14774
rect 22540 14710 22556 14774
rect 23179 14854 23275 14870
rect 23179 14790 23195 14854
rect 23259 14790 23275 14854
rect 23179 14774 23275 14790
rect 22728 14743 23048 14762
rect 22460 14694 22556 14710
rect 22460 14630 22476 14694
rect 22540 14630 22556 14694
rect 22460 14614 22556 14630
rect 22460 14550 22476 14614
rect 22540 14550 22556 14614
rect 22460 14534 22556 14550
rect 22460 14470 22476 14534
rect 22540 14470 22556 14534
rect 22460 14454 22556 14470
rect 22460 14390 22476 14454
rect 22540 14390 22556 14454
rect 22719 14734 23048 14743
rect 22719 14430 22728 14734
rect 23032 14430 23048 14734
rect 22719 14421 23048 14430
rect 22460 14374 22556 14390
rect 22460 14310 22476 14374
rect 22540 14310 22556 14374
rect 22460 14294 22556 14310
rect 21741 13994 21837 14010
rect 21741 13930 21757 13994
rect 21821 13930 21837 13994
rect 21741 13914 21837 13930
rect 21741 13850 21757 13914
rect 21821 13850 21837 13914
rect 21741 13834 21837 13850
rect 21741 13770 21757 13834
rect 21821 13770 21837 13834
rect 21741 13754 21837 13770
rect 21741 13690 21757 13754
rect 21821 13690 21837 13754
rect 22000 14034 22328 14043
rect 22000 13730 22009 14034
rect 22313 13730 22328 14034
rect 22000 13721 22328 13730
rect 21741 13674 21837 13690
rect 21741 13610 21757 13674
rect 21821 13610 21837 13674
rect 21741 13594 21837 13610
rect 22008 13482 22328 13721
rect 22460 14154 22556 14170
rect 22460 14090 22476 14154
rect 22540 14090 22556 14154
rect 22460 14074 22556 14090
rect 22460 14010 22476 14074
rect 22540 14010 22556 14074
rect 22728 14043 23048 14421
rect 23179 14710 23195 14774
rect 23259 14710 23275 14774
rect 23179 14694 23275 14710
rect 23179 14630 23195 14694
rect 23259 14630 23275 14694
rect 23179 14614 23275 14630
rect 23179 14550 23195 14614
rect 23259 14550 23275 14614
rect 23179 14534 23275 14550
rect 23179 14470 23195 14534
rect 23259 14470 23275 14534
rect 23179 14454 23275 14470
rect 23179 14390 23195 14454
rect 23259 14390 23275 14454
rect 23179 14374 23275 14390
rect 23179 14310 23195 14374
rect 23259 14310 23275 14374
rect 23179 14294 23275 14310
rect 22460 13994 22556 14010
rect 22460 13930 22476 13994
rect 22540 13930 22556 13994
rect 22460 13914 22556 13930
rect 22460 13850 22476 13914
rect 22540 13850 22556 13914
rect 22460 13834 22556 13850
rect 22460 13770 22476 13834
rect 22540 13770 22556 13834
rect 22460 13754 22556 13770
rect 22460 13690 22476 13754
rect 22540 13690 22556 13754
rect 22719 14034 23048 14043
rect 22719 13730 22728 14034
rect 23032 13730 23048 14034
rect 22719 13721 23048 13730
rect 22460 13674 22556 13690
rect 22460 13610 22476 13674
rect 22540 13610 22556 13674
rect 22460 13594 22556 13610
rect 22728 13482 23048 13721
rect 23179 14154 23275 14170
rect 23179 14090 23195 14154
rect 23259 14090 23275 14154
rect 23179 14074 23275 14090
rect 23179 14010 23195 14074
rect 23259 14010 23275 14074
rect 23179 13994 23275 14010
rect 23179 13930 23195 13994
rect 23259 13930 23275 13994
rect 23179 13914 23275 13930
rect 23179 13850 23195 13914
rect 23259 13850 23275 13914
rect 23179 13834 23275 13850
rect 23179 13770 23195 13834
rect 23259 13828 23275 13834
rect 23259 13770 23536 13828
rect 23179 13768 23536 13770
rect 23179 13754 23275 13768
rect 23179 13690 23195 13754
rect 23259 13690 23275 13754
rect 23179 13674 23275 13690
rect 23179 13610 23195 13674
rect 23259 13610 23275 13674
rect 23179 13594 23275 13610
rect 16110 13464 23278 13482
rect 16110 13454 17264 13464
rect 16110 13390 16138 13454
rect 16202 13390 16218 13454
rect 16282 13400 17264 13454
rect 17328 13400 23278 13464
rect 16282 13390 23278 13400
rect 16110 13362 23278 13390
rect 3348 11320 3372 11384
rect 3436 11320 3452 11384
rect 3516 11320 3532 11384
rect 3596 11320 3612 11384
rect 3676 11320 3692 11384
rect 3756 11320 3772 11384
rect 3836 11320 3852 11384
rect 3916 11320 3932 11384
rect 3996 11320 4012 11384
rect 4076 11320 4092 11384
rect 4156 11320 4172 11384
rect 4236 11320 4252 11384
rect 4316 11320 4332 11384
rect 4396 11320 4412 11384
rect 4476 11320 4492 11384
rect 4556 11320 4572 11384
rect 4636 11320 4652 11384
rect 4716 11320 4732 11384
rect 4796 11320 4812 11384
rect 4876 11320 4892 11384
rect 4956 11320 4980 11384
rect 3348 7624 4980 11320
rect 23476 11147 23536 13768
rect 43656 11384 45288 15080
rect 43656 11320 43680 11384
rect 43744 11320 43760 11384
rect 43824 11320 43840 11384
rect 43904 11320 43920 11384
rect 43984 11320 44000 11384
rect 44064 11320 44080 11384
rect 44144 11320 44160 11384
rect 44224 11320 44240 11384
rect 44304 11320 44320 11384
rect 44384 11320 44400 11384
rect 44464 11320 44480 11384
rect 44544 11320 44560 11384
rect 44624 11320 44640 11384
rect 44704 11320 44720 11384
rect 44784 11320 44800 11384
rect 44864 11320 44880 11384
rect 44944 11320 44960 11384
rect 45024 11320 45040 11384
rect 45104 11320 45120 11384
rect 45184 11320 45200 11384
rect 45264 11320 45288 11384
rect 23473 11146 23539 11147
rect 23473 11144 23474 11146
rect 23200 11110 23474 11144
rect 16708 11094 16804 11110
rect 16708 11030 16724 11094
rect 16788 11030 16804 11094
rect 16708 11014 16804 11030
rect 16248 10983 16568 11002
rect 16248 10974 16570 10983
rect 16248 10670 16257 10974
rect 16561 10670 16570 10974
rect 16248 10661 16570 10670
rect 16708 10950 16724 11014
rect 16788 10950 16804 11014
rect 17427 11094 17523 11110
rect 17427 11030 17443 11094
rect 17507 11030 17523 11094
rect 17427 11014 17523 11030
rect 16968 10983 17288 11002
rect 16708 10934 16804 10950
rect 16708 10870 16724 10934
rect 16788 10870 16804 10934
rect 16708 10854 16804 10870
rect 16708 10790 16724 10854
rect 16788 10790 16804 10854
rect 16708 10774 16804 10790
rect 16708 10710 16724 10774
rect 16788 10710 16804 10774
rect 16708 10694 16804 10710
rect 16248 10283 16568 10661
rect 16708 10630 16724 10694
rect 16788 10630 16804 10694
rect 16967 10974 17289 10983
rect 16967 10670 16976 10974
rect 17280 10670 17289 10974
rect 16967 10661 17289 10670
rect 17427 10950 17443 11014
rect 17507 10950 17523 11014
rect 18146 11094 18242 11110
rect 18146 11030 18162 11094
rect 18226 11030 18242 11094
rect 18146 11014 18242 11030
rect 17688 10983 18008 11002
rect 17427 10934 17523 10950
rect 17427 10870 17443 10934
rect 17507 10870 17523 10934
rect 17427 10854 17523 10870
rect 17427 10790 17443 10854
rect 17507 10790 17523 10854
rect 17427 10774 17523 10790
rect 17427 10710 17443 10774
rect 17507 10710 17523 10774
rect 17427 10694 17523 10710
rect 16708 10614 16804 10630
rect 16708 10550 16724 10614
rect 16788 10550 16804 10614
rect 16708 10534 16804 10550
rect 16708 10394 16804 10410
rect 16708 10330 16724 10394
rect 16788 10330 16804 10394
rect 16708 10314 16804 10330
rect 16248 10274 16570 10283
rect 16248 9970 16257 10274
rect 16561 9970 16570 10274
rect 16248 9961 16570 9970
rect 16708 10250 16724 10314
rect 16788 10250 16804 10314
rect 16968 10283 17288 10661
rect 17427 10630 17443 10694
rect 17507 10630 17523 10694
rect 17686 10974 18008 10983
rect 17686 10670 17695 10974
rect 17999 10670 18008 10974
rect 17686 10661 18008 10670
rect 17427 10614 17523 10630
rect 17427 10550 17443 10614
rect 17507 10550 17523 10614
rect 17427 10534 17523 10550
rect 17427 10394 17523 10410
rect 17427 10330 17443 10394
rect 17507 10330 17523 10394
rect 17427 10314 17523 10330
rect 16708 10234 16804 10250
rect 16708 10170 16724 10234
rect 16788 10170 16804 10234
rect 16708 10154 16804 10170
rect 16708 10090 16724 10154
rect 16788 10090 16804 10154
rect 16708 10074 16804 10090
rect 16708 10010 16724 10074
rect 16788 10010 16804 10074
rect 16708 9994 16804 10010
rect 16248 9722 16568 9961
rect 16708 9930 16724 9994
rect 16788 9930 16804 9994
rect 16967 10274 17289 10283
rect 16967 9970 16976 10274
rect 17280 9970 17289 10274
rect 16967 9961 17289 9970
rect 17427 10250 17443 10314
rect 17507 10250 17523 10314
rect 17688 10283 18008 10661
rect 18146 10950 18162 11014
rect 18226 10950 18242 11014
rect 18865 11094 18961 11110
rect 18865 11030 18881 11094
rect 18945 11030 18961 11094
rect 18865 11014 18961 11030
rect 18408 10983 18728 11002
rect 18146 10934 18242 10950
rect 18146 10870 18162 10934
rect 18226 10870 18242 10934
rect 18146 10854 18242 10870
rect 18146 10790 18162 10854
rect 18226 10790 18242 10854
rect 18146 10774 18242 10790
rect 18146 10710 18162 10774
rect 18226 10710 18242 10774
rect 18146 10694 18242 10710
rect 18146 10630 18162 10694
rect 18226 10630 18242 10694
rect 18405 10974 18728 10983
rect 18405 10670 18414 10974
rect 18718 10670 18728 10974
rect 18405 10661 18728 10670
rect 18146 10614 18242 10630
rect 18146 10550 18162 10614
rect 18226 10550 18242 10614
rect 18146 10534 18242 10550
rect 17427 10234 17523 10250
rect 17427 10170 17443 10234
rect 17507 10170 17523 10234
rect 17427 10154 17523 10170
rect 17427 10090 17443 10154
rect 17507 10090 17523 10154
rect 17427 10074 17523 10090
rect 17427 10010 17443 10074
rect 17507 10010 17523 10074
rect 17427 9994 17523 10010
rect 16708 9914 16804 9930
rect 16708 9850 16724 9914
rect 16788 9850 16804 9914
rect 16708 9834 16804 9850
rect 16968 9722 17288 9961
rect 17427 9930 17443 9994
rect 17507 9930 17523 9994
rect 17686 10274 18008 10283
rect 17686 9970 17695 10274
rect 17999 9970 18008 10274
rect 17686 9961 18008 9970
rect 17427 9914 17523 9930
rect 17427 9850 17443 9914
rect 17507 9850 17523 9914
rect 17427 9834 17523 9850
rect 17688 9722 18008 9961
rect 18146 10394 18242 10410
rect 18146 10330 18162 10394
rect 18226 10330 18242 10394
rect 18146 10314 18242 10330
rect 18146 10250 18162 10314
rect 18226 10250 18242 10314
rect 18408 10283 18728 10661
rect 18865 10950 18881 11014
rect 18945 10950 18961 11014
rect 19584 11094 19680 11110
rect 19584 11030 19600 11094
rect 19664 11030 19680 11094
rect 19584 11014 19680 11030
rect 19128 10983 19448 11002
rect 18865 10934 18961 10950
rect 18865 10870 18881 10934
rect 18945 10870 18961 10934
rect 18865 10854 18961 10870
rect 18865 10790 18881 10854
rect 18945 10790 18961 10854
rect 18865 10774 18961 10790
rect 18865 10710 18881 10774
rect 18945 10710 18961 10774
rect 18865 10694 18961 10710
rect 18865 10630 18881 10694
rect 18945 10630 18961 10694
rect 19124 10974 19448 10983
rect 19124 10670 19133 10974
rect 19437 10670 19448 10974
rect 19124 10661 19448 10670
rect 18865 10614 18961 10630
rect 18865 10550 18881 10614
rect 18945 10550 18961 10614
rect 18865 10534 18961 10550
rect 18146 10234 18242 10250
rect 18146 10170 18162 10234
rect 18226 10170 18242 10234
rect 18146 10154 18242 10170
rect 18146 10090 18162 10154
rect 18226 10090 18242 10154
rect 18146 10074 18242 10090
rect 18146 10010 18162 10074
rect 18226 10010 18242 10074
rect 18146 9994 18242 10010
rect 18146 9930 18162 9994
rect 18226 9930 18242 9994
rect 18405 10274 18728 10283
rect 18405 9970 18414 10274
rect 18718 9970 18728 10274
rect 18405 9961 18728 9970
rect 18146 9914 18242 9930
rect 18146 9850 18162 9914
rect 18226 9850 18242 9914
rect 18146 9834 18242 9850
rect 18408 9722 18728 9961
rect 18865 10394 18961 10410
rect 18865 10330 18881 10394
rect 18945 10330 18961 10394
rect 18865 10314 18961 10330
rect 18865 10250 18881 10314
rect 18945 10250 18961 10314
rect 19128 10283 19448 10661
rect 19584 10950 19600 11014
rect 19664 10950 19680 11014
rect 20303 11094 20399 11110
rect 20303 11030 20319 11094
rect 20383 11030 20399 11094
rect 20303 11014 20399 11030
rect 19848 10983 20168 11002
rect 19584 10934 19680 10950
rect 19584 10870 19600 10934
rect 19664 10870 19680 10934
rect 19584 10854 19680 10870
rect 19584 10790 19600 10854
rect 19664 10790 19680 10854
rect 19584 10774 19680 10790
rect 19584 10710 19600 10774
rect 19664 10710 19680 10774
rect 19584 10694 19680 10710
rect 19584 10630 19600 10694
rect 19664 10630 19680 10694
rect 19843 10974 20168 10983
rect 19843 10670 19852 10974
rect 20156 10670 20168 10974
rect 19843 10661 20168 10670
rect 19584 10614 19680 10630
rect 19584 10550 19600 10614
rect 19664 10550 19680 10614
rect 19584 10534 19680 10550
rect 18865 10234 18961 10250
rect 18865 10170 18881 10234
rect 18945 10170 18961 10234
rect 18865 10154 18961 10170
rect 18865 10090 18881 10154
rect 18945 10090 18961 10154
rect 18865 10074 18961 10090
rect 18865 10010 18881 10074
rect 18945 10010 18961 10074
rect 18865 9994 18961 10010
rect 18865 9930 18881 9994
rect 18945 9930 18961 9994
rect 19124 10274 19448 10283
rect 19124 9970 19133 10274
rect 19437 9970 19448 10274
rect 19124 9961 19448 9970
rect 18865 9914 18961 9930
rect 18865 9850 18881 9914
rect 18945 9850 18961 9914
rect 18865 9834 18961 9850
rect 19128 9722 19448 9961
rect 19584 10394 19680 10410
rect 19584 10330 19600 10394
rect 19664 10330 19680 10394
rect 19584 10314 19680 10330
rect 19584 10250 19600 10314
rect 19664 10250 19680 10314
rect 19848 10283 20168 10661
rect 20303 10950 20319 11014
rect 20383 10950 20399 11014
rect 21022 11094 21118 11110
rect 21022 11030 21038 11094
rect 21102 11030 21118 11094
rect 21022 11014 21118 11030
rect 20568 10983 20888 11002
rect 20303 10934 20399 10950
rect 20303 10870 20319 10934
rect 20383 10870 20399 10934
rect 20303 10854 20399 10870
rect 20303 10790 20319 10854
rect 20383 10790 20399 10854
rect 20303 10774 20399 10790
rect 20303 10710 20319 10774
rect 20383 10710 20399 10774
rect 20303 10694 20399 10710
rect 20303 10630 20319 10694
rect 20383 10630 20399 10694
rect 20562 10974 20888 10983
rect 20562 10670 20571 10974
rect 20875 10670 20888 10974
rect 20562 10661 20888 10670
rect 20303 10614 20399 10630
rect 20303 10550 20319 10614
rect 20383 10550 20399 10614
rect 20303 10534 20399 10550
rect 19584 10234 19680 10250
rect 19584 10170 19600 10234
rect 19664 10170 19680 10234
rect 19584 10154 19680 10170
rect 19584 10090 19600 10154
rect 19664 10090 19680 10154
rect 19584 10074 19680 10090
rect 19584 10010 19600 10074
rect 19664 10010 19680 10074
rect 19584 9994 19680 10010
rect 19584 9930 19600 9994
rect 19664 9930 19680 9994
rect 19843 10274 20168 10283
rect 19843 9970 19852 10274
rect 20156 9970 20168 10274
rect 19843 9961 20168 9970
rect 19584 9914 19680 9930
rect 19584 9850 19600 9914
rect 19664 9850 19680 9914
rect 19584 9834 19680 9850
rect 19848 9722 20168 9961
rect 20303 10394 20399 10410
rect 20303 10330 20319 10394
rect 20383 10330 20399 10394
rect 20303 10314 20399 10330
rect 20303 10250 20319 10314
rect 20383 10250 20399 10314
rect 20568 10283 20888 10661
rect 21022 10950 21038 11014
rect 21102 10950 21118 11014
rect 21741 11094 21837 11110
rect 21741 11030 21757 11094
rect 21821 11030 21837 11094
rect 21741 11014 21837 11030
rect 21288 10983 21608 11002
rect 21022 10934 21118 10950
rect 21022 10870 21038 10934
rect 21102 10870 21118 10934
rect 21022 10854 21118 10870
rect 21022 10790 21038 10854
rect 21102 10790 21118 10854
rect 21022 10774 21118 10790
rect 21022 10710 21038 10774
rect 21102 10710 21118 10774
rect 21022 10694 21118 10710
rect 21022 10630 21038 10694
rect 21102 10630 21118 10694
rect 21281 10974 21608 10983
rect 21281 10670 21290 10974
rect 21594 10670 21608 10974
rect 21281 10661 21608 10670
rect 21022 10614 21118 10630
rect 21022 10550 21038 10614
rect 21102 10550 21118 10614
rect 21022 10534 21118 10550
rect 20303 10234 20399 10250
rect 20303 10170 20319 10234
rect 20383 10170 20399 10234
rect 20303 10154 20399 10170
rect 20303 10090 20319 10154
rect 20383 10090 20399 10154
rect 20303 10074 20399 10090
rect 20303 10010 20319 10074
rect 20383 10010 20399 10074
rect 20303 9994 20399 10010
rect 20303 9930 20319 9994
rect 20383 9930 20399 9994
rect 20562 10274 20888 10283
rect 20562 9970 20571 10274
rect 20875 9970 20888 10274
rect 20562 9961 20888 9970
rect 20303 9914 20399 9930
rect 20303 9850 20319 9914
rect 20383 9850 20399 9914
rect 20303 9834 20399 9850
rect 20568 9722 20888 9961
rect 21022 10394 21118 10410
rect 21022 10330 21038 10394
rect 21102 10330 21118 10394
rect 21022 10314 21118 10330
rect 21022 10250 21038 10314
rect 21102 10250 21118 10314
rect 21288 10283 21608 10661
rect 21741 10950 21757 11014
rect 21821 10950 21837 11014
rect 22460 11094 22556 11110
rect 22460 11030 22476 11094
rect 22540 11030 22556 11094
rect 22460 11014 22556 11030
rect 22008 10983 22328 11002
rect 21741 10934 21837 10950
rect 21741 10870 21757 10934
rect 21821 10870 21837 10934
rect 21741 10854 21837 10870
rect 21741 10790 21757 10854
rect 21821 10790 21837 10854
rect 21741 10774 21837 10790
rect 21741 10710 21757 10774
rect 21821 10710 21837 10774
rect 21741 10694 21837 10710
rect 21741 10630 21757 10694
rect 21821 10630 21837 10694
rect 22000 10974 22328 10983
rect 22000 10670 22009 10974
rect 22313 10670 22328 10974
rect 22000 10661 22328 10670
rect 21741 10614 21837 10630
rect 21741 10550 21757 10614
rect 21821 10550 21837 10614
rect 21741 10534 21837 10550
rect 21022 10234 21118 10250
rect 21022 10170 21038 10234
rect 21102 10170 21118 10234
rect 21022 10154 21118 10170
rect 21022 10090 21038 10154
rect 21102 10090 21118 10154
rect 21022 10074 21118 10090
rect 21022 10010 21038 10074
rect 21102 10010 21118 10074
rect 21022 9994 21118 10010
rect 21022 9930 21038 9994
rect 21102 9930 21118 9994
rect 21281 10274 21608 10283
rect 21281 9970 21290 10274
rect 21594 9970 21608 10274
rect 21281 9961 21608 9970
rect 21022 9914 21118 9930
rect 21022 9850 21038 9914
rect 21102 9850 21118 9914
rect 21022 9834 21118 9850
rect 21288 9722 21608 9961
rect 21741 10394 21837 10410
rect 21741 10330 21757 10394
rect 21821 10330 21837 10394
rect 21741 10314 21837 10330
rect 21741 10250 21757 10314
rect 21821 10250 21837 10314
rect 22008 10283 22328 10661
rect 22460 10950 22476 11014
rect 22540 10950 22556 11014
rect 23179 11094 23474 11110
rect 23179 11030 23195 11094
rect 23259 11084 23474 11094
rect 23259 11030 23275 11084
rect 23473 11082 23474 11084
rect 23538 11082 23539 11146
rect 23473 11081 23539 11082
rect 23179 11014 23275 11030
rect 22728 10983 23048 11002
rect 22460 10934 22556 10950
rect 22460 10870 22476 10934
rect 22540 10870 22556 10934
rect 22460 10854 22556 10870
rect 22460 10790 22476 10854
rect 22540 10790 22556 10854
rect 22460 10774 22556 10790
rect 22460 10710 22476 10774
rect 22540 10710 22556 10774
rect 22460 10694 22556 10710
rect 22460 10630 22476 10694
rect 22540 10630 22556 10694
rect 22719 10974 23048 10983
rect 22719 10670 22728 10974
rect 23032 10670 23048 10974
rect 22719 10661 23048 10670
rect 22460 10614 22556 10630
rect 22460 10550 22476 10614
rect 22540 10550 22556 10614
rect 22460 10534 22556 10550
rect 21741 10234 21837 10250
rect 21741 10170 21757 10234
rect 21821 10170 21837 10234
rect 21741 10154 21837 10170
rect 21741 10090 21757 10154
rect 21821 10090 21837 10154
rect 21741 10074 21837 10090
rect 21741 10010 21757 10074
rect 21821 10010 21837 10074
rect 21741 9994 21837 10010
rect 21741 9930 21757 9994
rect 21821 9930 21837 9994
rect 22000 10274 22328 10283
rect 22000 9970 22009 10274
rect 22313 9970 22328 10274
rect 22000 9961 22328 9970
rect 21741 9914 21837 9930
rect 21741 9850 21757 9914
rect 21821 9850 21837 9914
rect 21741 9834 21837 9850
rect 22008 9722 22328 9961
rect 22460 10394 22556 10410
rect 22460 10330 22476 10394
rect 22540 10330 22556 10394
rect 22460 10314 22556 10330
rect 22460 10250 22476 10314
rect 22540 10250 22556 10314
rect 22728 10283 23048 10661
rect 23179 10950 23195 11014
rect 23259 10950 23275 11014
rect 23179 10934 23275 10950
rect 23179 10870 23195 10934
rect 23259 10870 23275 10934
rect 23179 10854 23275 10870
rect 23179 10790 23195 10854
rect 23259 10790 23275 10854
rect 23179 10774 23275 10790
rect 23179 10710 23195 10774
rect 23259 10710 23275 10774
rect 23179 10694 23275 10710
rect 23179 10630 23195 10694
rect 23259 10630 23275 10694
rect 23179 10614 23275 10630
rect 23179 10550 23195 10614
rect 23259 10550 23275 10614
rect 23179 10534 23275 10550
rect 22460 10234 22556 10250
rect 22460 10170 22476 10234
rect 22540 10170 22556 10234
rect 22460 10154 22556 10170
rect 22460 10090 22476 10154
rect 22540 10090 22556 10154
rect 22460 10074 22556 10090
rect 22460 10010 22476 10074
rect 22540 10010 22556 10074
rect 22460 9994 22556 10010
rect 22460 9930 22476 9994
rect 22540 9930 22556 9994
rect 22719 10274 23048 10283
rect 22719 9970 22728 10274
rect 23032 9970 23048 10274
rect 22719 9961 23048 9970
rect 22460 9914 22556 9930
rect 22460 9850 22476 9914
rect 22540 9850 22556 9914
rect 22460 9834 22556 9850
rect 22728 9722 23048 9961
rect 23179 10394 23275 10410
rect 23179 10330 23195 10394
rect 23259 10330 23275 10394
rect 23179 10314 23275 10330
rect 23179 10250 23195 10314
rect 23259 10250 23275 10314
rect 23179 10234 23275 10250
rect 23179 10170 23195 10234
rect 23259 10170 23275 10234
rect 23179 10154 23275 10170
rect 23179 10090 23195 10154
rect 23259 10090 23275 10154
rect 23179 10074 23275 10090
rect 23179 10010 23195 10074
rect 23259 10010 23275 10074
rect 23179 9994 23275 10010
rect 23179 9930 23195 9994
rect 23259 9930 23275 9994
rect 23179 9914 23275 9930
rect 23179 9850 23195 9914
rect 23259 9850 23275 9914
rect 23179 9834 23275 9850
rect 16110 9694 23278 9722
rect 16110 9630 16138 9694
rect 16202 9630 16218 9694
rect 16282 9682 23278 9694
rect 16282 9630 17264 9682
rect 16110 9618 17264 9630
rect 17328 9618 23278 9682
rect 16110 9602 23278 9618
rect 3348 7560 3372 7624
rect 3436 7560 3452 7624
rect 3516 7560 3532 7624
rect 3596 7560 3612 7624
rect 3676 7560 3692 7624
rect 3756 7560 3772 7624
rect 3836 7560 3852 7624
rect 3916 7560 3932 7624
rect 3996 7560 4012 7624
rect 4076 7560 4092 7624
rect 4156 7560 4172 7624
rect 4236 7560 4252 7624
rect 4316 7560 4332 7624
rect 4396 7560 4412 7624
rect 4476 7560 4492 7624
rect 4556 7560 4572 7624
rect 4636 7560 4652 7624
rect 4716 7560 4732 7624
rect 4796 7560 4812 7624
rect 4876 7560 4892 7624
rect 4956 7560 4980 7624
rect 3348 4838 4980 7560
rect 3348 3322 3406 4838
rect 4922 3322 4980 4838
rect 3348 0 4980 3322
rect 43656 7624 45288 11320
rect 43656 7560 43680 7624
rect 43744 7560 43760 7624
rect 43824 7560 43840 7624
rect 43904 7560 43920 7624
rect 43984 7560 44000 7624
rect 44064 7560 44080 7624
rect 44144 7560 44160 7624
rect 44224 7560 44240 7624
rect 44304 7560 44320 7624
rect 44384 7560 44400 7624
rect 44464 7560 44480 7624
rect 44544 7560 44560 7624
rect 44624 7560 44640 7624
rect 44704 7560 44720 7624
rect 44784 7560 44800 7624
rect 44864 7560 44880 7624
rect 44944 7560 44960 7624
rect 45024 7560 45040 7624
rect 45104 7560 45120 7624
rect 45184 7560 45200 7624
rect 45264 7560 45288 7624
rect 43656 4838 45288 7560
rect 43656 3322 43714 4838
rect 45230 3322 45288 4838
rect 43656 0 45288 3322
rect 46104 46270 47736 47192
rect 46104 44754 46162 46270
rect 47678 44754 47736 46270
rect 46104 39584 47736 44754
rect 46104 39520 46128 39584
rect 46192 39520 46208 39584
rect 46272 39520 46288 39584
rect 46352 39520 46368 39584
rect 46432 39520 46448 39584
rect 46512 39520 46528 39584
rect 46592 39520 46608 39584
rect 46672 39520 46688 39584
rect 46752 39520 46768 39584
rect 46832 39520 46848 39584
rect 46912 39520 46928 39584
rect 46992 39520 47008 39584
rect 47072 39520 47088 39584
rect 47152 39520 47168 39584
rect 47232 39520 47248 39584
rect 47312 39520 47328 39584
rect 47392 39520 47408 39584
rect 47472 39520 47488 39584
rect 47552 39520 47568 39584
rect 47632 39520 47648 39584
rect 47712 39520 47736 39584
rect 46104 35824 47736 39520
rect 46104 35760 46128 35824
rect 46192 35760 46208 35824
rect 46272 35760 46288 35824
rect 46352 35760 46368 35824
rect 46432 35760 46448 35824
rect 46512 35760 46528 35824
rect 46592 35760 46608 35824
rect 46672 35760 46688 35824
rect 46752 35760 46768 35824
rect 46832 35760 46848 35824
rect 46912 35760 46928 35824
rect 46992 35760 47008 35824
rect 47072 35760 47088 35824
rect 47152 35760 47168 35824
rect 47232 35760 47248 35824
rect 47312 35760 47328 35824
rect 47392 35760 47408 35824
rect 47472 35760 47488 35824
rect 47552 35760 47568 35824
rect 47632 35760 47648 35824
rect 47712 35760 47736 35824
rect 46104 32064 47736 35760
rect 46104 32000 46128 32064
rect 46192 32000 46208 32064
rect 46272 32000 46288 32064
rect 46352 32000 46368 32064
rect 46432 32000 46448 32064
rect 46512 32000 46528 32064
rect 46592 32000 46608 32064
rect 46672 32000 46688 32064
rect 46752 32000 46768 32064
rect 46832 32000 46848 32064
rect 46912 32000 46928 32064
rect 46992 32000 47008 32064
rect 47072 32000 47088 32064
rect 47152 32000 47168 32064
rect 47232 32000 47248 32064
rect 47312 32000 47328 32064
rect 47392 32000 47408 32064
rect 47472 32000 47488 32064
rect 47552 32000 47568 32064
rect 47632 32000 47648 32064
rect 47712 32000 47736 32064
rect 46104 28304 47736 32000
rect 46104 28240 46128 28304
rect 46192 28240 46208 28304
rect 46272 28240 46288 28304
rect 46352 28240 46368 28304
rect 46432 28240 46448 28304
rect 46512 28240 46528 28304
rect 46592 28240 46608 28304
rect 46672 28240 46688 28304
rect 46752 28240 46768 28304
rect 46832 28240 46848 28304
rect 46912 28240 46928 28304
rect 46992 28240 47008 28304
rect 47072 28240 47088 28304
rect 47152 28240 47168 28304
rect 47232 28240 47248 28304
rect 47312 28240 47328 28304
rect 47392 28240 47408 28304
rect 47472 28240 47488 28304
rect 47552 28240 47568 28304
rect 47632 28240 47648 28304
rect 47712 28240 47736 28304
rect 46104 24544 47736 28240
rect 46104 24480 46128 24544
rect 46192 24480 46208 24544
rect 46272 24480 46288 24544
rect 46352 24480 46368 24544
rect 46432 24480 46448 24544
rect 46512 24480 46528 24544
rect 46592 24480 46608 24544
rect 46672 24480 46688 24544
rect 46752 24480 46768 24544
rect 46832 24480 46848 24544
rect 46912 24480 46928 24544
rect 46992 24480 47008 24544
rect 47072 24480 47088 24544
rect 47152 24480 47168 24544
rect 47232 24480 47248 24544
rect 47312 24480 47328 24544
rect 47392 24480 47408 24544
rect 47472 24480 47488 24544
rect 47552 24480 47568 24544
rect 47632 24480 47648 24544
rect 47712 24480 47736 24544
rect 46104 20784 47736 24480
rect 46104 20720 46128 20784
rect 46192 20720 46208 20784
rect 46272 20720 46288 20784
rect 46352 20720 46368 20784
rect 46432 20720 46448 20784
rect 46512 20720 46528 20784
rect 46592 20720 46608 20784
rect 46672 20720 46688 20784
rect 46752 20720 46768 20784
rect 46832 20720 46848 20784
rect 46912 20720 46928 20784
rect 46992 20720 47008 20784
rect 47072 20720 47088 20784
rect 47152 20720 47168 20784
rect 47232 20720 47248 20784
rect 47312 20720 47328 20784
rect 47392 20720 47408 20784
rect 47472 20720 47488 20784
rect 47552 20720 47568 20784
rect 47632 20720 47648 20784
rect 47712 20720 47736 20784
rect 46104 17024 47736 20720
rect 46104 16960 46128 17024
rect 46192 16960 46208 17024
rect 46272 16960 46288 17024
rect 46352 16960 46368 17024
rect 46432 16960 46448 17024
rect 46512 16960 46528 17024
rect 46592 16960 46608 17024
rect 46672 16960 46688 17024
rect 46752 16960 46768 17024
rect 46832 16960 46848 17024
rect 46912 16960 46928 17024
rect 46992 16960 47008 17024
rect 47072 16960 47088 17024
rect 47152 16960 47168 17024
rect 47232 16960 47248 17024
rect 47312 16960 47328 17024
rect 47392 16960 47408 17024
rect 47472 16960 47488 17024
rect 47552 16960 47568 17024
rect 47632 16960 47648 17024
rect 47712 16960 47736 17024
rect 46104 13264 47736 16960
rect 46104 13200 46128 13264
rect 46192 13200 46208 13264
rect 46272 13200 46288 13264
rect 46352 13200 46368 13264
rect 46432 13200 46448 13264
rect 46512 13200 46528 13264
rect 46592 13200 46608 13264
rect 46672 13200 46688 13264
rect 46752 13200 46768 13264
rect 46832 13200 46848 13264
rect 46912 13200 46928 13264
rect 46992 13200 47008 13264
rect 47072 13200 47088 13264
rect 47152 13200 47168 13264
rect 47232 13200 47248 13264
rect 47312 13200 47328 13264
rect 47392 13200 47408 13264
rect 47472 13200 47488 13264
rect 47552 13200 47568 13264
rect 47632 13200 47648 13264
rect 47712 13200 47736 13264
rect 46104 9504 47736 13200
rect 46104 9440 46128 9504
rect 46192 9440 46208 9504
rect 46272 9440 46288 9504
rect 46352 9440 46368 9504
rect 46432 9440 46448 9504
rect 46512 9440 46528 9504
rect 46592 9440 46608 9504
rect 46672 9440 46688 9504
rect 46752 9440 46768 9504
rect 46832 9440 46848 9504
rect 46912 9440 46928 9504
rect 46992 9440 47008 9504
rect 47072 9440 47088 9504
rect 47152 9440 47168 9504
rect 47232 9440 47248 9504
rect 47312 9440 47328 9504
rect 47392 9440 47408 9504
rect 47472 9440 47488 9504
rect 47552 9440 47568 9504
rect 47632 9440 47648 9504
rect 47712 9440 47736 9504
rect 46104 5744 47736 9440
rect 46104 5680 46128 5744
rect 46192 5680 46208 5744
rect 46272 5680 46288 5744
rect 46352 5680 46368 5744
rect 46432 5680 46448 5744
rect 46512 5680 46528 5744
rect 46592 5680 46608 5744
rect 46672 5680 46688 5744
rect 46752 5680 46768 5744
rect 46832 5680 46848 5744
rect 46912 5680 46928 5744
rect 46992 5680 47008 5744
rect 47072 5680 47088 5744
rect 47152 5680 47168 5744
rect 47232 5680 47248 5744
rect 47312 5680 47328 5744
rect 47392 5680 47408 5744
rect 47472 5680 47488 5744
rect 47552 5680 47568 5744
rect 47632 5680 47648 5744
rect 47712 5680 47736 5744
rect 46104 2390 47736 5680
rect 46104 874 46162 2390
rect 47678 874 47736 2390
rect 46104 0 47736 874
<< via4 >>
rect 958 44754 2474 46270
rect 958 874 2474 2390
rect 3406 42306 4922 43822
rect 43714 42306 45230 43822
rect 3406 3322 4922 4838
rect 43714 3322 45230 4838
rect 46162 44754 47678 46270
rect 46162 874 47678 2390
<< metal5 >>
rect 0 46270 48668 46328
rect 0 44754 958 46270
rect 2474 44754 46162 46270
rect 47678 44754 48668 46270
rect 0 44696 48668 44754
rect 0 43822 48668 43880
rect 0 42306 3406 43822
rect 4922 42306 43714 43822
rect 45230 42306 48668 43822
rect 0 42248 48668 42306
rect 0 4838 48668 4896
rect 0 3322 3406 4838
rect 4922 3322 43714 4838
rect 45230 3322 48668 4838
rect 0 3264 48668 3322
rect 0 2390 48668 2448
rect 0 874 958 2390
rect 2474 874 46162 2390
rect 47678 874 48668 2390
rect 0 816 48668 874
<< labels >>
rlabel metal1 s 0 17292 119 17320 4 porst
port 1 nsew
rlabel metal2 s 27448 47095 27476 47192 4 vbg
port 2 nsew
rlabel metal5 s 0 816 1632 2448 4 VSS
port 3 nsew
rlabel metal5 s 0 3264 1632 4896 4 VDD
port 4 nsew
flabel metal1 8016 7012 8136 7132 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_1/Rin
flabel metal1 8016 6052 8136 6172 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_1/Rout
flabel metal1 7896 7562 7956 7622 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_1/VPWR
flabel metal1 7896 5682 7956 5742 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_1/VGND
flabel metal1 14387 7012 14507 7132 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_2_1/Rin
flabel metal1 14387 6052 14507 6172 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_2_1/Rout
flabel metal1 14268 7562 14328 7622 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_2_1/VPWR
flabel metal1 14268 5682 14328 5742 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_2_1/VGND
flabel metal1 17718 7012 17838 7132 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_27/Rin
flabel metal1 17718 6052 17838 6172 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_27/Rout
flabel metal1 17598 7562 17658 7622 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_27/VPWR
flabel metal1 17598 5682 17658 5742 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_27/VGND
flabel metal1 20462 7012 20582 7132 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_25/Rin
flabel metal1 20462 6052 20582 6172 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_25/Rout
flabel metal1 20342 7562 20402 7622 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_25/VPWR
flabel metal1 20342 5682 20402 5742 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_25/VGND
flabel metal1 23206 7012 23326 7132 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_23/Rin
flabel metal1 23206 6052 23326 6172 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_23/Rout
flabel metal1 23086 7562 23146 7622 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_23/VPWR
flabel metal1 23086 5682 23146 5742 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_23/VGND
flabel metal1 25950 7012 26070 7132 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_26/Rin
flabel metal1 25950 6052 26070 6172 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_26/Rout
flabel metal1 25830 7562 25890 7622 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_26/VPWR
flabel metal1 25830 5682 25890 5742 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_26/VGND
flabel metal1 28694 7012 28814 7132 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_28/Rin
flabel metal1 28694 6052 28814 6172 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_28/Rout
flabel metal1 28574 7562 28634 7622 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_28/VPWR
flabel metal1 28574 5682 28634 5742 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_28/VGND
flabel metal1 31438 7012 31558 7132 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_13/Rin
flabel metal1 31438 6052 31558 6172 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_13/Rout
flabel metal1 31318 7562 31378 7622 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_13/VPWR
flabel metal1 31318 5682 31378 5742 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_13/VGND
flabel metal1 35260 7012 35380 7132 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_11/Rin
flabel metal1 35260 6052 35380 6172 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_11/Rout
flabel metal1 35140 7562 35200 7622 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_11/VPWR
flabel metal1 35140 5682 35200 5742 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_11/VGND
flabel metal1 38004 7012 38124 7132 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_15/Rin
flabel metal1 38004 6052 38124 6172 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_15/Rout
flabel metal1 37884 7562 37944 7622 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_15/VPWR
flabel metal1 37884 5682 37944 5742 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_15/VGND
flabel metal1 8016 10772 8136 10892 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_3/Rin
flabel metal1 8016 9812 8136 9932 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_3/Rout
flabel metal1 7896 11322 7956 11382 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_3/VPWR
flabel metal1 7896 9442 7956 9502 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_3/VGND
flabel metal1 10760 10772 10880 10892 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_24/Rin
flabel metal1 10760 9812 10880 9932 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_24/Rout
flabel metal1 10640 11322 10700 11382 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_24/VPWR
flabel metal1 10640 9442 10700 9502 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_24/VGND
flabel metal1 13504 10772 13624 10892 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_21/Rin
flabel metal1 13504 9812 13624 9932 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_21/Rout
flabel metal1 13384 11322 13444 11382 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_21/VPWR
flabel metal1 13384 9442 13444 9502 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_21/VGND
flabel metal2 16108 11042 16308 11122 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_8/Cin
flabel metal4 16130 9612 16290 9712 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_8/Cout
flabel metal1 16110 11322 16170 11382 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_8/VPWR
flabel metal1 16110 9442 16170 9502 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_8/VGND
flabel metal1 23697 10772 23817 10892 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_2_0/Rin
flabel metal1 23697 9812 23817 9932 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_2_0/Rout
flabel metal1 23578 11322 23638 11382 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_2_0/VPWR
flabel metal1 23578 9442 23638 9502 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_2_0/VGND
flabel metal1 27028 10772 27148 10892 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_29/Rin
flabel metal1 27028 9812 27148 9932 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_29/Rout
flabel metal1 26908 11322 26968 11382 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_29/VPWR
flabel metal1 26908 9442 26968 9502 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_29/VGND
flabel metal1 29772 10772 29892 10892 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_30/Rin
flabel metal1 29772 9812 29892 9932 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_30/Rout
flabel metal1 29652 11322 29712 11382 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_30/VPWR
flabel metal1 29652 9442 29712 9502 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_30/VGND
flabel metal1 35260 10772 35380 10892 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_14/Rin
flabel metal1 35260 9812 35380 9932 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_14/Rout
flabel metal1 35140 11322 35200 11382 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_14/VPWR
flabel metal1 35140 9442 35200 9502 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_14/VGND
flabel metal1 32516 10772 32636 10892 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_10/Rin
flabel metal1 32516 9812 32636 9932 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_10/Rout
flabel metal1 32396 11322 32456 11382 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_10/VPWR
flabel metal1 32396 9442 32456 9502 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_10/VGND
flabel metal1 38004 10772 38124 10892 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_12/Rin
flabel metal1 38004 9812 38124 9932 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_12/Rout
flabel metal1 37884 11322 37944 11382 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_12/VPWR
flabel metal1 37884 9442 37944 9502 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_12/VGND
flabel metal1 8016 14532 8136 14652 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_4/Rin
flabel metal1 8016 13572 8136 13692 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_4/Rout
flabel metal1 7896 15082 7956 15142 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_4/VPWR
flabel metal1 7896 13202 7956 13262 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_4/VGND
flabel metal1 10760 14532 10880 14652 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_2/Rin
flabel metal1 10760 13572 10880 13692 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_2/Rout
flabel metal1 10640 15082 10700 15142 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_2/VPWR
flabel metal1 10640 13202 10700 13262 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_2/VGND
flabel metal2 16108 14802 16308 14882 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_6/Cin
flabel metal4 16130 13372 16290 13472 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_6/Cout
flabel metal1 16110 15082 16170 15142 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_6/VPWR
flabel metal1 16110 13202 16170 13262 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_6/VGND
flabel metal1 13504 14532 13624 14652 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_9/Rin
flabel metal1 13504 13572 13624 13692 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_9/Rout
flabel metal1 13384 15082 13444 15142 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_9/VPWR
flabel metal1 13384 13202 13444 13262 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_9/VGND
flabel locali 38194 14128 38442 14232 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Emitter
flabel locali 38253 14754 38354 14803 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Collector
flabel locali 38230 14604 38348 14644 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Base
flabel locali 36854 14128 37102 14232 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Emitter
flabel locali 36913 14754 37014 14803 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector
flabel locali 36890 14604 37008 14644 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Base
flabel locali 35514 14128 35762 14232 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Emitter
flabel locali 35573 14754 35674 14803 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector
flabel locali 35550 14604 35668 14644 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Base
flabel locali 34174 14128 34422 14232 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Emitter
flabel locali 34233 14754 34334 14803 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector
flabel locali 34210 14604 34328 14644 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Base
flabel locali 32834 14128 33082 14232 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Emitter
flabel locali 32893 14754 32994 14803 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector
flabel locali 32870 14604 32988 14644 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Base
flabel locali 31494 14128 31742 14232 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Emitter
flabel locali 31553 14754 31654 14803 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector
flabel locali 31530 14604 31648 14644 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Base
flabel locali 30154 14128 30402 14232 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter
flabel locali 30213 14754 30314 14803 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector
flabel locali 30190 14604 30308 14644 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Base
flabel locali 28814 14128 29062 14232 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/xm1/Emitter
flabel locali 28873 14754 28974 14803 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/xm1/Collector
flabel locali 28850 14604 28968 14644 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/xm1/Base
flabel metal1 28800 14242 29040 14372 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/Emitter
flabel metal1 28450 14604 28690 14644 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/Base
flabel metal1 28286 14756 28526 14796 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/Collector
flabel metal1 28260 15082 28320 15142 1 FreeSans 1000 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/VPWR
flabel metal1 28260 13202 28320 13262 1 FreeSans 1000 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_3/VGND
flabel metal1 23696 14532 23816 14652 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_22/Rin
flabel metal1 23696 13572 23816 13692 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_22/Rout
flabel metal1 23576 15082 23636 15142 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_22/VPWR
flabel metal1 23576 13202 23636 13262 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_22/VGND
flabel metal1 39376 14532 39496 14652 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_16/Rin
flabel metal1 39376 13572 39496 13692 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_16/Rout
flabel metal1 39256 15082 39316 15142 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_16/VPWR
flabel metal1 39256 13202 39316 13262 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_16/VGND
flabel locali 10134 17296 10194 17356 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_9_0/GATE
flabel locali 10134 18682 10194 18742 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_9_0/SOURCE
flabel locali 10134 17462 10194 17522 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_9_0/DRAIN
flabel metal1 6014 18842 6074 18902 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_9_0/VPWR
flabel metal1 6014 16962 6074 17022 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_9_0/VGND
flabel metal1 10760 18292 10880 18412 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_5/Rin
flabel metal1 10760 17332 10880 17452 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_5/Rout
flabel metal1 10640 18842 10700 18902 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_5/VPWR
flabel metal1 10640 16962 10700 17022 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_5/VGND
flabel metal2 16108 18562 16308 18642 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_7/Cin
flabel metal4 16130 17132 16290 17232 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_7/Cout
flabel metal1 16110 18842 16170 18902 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_7/VPWR
flabel metal1 16110 16962 16170 17022 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_7/VGND
flabel metal1 13504 18292 13624 18412 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_6/Rin
flabel metal1 13504 17332 13624 17452 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_6/Rout
flabel metal1 13384 18842 13444 18902 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_6/VPWR
flabel metal1 13384 16962 13444 17022 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_6/VGND
flabel locali 26764 17096 26824 17156 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_6_0/GATE
flabel locali 26764 18682 26824 18722 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_6_0/SOURCE
flabel locali 26764 17202 26824 17262 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_6_0/DRAIN
flabel nwell 23850 18842 23910 18902 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_6_0/VPWR
flabel metal1 23850 16962 24008 17022 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_6_0/VGND
flabel locali 38194 17888 38442 17992 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Emitter
flabel locali 38253 18514 38354 18563 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Collector
flabel locali 38230 18364 38348 18404 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Base
flabel locali 36854 17888 37102 17992 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Emitter
flabel locali 36913 18514 37014 18563 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector
flabel locali 36890 18364 37008 18404 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Base
flabel locali 35514 17888 35762 17992 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Emitter
flabel locali 35573 18514 35674 18563 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector
flabel locali 35550 18364 35668 18404 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Base
flabel locali 34174 17888 34422 17992 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Emitter
flabel locali 34233 18514 34334 18563 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector
flabel locali 34210 18364 34328 18404 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Base
flabel locali 32834 17888 33082 17992 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Emitter
flabel locali 32893 18514 32994 18563 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector
flabel locali 32870 18364 32988 18404 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Base
flabel locali 31494 17888 31742 17992 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Emitter
flabel locali 31553 18514 31654 18563 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector
flabel locali 31530 18364 31648 18404 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Base
flabel locali 30154 17888 30402 17992 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter
flabel locali 30213 18514 30314 18563 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector
flabel locali 30190 18364 30308 18404 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Base
flabel locali 28814 17888 29062 17992 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/xm1/Emitter
flabel locali 28873 18514 28974 18563 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/xm1/Collector
flabel locali 28850 18364 28968 18404 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/xm1/Base
flabel metal1 28800 18002 29040 18132 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/Emitter
flabel metal1 28450 18364 28690 18404 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/Base
flabel metal1 28286 18516 28526 18556 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/Collector
flabel metal1 28260 18842 28320 18902 1 FreeSans 1000 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/VPWR
flabel metal1 28260 16962 28320 17022 1 FreeSans 1000 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_0/VGND
flabel metal1 39376 18292 39496 18412 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_17/Rin
flabel metal1 39376 17332 39496 17452 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_17/Rout
flabel metal1 39256 18842 39316 18902 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_17/VPWR
flabel metal1 39256 16962 39316 17022 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_17/VGND
flabel locali 13244 20856 13304 20916 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_12_0/GATE
flabel locali 13244 22442 13304 22482 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_12_0/SOURCE
flabel locali 13244 20962 13304 21022 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_12_0/DRAIN
flabel nwell 7582 22602 7642 22662 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_12_0/VPWR
flabel metal1 7582 20722 7740 20782 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_12_0/VGND
flabel metal2 13560 22322 13760 22402 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_5/Cin
flabel metal4 13582 20892 13742 20992 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_5/Cout
flabel metal1 13562 22602 13622 22662 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_5/VPWR
flabel metal1 13562 20722 13622 20782 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_5/VGND
flabel locali 21562 21648 21810 21752 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_1_0/xm1/Emitter
flabel locali 21621 22274 21722 22323 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_1_0/xm1/Collector
flabel locali 21598 22124 21716 22164 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_1_0/xm1/Base
flabel locali 21570 21762 21798 21892 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_1_0/Emitter
flabel locali 21782 22124 21902 22164 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_1_0/Base
flabel locali 21818 22276 21938 22316 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_1_0/Collector
flabel metal1 21008 22602 21068 22662 1 FreeSans 1000 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_1_0/VPWR
flabel metal1 21008 20722 21068 20782 1 FreeSans 1000 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_1_0/VGND
flabel locali 38194 21648 38442 21752 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Emitter
flabel locali 38253 22274 38354 22323 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Collector
flabel locali 38230 22124 38348 22164 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Base
flabel locali 36854 21648 37102 21752 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Emitter
flabel locali 36913 22274 37014 22323 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector
flabel locali 36890 22124 37008 22164 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Base
flabel locali 35514 21648 35762 21752 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Emitter
flabel locali 35573 22274 35674 22323 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector
flabel locali 35550 22124 35668 22164 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Base
flabel locali 34174 21648 34422 21752 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Emitter
flabel locali 34233 22274 34334 22323 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector
flabel locali 34210 22124 34328 22164 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Base
flabel locali 32834 21648 33082 21752 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Emitter
flabel locali 32893 22274 32994 22323 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector
flabel locali 32870 22124 32988 22164 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Base
flabel locali 31494 21648 31742 21752 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Emitter
flabel locali 31553 22274 31654 22323 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector
flabel locali 31530 22124 31648 22164 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Base
flabel locali 30154 21648 30402 21752 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter
flabel locali 30213 22274 30314 22323 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector
flabel locali 30190 22124 30308 22164 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Base
flabel locali 28814 21648 29062 21752 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/xm1/Emitter
flabel locali 28873 22274 28974 22323 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/xm1/Collector
flabel locali 28850 22124 28968 22164 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/xm1/Base
flabel metal1 28800 21762 29040 21892 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/Emitter
flabel metal1 28450 22124 28690 22164 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/Base
flabel metal1 28286 22276 28526 22316 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/Collector
flabel metal1 28260 22602 28320 22662 1 FreeSans 1000 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/VPWR
flabel metal1 28260 20722 28320 20782 1 FreeSans 1000 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_1/VGND
flabel locali 27088 21056 27148 21116 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_9_2/GATE
flabel locali 27088 22442 27148 22502 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_9_2/SOURCE
flabel locali 27088 21222 27148 21282 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_9_2/DRAIN
flabel metal1 22968 22602 23028 22662 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_9_2/VPWR
flabel metal1 22968 20722 23028 20782 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_9_2/VGND
flabel metal1 39866 22052 39986 22172 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_8/Rin
flabel metal1 39866 21092 39986 21212 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_8/Rout
flabel metal1 39746 22602 39806 22662 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_8/VPWR
flabel metal1 39746 20722 39806 20782 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_8/VGND
flabel metal1 6840 25812 6960 25932 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_7/Rin
flabel metal1 6840 24852 6960 24972 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_7/Rout
flabel metal1 6720 26362 6780 26422 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_7/VPWR
flabel metal1 6720 24482 6780 24542 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_7/VGND
flabel locali 15106 24616 15166 24676 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_12_1/GATE
flabel locali 15106 26202 15166 26242 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_12_1/SOURCE
flabel locali 15106 24722 15166 24782 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_12_1/DRAIN
flabel nwell 9444 26362 9504 26422 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_12_1/VPWR
flabel metal1 9444 24482 9602 24542 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_12_1/VGND
flabel metal2 15422 26082 15622 26162 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_9/Cin
flabel metal4 15444 24652 15604 24752 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_9/Cout
flabel metal1 15424 26362 15484 26422 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_9/VPWR
flabel metal1 15424 24482 15484 24542 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_9/VGND
flabel locali 38194 25408 38442 25512 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Emitter
flabel locali 38253 26034 38354 26083 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Collector
flabel locali 38230 25884 38348 25924 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Base
flabel locali 36854 25408 37102 25512 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Emitter
flabel locali 36913 26034 37014 26083 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector
flabel locali 36890 25884 37008 25924 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Base
flabel locali 35514 25408 35762 25512 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Emitter
flabel locali 35573 26034 35674 26083 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector
flabel locali 35550 25884 35668 25924 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Base
flabel locali 34174 25408 34422 25512 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Emitter
flabel locali 34233 26034 34334 26083 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector
flabel locali 34210 25884 34328 25924 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Base
flabel locali 32834 25408 33082 25512 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Emitter
flabel locali 32893 26034 32994 26083 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector
flabel locali 32870 25884 32988 25924 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Base
flabel locali 31494 25408 31742 25512 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Emitter
flabel locali 31553 26034 31654 26083 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector
flabel locali 31530 25884 31648 25924 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Base
flabel locali 30154 25408 30402 25512 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter
flabel locali 30213 26034 30314 26083 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector
flabel locali 30190 25884 30308 25924 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Base
flabel locali 28814 25408 29062 25512 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/xm1/Emitter
flabel locali 28873 26034 28974 26083 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/xm1/Collector
flabel locali 28850 25884 28968 25924 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/xm1/Base
flabel metal1 28800 25522 29040 25652 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/Emitter
flabel metal1 28450 25884 28690 25924 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/Base
flabel metal1 28286 26036 28526 26076 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/Collector
flabel metal1 28260 26362 28320 26422 1 FreeSans 1000 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/VPWR
flabel metal1 28260 24482 28320 24542 1 FreeSans 1000 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_8_2/VGND
flabel locali 27088 24816 27148 24876 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_9_1/GATE
flabel locali 27088 26202 27148 26262 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_9_1/SOURCE
flabel locali 27088 24982 27148 25042 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_9_1/DRAIN
flabel metal1 22968 26362 23028 26422 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_9_1/VPWR
flabel metal1 22968 24482 23028 24542 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_9_1/VGND
flabel metal1 39866 25812 39986 25932 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_0/Rin
flabel metal1 39866 24852 39986 24972 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_0/Rout
flabel metal1 39746 26362 39806 26422 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_0/VPWR
flabel metal1 39746 24482 39806 24542 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_0/VGND
flabel metal1 37514 29572 37634 29692 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_20/Rin
flabel metal1 37514 28612 37634 28732 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_20/Rout
flabel metal1 37394 30122 37454 30182 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_20/VPWR
flabel metal1 37394 28242 37454 28302 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_20/VGND
flabel metal1 40258 29572 40378 29692 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_18/Rin
flabel metal1 40258 28612 40378 28732 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_18/Rout
flabel metal1 40138 30122 40198 30182 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_18/VPWR
flabel metal1 40138 28242 40198 28302 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_18/VGND
flabel locali 36858 28376 36918 28436 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_6_1/GATE
flabel locali 36858 29962 36918 30002 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_6_1/SOURCE
flabel locali 36858 28482 36918 28542 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_6_1/DRAIN
flabel nwell 33944 30122 34004 30182 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_6_1/VPWR
flabel metal1 33944 28242 34102 28302 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_6_1/VGND
flabel locali 33562 28376 33622 28436 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_60_2/GATE
flabel locali 33562 29962 33622 30002 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_60_2/SOURCE
flabel locali 33562 28482 33622 28542 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_60_2/DRAIN
flabel nwell 5916 30122 5976 30182 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_60_2/VPWR
flabel metal1 5916 28242 6074 28302 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_60_2/VGND
flabel metal2 6602 33602 6802 33682 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_2/Cin
flabel metal4 6624 32172 6784 32272 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_2/Cout
flabel metal1 6604 33882 6664 33942 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_2/VPWR
flabel metal1 6604 32002 6664 32062 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_2/VGND
flabel locali 41696 32136 41756 32196 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_60_1/GATE
flabel locali 41696 33722 41756 33762 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_60_1/SOURCE
flabel locali 41696 32242 41756 32302 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_60_1/DRAIN
flabel nwell 14050 33882 14110 33942 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_60_1/VPWR
flabel metal1 14050 32002 14208 32062 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_60_1/VGND
flabel metal2 5916 37362 6116 37442 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_1/Cin
flabel metal4 5938 35932 6098 36032 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_1/Cout
flabel metal1 5918 37642 5978 37702 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_1/VPWR
flabel metal1 5918 35762 5978 35822 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_1/VGND
flabel metal2 13364 37362 13564 37442 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_3/Cin
flabel metal4 13386 35932 13546 36032 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_3/Cout
flabel metal1 13366 37642 13426 37702 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_3/VPWR
flabel metal1 13366 35762 13426 35822 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_3/VGND
flabel metal2 20812 37362 21012 37442 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_0/Cin
flabel metal4 20834 35932 20994 36032 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_0/Cout
flabel metal1 20814 37642 20874 37702 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_0/VPWR
flabel metal1 20814 35762 20874 35822 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_0/VGND
flabel locali 28784 35936 28844 35996 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_1_1/GATE
flabel locali 28784 37482 28844 37542 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_1_1/SOURCE
flabel locali 28784 36162 28844 36222 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_1_1/DRAIN
flabel metal1 28328 37642 28388 37702 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_1_1/VPWR
flabel metal1 28328 35762 28388 35822 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_1_1/VGND
flabel locali 38618 36688 38866 36792 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Emitter
flabel locali 38677 37314 38778 37363 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector
flabel locali 38654 37164 38772 37204 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Base
flabel locali 37278 36688 37526 36792 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Emitter
flabel locali 37337 37314 37438 37363 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector
flabel locali 37314 37164 37432 37204 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Base
flabel locali 35938 36688 36186 36792 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Emitter
flabel locali 35997 37314 36098 37363 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector
flabel locali 35974 37164 36092 37204 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Base
flabel locali 34598 36688 34846 36792 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Emitter
flabel locali 34657 37314 34758 37363 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector
flabel locali 34634 37164 34752 37204 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Base
flabel locali 33258 36688 33506 36792 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Emitter
flabel locali 33317 37314 33418 37363 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector
flabel locali 33294 37164 33412 37204 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Base
flabel locali 31918 36688 32166 36792 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Emitter
flabel locali 31977 37314 32078 37363 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector
flabel locali 31954 37164 32072 37204 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Base
flabel locali 30578 36688 30826 36792 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/xm1/Emitter
flabel locali 30637 37314 30738 37363 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/xm1/Collector
flabel locali 30614 37164 30732 37204 0 FreeSans 500 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/xm1/Base
flabel metal1 30564 36802 30804 36932 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/Emitter
flabel metal1 30214 37164 30454 37204 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/Base
flabel metal1 30050 37316 30290 37356 1 FreeSans 600 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/Collector
flabel metal1 30024 37642 30084 37702 1 FreeSans 1000 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/VPWR
flabel metal1 30024 35762 30084 35822 1 FreeSans 1000 0 0 0 sky130_asc_pnp_05v5_W3p40L3p40_7_0/VGND
flabel metal1 39866 37092 39986 37212 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_19/Rin
flabel metal1 39866 36132 39986 36252 1 FreeSans 600 0 0 0 sky130_asc_res_xhigh_po_2p85_1_19/Rout
flabel metal1 39746 37642 39806 37702 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_19/VPWR
flabel metal1 39746 35762 39806 35822 1 FreeSans 1000 0 0 0 sky130_asc_res_xhigh_po_2p85_1_19/VGND
flabel metal2 6798 41122 6998 41202 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_4/Cin
flabel metal4 6820 39692 6980 39792 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_4/Cout
flabel metal1 6800 41402 6860 41462 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_4/VPWR
flabel metal1 6800 39522 6860 39582 1 FreeSans 1000 0 0 0 sky130_asc_cap_mim_m3_1_4/VGND
flabel locali 6440 39696 6500 39756 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_1_0/GATE
flabel locali 6440 41242 6500 41302 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_1_0/SOURCE
flabel locali 6440 39922 6500 39982 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_1_0/DRAIN
flabel metal1 5984 41402 6044 41462 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_1_0/VPWR
flabel metal1 5984 39522 6044 39582 1 FreeSans 1000 0 0 0 sky130_asc_nfet_01v8_lvt_1_0/VGND
flabel locali 42578 39656 42638 39716 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_60_0/GATE
flabel locali 42578 41242 42638 41282 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_60_0/SOURCE
flabel locali 42578 39762 42638 39822 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_60_0/DRAIN
flabel nwell 14932 41402 14992 41462 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_60_0/VPWR
flabel metal1 14932 39522 15090 39582 1 FreeSans 1000 0 0 0 sky130_asc_pfet_01v8_lvt_60_0/VGND
<< end >>
