SIMPLE DIFFERENTIAL PAIR
VCC 7 0 12
VEE 8 0 -12
VIN 1 0 AC 1 DC 0
RS1 1 2 1K
RS2 6 0 1K
Q1 3 2 4 MOD1
Q2 5 6 4 MOD1
RC1 7 3 10K
RC2 7 5 10K
RE 4 8 10K
.MODEL MOD1 NPN BF=50 VAF=50 IS=1.E-12 RB=100 CJC=.5PF TF=.6NS
.ic v(1)=0 v(2)=-0.009996365874665257 v(3)=6.36449558290397 v(4)=-0.5290639756045419 v(5)=6.36449558290401
+ v(6)=-0.009996365874665384 v(7)=12.0 v(8)=-12.0 
.op
.save all
.TF V(2) VIN
* .control 
*     save all
*     tran 10ns 20us 0us
*     run
*     write ../raw-result/test_all.raw all
* .endc
.END