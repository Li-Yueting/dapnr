* NGSPICE file created from bgr_top_flat.ext - technology: sky130A

.subckt bgr_top_flat porst vbg VSS VDD
X0 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.t24 VDD.t439 VDD.t438 sky130_fd_pr__pfet_01v8_lvt ad=8.2639e+13p pd=5.2584e+08u as=0p ps=0u w=6.45e+06u l=2e+06u
X1 VSS.t94 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X2 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t8 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t62 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t14 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X3 VDD.t437 sky130_asc_pfet_01v8_lvt_60_0/GATE.t25 vbg.t59 VDD.t436 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X4 sky130_asc_pfet_01v8_lvt_60_0/GATE.t26 VDD.t143 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X5 sky130_asc_pfet_01v8_lvt_60_0/GATE.t27 VDD.t167 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X6 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t11 sky130_asc_pfet_01v8_lvt_60_0/GATE.t28 VDD.t435 VDD.t434 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X7 VDD.t433 sky130_asc_pfet_01v8_lvt_60_0/GATE.t29 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t60 VDD.t432 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X8 VDD.t431 sky130_asc_pfet_01v8_lvt_60_0/GATE.t30 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t10 VDD.t430 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X9 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t59 sky130_asc_pfet_01v8_lvt_60_0/GATE.t31 VDD.t429 VDD.t428 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X10 VSS.t95 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X11 sky130_asc_res_xhigh_po_2p85_1_21/Rout a_15392_9587.t0 VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X12 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.t32 VDD.t427 VDD.t426 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X13 sky130_asc_pfet_01v8_lvt_60_0/GATE.t33 VDD.t140 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X14 VSS VSS.t92 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X15 sky130_asc_pfet_01v8_lvt_60_0/GATE.t34 VDD.t349 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X16 VDD.t425 sky130_asc_pfet_01v8_lvt_60_0/GATE.t35 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t58 VDD.t424 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X17 VSS.t97 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X18 sky130_asc_pfet_01v8_lvt_60_0/GATE.t36 VDD.t348 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X19 VSS.t98 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X20 sky130_asc_res_xhigh_po_2p85_1_19/Rin.t0 a_39402_28387.t0 VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X21 VSS.t99 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X22 VDD.t423 sky130_asc_pfet_01v8_lvt_60_0/GATE.t37 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t9 VDD.t422 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X23 sky130_asc_pfet_01v8_lvt_60_0/GATE.t38 VDD.t142 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X24 VDD.t421 sky130_asc_pfet_01v8_lvt_60_0/GATE.t39 vbg.t58 VDD.t420 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X25 VSS VSS.t90 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X26 sky130_asc_pfet_01v8_lvt_60_0/GATE.t40 VDD.t343 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X27 sky130_asc_res_xhigh_po_2p85_1_17/Rout a_41264_17107.t0 VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X28 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.t41 VDD.t419 VDD.t418 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X29 sky130_asc_res_xhigh_po_2p85_1_14/Rin.t0 a_37148_9587.t1 VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X30 VSS VSS.t88 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X31 sky130_asc_res_xhigh_po_2p85_1_2/Rin.t0 a_9904_9587# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X32 VDD.t397 sky130_asc_pfet_01v8_lvt_60_0/GATE.t42 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t396 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X33 sky130_asc_pfet_01v8_lvt_60_0/GATE.t43 VDD.t107 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X34 sky130_asc_pfet_01v8_lvt_60_0/GATE.t44 VDD.t334 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X35 VDD.t417 sky130_asc_pfet_01v8_lvt_60_0/GATE.t45 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t8 VDD.t416 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X36 VSS.t102 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X37 sky130_asc_pfet_01v8_lvt_60_0/GATE.t46 VDD.t340 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X38 VDD.t413 sky130_asc_pfet_01v8_lvt_60_0/GATE.t47 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t7 VDD.t412 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X39 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t57 sky130_asc_pfet_01v8_lvt_60_0/GATE.t48 VDD.t415 VDD.t414 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X40 VSS.t103 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X41 VDD.t411 sky130_asc_pfet_01v8_lvt_60_0/GATE.t49 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t56 VDD.t410 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X42 sky130_asc_pfet_01v8_lvt_60_0/GATE.t50 VDD.t88 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X43 sky130_asc_pfet_01v8_lvt_60_0/GATE.t51 VDD.t325 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X44 sky130_asc_pfet_01v8_lvt_60_0/GATE.t33 VDD.t335 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X45 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t13 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t63 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t7 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X46 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t6 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t64 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t12 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X47 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t55 sky130_asc_pfet_01v8_lvt_60_0/GATE.t52 VDD.t409 VDD.t408 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X48 VDD.t407 sky130_asc_pfet_01v8_lvt_60_0/GATE.t53 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t54 VDD.t406 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X49 sky130_asc_res_xhigh_po_2p85_1_19/Rout a_41754_35907# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X50 sky130_asc_pfet_01v8_lvt_60_0/GATE.t54 VDD.t91 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X51 sky130_asc_res_xhigh_po_2p85_1_1/Rout a_9904_5827# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X52 VSS.t104 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X53 VSS.t105 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X54 sky130_asc_pfet_01v8_lvt_60_0/GATE.t55 VDD.t87 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X55 VSS.t106 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X56 VDD.t405 sky130_asc_pfet_01v8_lvt_60_0/GATE.t56 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t404 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X57 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.t57 VDD.t403 VDD.t402 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X58 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t11 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t65 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t5 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X59 VDD.t401 sky130_asc_pfet_01v8_lvt_60_0/GATE.t58 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t400 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X60 sky130_asc_pfet_01v8_lvt_60_0/GATE.t44 VDD.t98 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X61 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.t59 VDD.t399 VDD.t398 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X62 VSS.t107 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X63 VSS.t108 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X64 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t4 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t66 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t9 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X65 VSS.t109 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X66 VSS.t13 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t14 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t18 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X67 VSS.t110 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X68 sky130_asc_pfet_01v8_lvt_60_0/GATE.t43 VDD.t312 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X69 VSS VSS.t86 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X70 VSS.t112 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X71 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.t60 VDD.t395 VDD.t394 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X72 VDD.t393 sky130_asc_pfet_01v8_lvt_60_0/GATE.t61 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t53 VDD.t392 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X73 VSS.t113 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X74 VSS.t114 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X75 vbg.t57 sky130_asc_pfet_01v8_lvt_60_0/GATE.t62 VDD.t391 VDD.t390 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X76 VSS.t115 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X77 VSS.t116 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X78 sky130_asc_pfet_01v8_lvt_60_0/GATE.t26 VDD.t23 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X79 sky130_asc_res_xhigh_po_2p85_1_29/Rout.t0 a_30582_5827# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X80 VDD.t389 sky130_asc_pfet_01v8_lvt_60_0/GATE.t63 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t52 VDD.t388 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X81 VSS.t117 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X82 VSS.t118 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X83 sky130_asc_cap_mim_m3_1_3/Cout VDD.t20 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X84 VSS VSS.t84 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X85 VSS.t120 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X86 sky130_asc_res_xhigh_po_2p85_1_26/Rin a_27838_5827.t1 VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X87 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t6 sky130_asc_pfet_01v8_lvt_60_0/GATE.t64 VDD.t387 VDD.t386 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X88 vbg.t56 sky130_asc_pfet_01v8_lvt_60_0/GATE.t65 VDD.t385 VDD.t384 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X89 VSS.t121 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X90 sky130_asc_res_xhigh_po_2p85_1_24/Rin a_12648_9587# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X91 sky130_asc_res_xhigh_po_2p85_1_9/Rout a_15392_13347.t0 VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X92 vbg.t55 sky130_asc_pfet_01v8_lvt_60_0/GATE.t66 VDD.t383 VDD.t382 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X93 VSS.t122 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X94 sky130_asc_pfet_01v8_lvt_60_0/GATE.t54 VDD.t309 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X95 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.t67 VDD.t381 VDD.t380 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X96 sky130_asc_pfet_01v8_lvt_60_0/GATE.t55 VDD.t304 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X97 VDD.t379 sky130_asc_pfet_01v8_lvt_60_0/GATE.t68 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t378 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X98 VSS.t123 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X99 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.t69 VDD.t377 VDD.t376 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X100 VSS VSS.t82 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X101 VDD.t375 sky130_asc_pfet_01v8_lvt_60_0/GATE.t70 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t51 VDD.t374 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X102 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t50 sky130_asc_pfet_01v8_lvt_60_0/GATE.t71 VDD.t373 VDD.t372 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X103 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t10 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t67 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t3 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X104 sky130_asc_pfet_01v8_lvt_60_0/GATE.t72 VDD.t37 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X105 VSS.t125 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X106 sky130_asc_res_xhigh_po_2p85_1_3/Rin a_9904_9587# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X107 sky130_asc_res_xhigh_po_2p85_1_15/Rin a_39892_5827# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X108 sky130_asc_res_xhigh_po_2p85_1_13/Rin a_33326_5827# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X109 sky130_asc_pfet_01v8_lvt_60_0/GATE.t73 VDD.t9 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X110 VSS.t126 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X111 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t49 sky130_asc_pfet_01v8_lvt_60_0/GATE.t74 VDD.t371 VDD.t370 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X112 VSS VSS.t80 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X113 sky130_asc_pfet_01v8_lvt_60_0/GATE.t75 VDD.t8 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X114 sky130_asc_res_xhigh_po_2p85_1_12/Rout.t0 a_37148_5827# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X115 VSS.t128 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X116 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t61 a_39402_28387.t1 VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X117 VDD.t369 sky130_asc_pfet_01v8_lvt_60_0/GATE.t76 vbg.t54 VDD.t368 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X118 VSS.t129 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X119 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t48 sky130_asc_pfet_01v8_lvt_60_0/GATE.t77 VDD.t367 VDD.t366 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X120 sky130_asc_res_xhigh_po_2p85_1_9/Rin a_34404_9587# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X121 VDD.t365 sky130_asc_pfet_01v8_lvt_60_0/GATE.t78 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t364 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X122 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t47 sky130_asc_pfet_01v8_lvt_60_0/GATE.t79 VDD.t363 VDD.t362 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X123 VDD.t361 sky130_asc_pfet_01v8_lvt_60_0/GATE.t80 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t360 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X124 sky130_asc_res_xhigh_po_2p85_1_18/Rout a_42146_28387# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X125 VSS VSS.t78 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X126 sky130_asc_pfet_01v8_lvt_60_0/GATE.t81 VDD.t10 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X127 sky130_asc_res_xhigh_po_2p85_1_7/Rin a_8728_24627# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X128 VSS.t131 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X129 VSS.t132 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X130 VSS.t133 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X131 sky130_asc_res_xhigh_po_2p85_1_22/Rin.t0 a_25094_5827# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X132 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t46 sky130_asc_pfet_01v8_lvt_60_0/GATE.t82 VDD.t359 VDD.t358 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X133 VDD.t357 sky130_asc_pfet_01v8_lvt_60_0/GATE.t83 vbg.t53 VDD.t356 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X134 VSS.t134 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X135 VSS.t135 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X136 sky130_asc_res_xhigh_po_2p85_1_10/Rin a_34404_9587# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X137 sky130_asc_res_xhigh_po_2p85_1_24/Rin.t0 a_22350_5827.t0 VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X138 sky130_asc_pfet_01v8_lvt_60_0/GATE.t34 VDD.t349 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X139 VDD.t351 sky130_asc_pfet_01v8_lvt_60_0/GATE.t84 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t350 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X140 VSS.t10 a_41754_24627.t0 VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X141 VDD.t355 sky130_asc_pfet_01v8_lvt_60_0/GATE.t85 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t45 VDD.t354 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X142 VSS.t136 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X143 sky130_asc_pfet_01v8_lvt_60_0/GATE.t36 VDD.t348 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X144 VSS.t137 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X145 VSS VSS.t76 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X146 VSS.t139 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X147 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t44 sky130_asc_pfet_01v8_lvt_60_0/GATE.t86 VDD.t353 VDD.t352 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X148 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t5 sky130_asc_pfet_01v8_lvt_60_0/GATE.t87 VDD.t347 VDD.t346 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X149 VDD.t345 sky130_asc_pfet_01v8_lvt_60_0/GATE.t88 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t43 VDD.t344 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X150 sky130_asc_pfet_01v8_lvt_60_0/GATE.t40 VDD.t343 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X151 sky130_asc_pfet_01v8_lvt_60_0/GATE.t81 VDD.t15 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X152 VSS.t7 a_16849_5827# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=1.075e+07u
X153 sky130_asc_pfet_01v8_lvt_60_0/GATE.t73 VDD.t265 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X154 sky130_asc_pfet_01v8_lvt_60_0/GATE.t89 VDD.t264 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X155 sky130_asc_pfet_01v8_lvt_60_0/GATE.t75 VDD.t18 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X156 VDD.t342 sky130_asc_pfet_01v8_lvt_60_0/GATE.t90 vbg.t52 VDD.t341 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X157 VSS.t140 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X158 VSS VSS.t74 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X159 VSS.t142 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X160 sky130_asc_res_xhigh_po_2p85_1_30/Rout.t0 a_28916_9587.t1 VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X161 sky130_asc_pfet_01v8_lvt_60_0/GATE.t46 VDD.t340 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X162 VDD.t339 sky130_asc_pfet_01v8_lvt_60_0/GATE.t91 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t42 VDD.t338 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X163 sky130_asc_pfet_01v8_lvt_60_0/GATE.t92 VDD.t17 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X164 VSS VSS.t72 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X165 sky130_asc_res_xhigh_po_2p85_1_7/Rout.t0 a_15392_17107.t1 VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X166 sky130_asc_pfet_01v8_lvt_60_0/GATE.t93 VDD.t16 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X167 VSS VSS.t70 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X168 VDD.t337 sky130_asc_pfet_01v8_lvt_60_0/GATE.t94 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t41 VDD.t336 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X169 VDD.t49 sky130_asc_pfet_01v8_lvt_60_0/GATE.t95 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t48 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X170 sky130_asc_pfet_01v8_lvt_60_0/GATE.t33 VDD.t335 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X171 sky130_asc_res_xhigh_po_2p85_1_16/Rout.t0 a_41264_13347# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X172 sky130_asc_pfet_01v8_lvt_60_0/GATE.t44 VDD.t334 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X173 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.t96 VDD.t333 VDD.t332 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X174 VSS VSS.t68 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X175 sky130_asc_res_xhigh_po_2p85_1_24/Rout.t0 a_12648_9587# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X176 sky130_asc_pfet_01v8_lvt_60_0/GATE.t97 VDD.t13 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X177 VDD.t331 sky130_asc_pfet_01v8_lvt_60_0/GATE.t98 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t40 VDD.t330 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X178 VSS.t4 a_26159_9587# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=1.075e+07u
X179 VSS.t146 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X180 sky130_asc_pfet_01v8_lvt_60_0/GATE.t40 VDD.t229 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X181 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t39 sky130_asc_pfet_01v8_lvt_60_0/GATE.t99 VDD.t329 VDD.t328 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X182 sky130_asc_pfet_01v8_lvt_60_0/GATE.t51 VDD.t325 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X183 VSS VSS.t66 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X184 VSS.t148 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X185 sky130_asc_res_xhigh_po_2p85_1_9/Rin a_15392_13347.t1 VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X186 vbg.t51 sky130_asc_pfet_01v8_lvt_60_0/GATE.t100 VDD.t327 VDD.t326 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X187 VDD.t324 sky130_asc_pfet_01v8_lvt_60_0/GATE.t101 vbg.t50 VDD.t323 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X188 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t8 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.t17 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X189 VSS.t149 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X190 sky130_asc_pfet_01v8_lvt_60_0/GATE.t43 VDD.t312 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X191 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t38 sky130_asc_pfet_01v8_lvt_60_0/GATE.t102 VDD.t322 VDD.t321 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X192 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.t103 VDD.t318 VDD.t317 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X193 VSS.t150 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X194 sky130_asc_res_xhigh_po_2p85_1_5/Rout.t0 a_12648_17107.t0 VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X195 VSS.t151 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X196 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t37 sky130_asc_pfet_01v8_lvt_60_0/GATE.t104 VDD.t320 VDD.t319 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X197 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t36 sky130_asc_pfet_01v8_lvt_60_0/GATE.t105 VDD.t316 VDD.t315 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X198 sky130_asc_pfet_01v8_lvt_60_0/GATE.t106 VDD.t144 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X199 VSS.t152 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X200 VDD.t314 sky130_asc_pfet_01v8_lvt_60_0/GATE.t107 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t313 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X201 sky130_asc_pfet_01v8_lvt_60_0/GATE.t26 VDD.t23 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X202 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t35 sky130_asc_pfet_01v8_lvt_60_0/GATE.t108 VDD.t311 VDD.t310 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X203 sky130_asc_pfet_01v8_lvt_60_0/GATE.t38 VDD.t22 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X204 sky130_asc_pfet_01v8_lvt_60_0/GATE.t93 VDD.t21 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X205 sky130_asc_res_xhigh_po_2p85_1_12/Rin.t0 a_39892_9587.t1 VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X206 VSS.t153 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X207 sky130_asc_cap_mim_m3_1_3/Cout VDD.t20 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X208 sky130_asc_pfet_01v8_lvt_60_0/GATE.t109 VDD.t202 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X209 VSS.t154 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X210 sky130_asc_pfet_01v8_lvt_60_0/GATE.t54 VDD.t309 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X211 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t0 a_42146_28387# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X212 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t34 sky130_asc_pfet_01v8_lvt_60_0/GATE.t110 VDD.t308 VDD.t307 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X213 VSS.t155 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X214 VSS.t156 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X215 sky130_asc_pfet_01v8_lvt_60_0/GATE.t55 VDD.t304 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X216 VSS.t157 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X217 VSS VSS.t64 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X218 VDD.t306 sky130_asc_pfet_01v8_lvt_60_0/GATE.t111 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t33 VDD.t305 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X219 VDD.t303 sky130_asc_pfet_01v8_lvt_60_0/GATE.t112 vbg.t49 VDD.t302 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X220 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t32 sky130_asc_pfet_01v8_lvt_60_0/GATE.t113 VDD.t301 VDD.t300 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X221 VSS.t159 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X222 VSS.t160 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X223 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t31 sky130_asc_pfet_01v8_lvt_60_0/GATE.t114 VDD.t299 VDD.t298 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X224 VSS.t161 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X225 VDD.t297 sky130_asc_pfet_01v8_lvt_60_0/GATE.t115 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t296 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X226 VSS VSS.t62 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X227 VDD.t295 sky130_asc_pfet_01v8_lvt_60_0/GATE.t116 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t30 VDD.t294 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X228 sky130_asc_res_xhigh_po_2p85_1_29/Rout a_28916_9587.t0 VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X229 VSS.t163 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X230 VSS.t164 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X231 sky130_asc_res_xhigh_po_2p85_1_18/Rout.t0 a_41264_17107.t1 VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X232 VSS VSS.t60 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X233 VSS VSS.t58 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X234 VSS.t167 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X235 VDD.t293 sky130_asc_pfet_01v8_lvt_60_0/GATE.t117 vbg.t48 VDD.t292 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X236 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t29 sky130_asc_pfet_01v8_lvt_60_0/GATE.t118 VDD.t291 VDD.t290 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X237 vbg.t47 sky130_asc_pfet_01v8_lvt_60_0/GATE.t119 VDD.t289 VDD.t288 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X238 VSS.t168 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X239 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t20 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t19 VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X240 VSS VSS.t56 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X241 sky130_asc_res_xhigh_po_2p85_1_26/Rin.t0 a_19606_5827# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X242 VDD.t493 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t17 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t18 VDD.t492 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X243 VDD.t285 sky130_asc_pfet_01v8_lvt_60_0/GATE.t120 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t28 VDD.t284 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X244 VSS.t170 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X245 VSS.t171 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X246 VDD.t287 sky130_asc_pfet_01v8_lvt_60_0/GATE.t121 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t27 VDD.t286 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X247 VSS VSS.t54 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X248 VDD.t283 sky130_asc_pfet_01v8_lvt_60_0/GATE.t122 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t282 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X249 VDD.t25 sky130_asc_pfet_01v8_lvt_60_0/GATE.t123 vbg.t46 VDD.t24 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X250 VSS.t173 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X251 VSS.t174 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X252 sky130_asc_cap_mim_m3_1_3/Cout VDD.t141 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X253 VDD.t279 sky130_asc_pfet_01v8_lvt_60_0/GATE.t124 vbg.t45 VDD.t278 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X254 VDD.t281 sky130_asc_pfet_01v8_lvt_60_0/GATE.t125 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t26 VDD.t280 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X255 sky130_asc_pfet_01v8_lvt_60_0/GATE.t27 VDD.t125 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X256 VDD.t277 sky130_asc_pfet_01v8_lvt_60_0/GATE.t126 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t25 VDD.t276 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X257 VSS.t175 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X258 sky130_asc_pfet_01v8_lvt_60_0/GATE.t109 VDD.t124 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X259 VDD.t275 sky130_asc_pfet_01v8_lvt_60_0/GATE.t127 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t274 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X260 VDD.t273 sky130_asc_pfet_01v8_lvt_60_0/GATE.t128 vbg.t44 VDD.t272 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X261 VSS VSS.t52 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X262 sky130_asc_res_xhigh_po_2p85_1_17/Rout.t0 a_41264_13347# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X263 sky130_asc_res_xhigh_po_2p85_1_19/Rin a_41754_35907# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X264 VDD.t271 sky130_asc_pfet_01v8_lvt_60_0/GATE.t129 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t24 VDD.t270 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X265 VSS.t177 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X266 sky130_asc_pfet_01v8_lvt_60_0/GATE.t130 VDD.t19 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X267 sky130_asc_res_xhigh_po_2p85_1_2/Rout.t0 a_9904_5827# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X268 VDD.t269 sky130_asc_pfet_01v8_lvt_60_0/GATE.t131 vbg.t43 VDD.t268 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X269 VSS.t178 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X270 VSS.t179 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X271 VSS VSS.t50 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X272 vbg.t42 sky130_asc_pfet_01v8_lvt_60_0/GATE.t132 VDD.t267 VDD.t266 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X273 sky130_asc_pfet_01v8_lvt_60_0/GATE.t73 VDD.t265 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X274 VSS.t181 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X275 VSS VSS.t48 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X276 sky130_asc_pfet_01v8_lvt_60_0/GATE.t89 VDD.t264 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X277 vbg.t41 sky130_asc_pfet_01v8_lvt_60_0/GATE.t133 VDD.t263 VDD.t262 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X278 sky130_asc_pfet_01v8_lvt_60_0/GATE.t75 VDD.t18 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X279 VDD.t261 sky130_asc_pfet_01v8_lvt_60_0/GATE.t134 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t23 VDD.t260 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X280 VDD.t259 sky130_asc_pfet_01v8_lvt_60_0/GATE.t135 vbg.t40 VDD.t258 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X281 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t22 sky130_asc_pfet_01v8_lvt_60_0/GATE.t136 VDD.t257 VDD.t256 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X282 VSS.t183 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X283 sky130_asc_pfet_01v8_lvt_60_0/GATE.t92 VDD.t17 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X284 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.t137 VDD.t47 VDD.t46 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X285 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t21 sky130_asc_pfet_01v8_lvt_60_0/GATE.t138 VDD.t255 VDD.t254 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X286 vbg.t39 sky130_asc_pfet_01v8_lvt_60_0/GATE.t139 VDD.t253 VDD.t252 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X287 VDD.t251 sky130_asc_pfet_01v8_lvt_60_0/GATE.t140 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t20 VDD.t250 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X288 VSS.t184 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X289 sky130_asc_res_xhigh_po_2p85_1_7/Rin a_41754_20867# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X290 sky130_asc_pfet_01v8_lvt_60_0/GATE.t93 VDD.t16 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X291 sky130_asc_pfet_01v8_lvt_60_0/GATE.t81 VDD.t15 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X292 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.t141 VDD.t249 VDD.t248 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X293 vbg.t38 sky130_asc_pfet_01v8_lvt_60_0/GATE.t142 VDD.t247 VDD.t246 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X294 sky130_asc_pfet_01v8_lvt_60_0/GATE.t34 VDD.t14 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X295 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t19 sky130_asc_pfet_01v8_lvt_60_0/GATE.t143 VDD.t245 VDD.t244 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X296 VSS.t185 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X297 sky130_asc_res_xhigh_po_2p85_1_30/Rout a_31660_9587.t0 VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X298 VDD.t29 sky130_asc_pfet_01v8_lvt_60_0/GATE.t144 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t18 VDD.t28 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X299 VSS VSS.t46 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X300 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t17 sky130_asc_pfet_01v8_lvt_60_0/GATE.t145 VDD.t243 VDD.t242 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X301 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.t146 VDD.t241 VDD.t240 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X302 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.t147 VDD.t239 VDD.t238 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X303 vbg.t37 sky130_asc_pfet_01v8_lvt_60_0/GATE.t148 VDD.t237 VDD.t236 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X304 VDD.t235 sky130_asc_pfet_01v8_lvt_60_0/GATE.t149 vbg.t36 VDD.t234 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X305 VSS VSS.t44 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X306 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t7 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.t9 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X307 sky130_asc_pfet_01v8_lvt_60_0/GATE.t97 VDD.t13 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X308 sky130_asc_pfet_01v8_lvt_60_0/GATE.t12 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t6 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X309 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t16 sky130_asc_pfet_01v8_lvt_60_0/GATE.t150 VDD.t27 VDD.t26 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X310 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.t151 VDD.t45 VDD.t44 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X311 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t15 sky130_asc_pfet_01v8_lvt_60_0/GATE.t152 VDD.t53 VDD.t52 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X312 VDD.t233 sky130_asc_pfet_01v8_lvt_60_0/GATE.t153 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t232 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X313 VSS VSS.t42 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X314 sky130_asc_pfet_01v8_lvt_60_0/GATE.t40 VDD.t229 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X315 VDD.t231 sky130_asc_pfet_01v8_lvt_60_0/GATE.t154 vbg.t35 VDD.t230 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X316 sky130_asc_pfet_01v8_lvt_60_0/GATE.t155 VDD.t58 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X317 sky130_asc_pfet_01v8_lvt_60_0/GATE.t23 porst.t0 VSS.t12 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X318 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.t156 VDD.t228 VDD.t227 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X319 VDD.t3 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t15 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t16 VDD.t2 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X320 sky130_asc_pfet_01v8_lvt_60_0/GATE.t89 VDD.t12 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X321 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t14 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t13 VDD.t487 VDD.t486 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X322 VSS.t189 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X323 VSS.t190 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X324 sky130_asc_pfet_01v8_lvt_60_0/GATE.t157 VDD.t11 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X325 VDD.t226 sky130_asc_pfet_01v8_lvt_60_0/GATE.t158 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t225 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X326 vbg.t34 sky130_asc_pfet_01v8_lvt_60_0/GATE.t159 VDD.t224 VDD.t223 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X327 VDD.t222 sky130_asc_pfet_01v8_lvt_60_0/GATE.t160 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t14 VDD.t221 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X328 VDD.t489 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t21 sky130_asc_pfet_01v8_lvt_60_0/GATE.t20 VDD.t488 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X329 VSS.t191 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X330 VDD.t220 sky130_asc_pfet_01v8_lvt_60_0/GATE.t161 vbg.t33 VDD.t219 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X331 sky130_asc_pfet_01v8_lvt_60_0/GATE.t50 VDD.t72 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X332 sky130_asc_pfet_01v8_lvt_60_0/GATE.t21 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t22 VDD.t491 VDD.t490 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X333 sky130_asc_pfet_01v8_lvt_60_0/GATE.t162 VDD.t63 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X334 VDD.t146 sky130_asc_pfet_01v8_lvt_60_0/GATE.t163 vbg.t32 VDD.t145 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X335 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.t164 VDD.t208 VDD.t207 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X336 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t13 sky130_asc_pfet_01v8_lvt_60_0/GATE.t165 VDD.t210 VDD.t209 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X337 VDD.t218 sky130_asc_pfet_01v8_lvt_60_0/GATE.t166 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t12 VDD.t217 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X338 sky130_asc_pfet_01v8_lvt_60_0/GATE.t162 VDD.t56 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X339 VDD.t216 sky130_asc_pfet_01v8_lvt_60_0/GATE.t167 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t215 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X340 VDD.t214 sky130_asc_pfet_01v8_lvt_60_0/GATE.t168 vbg.t31 VDD.t213 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X341 sky130_asc_pfet_01v8_lvt_60_0/GATE.t22 porst.t1 VSS.t11 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X342 VSS.t192 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X343 sky130_asc_pfet_01v8_lvt_60_0/GATE.t106 VDD.t144 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X344 VSS VSS.t40 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X345 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t11 sky130_asc_pfet_01v8_lvt_60_0/GATE.t169 VDD.t212 VDD.t211 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X346 VDD.t206 sky130_asc_pfet_01v8_lvt_60_0/GATE.t170 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t10 VDD.t205 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X347 VDD.t204 sky130_asc_pfet_01v8_lvt_60_0/GATE.t171 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t203 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X348 sky130_asc_pfet_01v8_lvt_60_0/GATE.t93 VDD.t21 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X349 VDD.t156 sky130_asc_pfet_01v8_lvt_60_0/GATE.t172 vbg.t30 VDD.t155 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X350 sky130_asc_pfet_01v8_lvt_60_0/GATE.t109 VDD.t202 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X351 VSS VSS.t38 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X352 sky130_asc_res_xhigh_po_2p85_1_22/Rout.t0 a_15392_9587.t1 VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X353 VSS.t1 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t12 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t13 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X354 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t479 VDD.t481 VDD.t480 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X355 sky130_asc_pfet_01v8_lvt_60_0/GATE.t15 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t5 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X356 VDD.t201 sky130_asc_pfet_01v8_lvt_60_0/GATE.t173 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t200 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X357 VDD.t478 VDD.t476 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t477 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X358 VDD.t199 sky130_asc_pfet_01v8_lvt_60_0/GATE.t174 vbg.t29 VDD.t198 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X359 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t9 sky130_asc_pfet_01v8_lvt_60_0/GATE.t175 VDD.t150 VDD.t149 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X360 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t15 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t68 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t2 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X361 vbg.t28 sky130_asc_pfet_01v8_lvt_60_0/GATE.t176 VDD.t154 VDD.t153 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X362 VDD.t191 sky130_asc_pfet_01v8_lvt_60_0/GATE.t177 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t190 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X363 VDD.t197 sky130_asc_pfet_01v8_lvt_60_0/GATE.t178 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t8 VDD.t196 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X364 sky130_asc_res_xhigh_po_2p85_1_23/Rin a_25094_5827# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X365 sky130_asc_pfet_01v8_lvt_60_0/GATE.t97 VDD.t57 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X366 VSS.t195 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X367 sky130_asc_res_xhigh_po_2p85_1_2/Rout a_12648_13347# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X368 VDD.t195 sky130_asc_pfet_01v8_lvt_60_0/GATE.t179 vbg.t27 VDD.t194 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X369 vbg.t26 sky130_asc_pfet_01v8_lvt_60_0/GATE.t180 VDD.t193 VDD.t192 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X370 sky130_asc_res_xhigh_po_2p85_1_26/Rout.t0 a_22350_5827.t1 VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X371 VSS.t196 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X372 sky130_asc_pfet_01v8_lvt_60_0/GATE.t181 VDD.t36 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X373 VSS.t8 porst.t2 sky130_asc_pfet_01v8_lvt_60_0/GATE.t5 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X374 VSS VSS.t36 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X375 sky130_asc_pfet_01v8_lvt_60_0/GATE.t38 VDD.t22 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X376 sky130_asc_res_xhigh_po_2p85_1_0/Rin.t0 a_41754_24627.t1 VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X377 VDD.t1 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t11 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t12 VDD.t0 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X378 VDD.t148 sky130_asc_pfet_01v8_lvt_60_0/GATE.t182 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t7 VDD.t147 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X379 VDD.t189 sky130_asc_pfet_01v8_lvt_60_0/GATE.t183 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t188 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X380 VDD.t187 sky130_asc_pfet_01v8_lvt_60_0/GATE.t184 vbg.t25 VDD.t186 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X381 sky130_asc_res_xhigh_po_2p85_1_4/Rout.t0 a_9904_13347# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X382 sky130_asc_res_xhigh_po_2p85_1_12/Rout a_39892_9587.t0 VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X383 vbg.t24 sky130_asc_pfet_01v8_lvt_60_0/GATE.t185 VDD.t185 VDD.t184 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X384 VSS.t198 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X385 VDD.t441 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t23 sky130_asc_pfet_01v8_lvt_60_0/GATE.t6 VDD.t440 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X386 VSS VSS.t34 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X387 vbg.t23 sky130_asc_pfet_01v8_lvt_60_0/GATE.t186 VDD.t183 VDD.t182 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X388 VSS.t200 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X389 sky130_asc_res_xhigh_po_2p85_1_21/Rout.t0 a_16849_5827# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=1.075e+07u
X390 VDD.t181 sky130_asc_pfet_01v8_lvt_60_0/GATE.t187 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t6 VDD.t180 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X391 VDD.t179 sky130_asc_pfet_01v8_lvt_60_0/GATE.t188 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t178 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X392 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t5 sky130_asc_pfet_01v8_lvt_60_0/GATE.t189 VDD.t177 VDD.t176 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X393 sky130_asc_pfet_01v8_lvt_60_0/GATE.t26 VDD.t143 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X394 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.t190 VDD.t175 VDD.t174 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X395 VSS.t201 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X396 sky130_asc_res_xhigh_po_2p85_1_14/Rout.t0 a_37148_9587.t0 VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X397 vbg.t22 sky130_asc_pfet_01v8_lvt_60_0/GATE.t191 VDD.t152 VDD.t151 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X398 sky130_asc_pfet_01v8_lvt_60_0/GATE.t27 VDD.t167 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X399 sky130_asc_res_xhigh_po_2p85_1_28/Rout a_30582_5827# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X400 sky130_asc_res_xhigh_po_2p85_1_22/Rout a_25584_13347# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X401 VSS VSS.t32 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X402 vbg.t21 sky130_asc_pfet_01v8_lvt_60_0/GATE.t192 VDD.t171 VDD.t170 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X403 VDD.t173 sky130_asc_pfet_01v8_lvt_60_0/GATE.t193 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t172 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X404 VSS.t203 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X405 sky130_asc_pfet_01v8_lvt_60_0/GATE.t7 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t24 VDD.t443 VDD.t442 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X406 VSS.t9 porst.t3 sky130_asc_pfet_01v8_lvt_60_0/GATE.t8 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X407 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.t194 VDD.t169 VDD.t168 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X408 vbg.t20 sky130_asc_pfet_01v8_lvt_60_0/GATE.t195 VDD.t166 VDD.t165 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X409 VDD.t475 VDD.t473 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t474 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X410 sky130_asc_res_xhigh_po_2p85_1_26/Rout a_27838_5827.t0 VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X411 sky130_asc_pfet_01v8_lvt_60_0/GATE.t38 VDD.t142 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X412 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t470 VDD.t472 VDD.t471 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X413 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t467 VDD.t469 VDD.t468 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X414 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.t196 VDD.t164 VDD.t163 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X415 VSS VSS.t14 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__pnp_05v5_W3p40L3p40
X416 vbg.t19 sky130_asc_pfet_01v8_lvt_60_0/GATE.t197 VDD.t162 VDD.t161 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X417 VDD.t160 sky130_asc_pfet_01v8_lvt_60_0/GATE.t198 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t4 VDD.t159 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X418 VSS.t205 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X419 VSS.t206 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X420 sky130_asc_cap_mim_m3_1_3/Cout VDD.t141 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X421 sky130_asc_pfet_01v8_lvt_60_0/GATE.t33 VDD.t140 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X422 vbg.t18 sky130_asc_pfet_01v8_lvt_60_0/GATE.t199 VDD.t158 VDD.t157 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X423 VSS.t207 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X424 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t3 sky130_asc_pfet_01v8_lvt_60_0/GATE.t200 VDD.t139 VDD.t138 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X425 vbg.t60 a_41754_20867# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X426 VSS VSS.t30 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X427 vbg.t17 sky130_asc_pfet_01v8_lvt_60_0/GATE.t201 VDD.t137 VDD.t136 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X428 sky130_asc_pfet_01v8_lvt_60_0/GATE.t27 VDD.t125 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X429 sky130_asc_pfet_01v8_lvt_60_0/GATE.t109 VDD.t124 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X430 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t4 sky130_asc_pfet_01v8_lvt_60_0/GATE.t202 VDD.t135 VDD.t134 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X431 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.t203 VDD.t133 VDD.t132 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X432 VSS VSS.t28 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X433 vbg.t16 sky130_asc_pfet_01v8_lvt_60_0/GATE.t204 VDD.t127 VDD.t126 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X434 sky130_asc_pfet_01v8_lvt_60_2/DRAIN a_31660_9587.t1 VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X435 VDD.t129 sky130_asc_pfet_01v8_lvt_60_0/GATE.t205 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t2 VDD.t128 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X436 sky130_asc_res_xhigh_po_2p85_1_15/Rout a_39892_5827# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X437 VSS.t0 porst.t4 sky130_asc_pfet_01v8_lvt_60_0/GATE.t0 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X438 VDD.t131 sky130_asc_pfet_01v8_lvt_60_0/GATE.t206 vbg.t15 VDD.t130 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X439 VSS.t210 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X440 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.t207 VDD.t123 VDD.t122 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X441 sky130_asc_res_xhigh_po_2p85_1_13/Rout a_33326_5827# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X442 VDD.t466 VDD.t464 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t465 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X443 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t461 VDD.t463 VDD.t462 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X444 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.t208 VDD.t121 VDD.t120 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X445 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t1 sky130_asc_pfet_01v8_lvt_60_0/GATE.t209 VDD.t119 VDD.t118 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X446 vbg.t14 sky130_asc_pfet_01v8_lvt_60_0/GATE.t210 VDD.t117 VDD.t116 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X447 sky130_asc_pfet_01v8_lvt_60_0/GATE.t130 VDD.t19 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X448 VDD.t115 sky130_asc_pfet_01v8_lvt_60_0/GATE.t211 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t114 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X449 sky130_asc_res_xhigh_po_2p85_1_10/Rin.t0 a_37148_5827# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X450 VSS VSS.t26 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X451 VSS.t212 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X452 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t4 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.t11 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X453 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t458 VDD.t460 VDD.t459 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X454 sky130_asc_pfet_01v8_lvt_60_0/GATE.t13 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t3 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X455 VDD.t113 sky130_asc_pfet_01v8_lvt_60_0/GATE.t212 vbg.t13 VDD.t112 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X456 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.t213 VDD.t111 VDD.t110 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X457 sky130_asc_pfet_01v8_lvt_60_0/GATE.t43 VDD.t107 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X458 VSS.t213 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X459 vbg.t12 sky130_asc_pfet_01v8_lvt_60_0/GATE.t214 VDD.t109 VDD.t108 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X460 sky130_asc_res_xhigh_po_2p85_1_7/Rout a_8728_24627# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X461 VDD.t106 sky130_asc_pfet_01v8_lvt_60_0/GATE.t215 vbg.t11 VDD.t105 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X462 VSS.t214 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X463 sky130_asc_pfet_01v8_lvt_60_0/GATE.t2 porst.t5 VSS.t3 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X464 VSS.t215 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X465 VSS.t216 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X466 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t2 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.t10 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X467 sky130_asc_pfet_01v8_lvt_60_0/GATE.t14 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X468 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.t216 VDD.t104 VDD.t103 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X469 sky130_asc_res_xhigh_po_2p85_1_6/Rout.t0 a_12648_17107.t1 VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X470 VDD.t102 sky130_asc_pfet_01v8_lvt_60_0/GATE.t217 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t101 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X471 VDD.t100 sky130_asc_pfet_01v8_lvt_60_0/GATE.t218 vbg.t10 VDD.t99 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X472 sky130_asc_pfet_01v8_lvt_60_0/GATE.t50 VDD.t88 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X473 sky130_asc_pfet_01v8_lvt_60_0/GATE.t34 VDD.t14 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X474 sky130_asc_pfet_01v8_lvt_60_0/GATE.t44 VDD.t98 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X475 VSS.t217 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X476 VDD.t97 sky130_asc_pfet_01v8_lvt_60_0/GATE.t219 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t3 VDD.t96 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X477 VDD.t95 sky130_asc_pfet_01v8_lvt_60_0/GATE.t220 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t94 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X478 VDD.t93 sky130_asc_pfet_01v8_lvt_60_0/GATE.t221 vbg.t9 VDD.t92 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X479 VSS.t6 porst.t6 sky130_asc_pfet_01v8_lvt_60_0/GATE.t4 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X480 sky130_asc_pfet_01v8_lvt_60_0/GATE.t3 porst.t7 VSS.t5 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X481 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t10 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t9 VDD.t445 VDD.t444 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X482 sky130_asc_pfet_01v8_lvt_60_0/GATE.t54 VDD.t91 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X483 VDD.t90 sky130_asc_pfet_01v8_lvt_60_0/GATE.t222 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t89 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X484 sky130_asc_pfet_01v8_lvt_60_0/GATE.t55 VDD.t87 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X485 VDD.t483 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t25 sky130_asc_pfet_01v8_lvt_60_0/GATE.t18 VDD.t482 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X486 VDD.t86 sky130_asc_pfet_01v8_lvt_60_0/GATE.t223 vbg.t8 VDD.t85 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X487 VSS.t218 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X488 sky130_asc_pfet_01v8_lvt_60_0/GATE.t19 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t26 VDD.t485 VDD.t484 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X489 VSS VSS.t24 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X490 VDD.t84 sky130_asc_pfet_01v8_lvt_60_0/GATE.t224 vbg.t7 VDD.t83 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X491 VSS.t220 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X492 VDD.t457 VDD.t455 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t456 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X493 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.t225 VDD.t82 VDD.t81 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X494 VDD.t80 sky130_asc_pfet_01v8_lvt_60_0/GATE.t226 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t2 VDD.t79 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X495 vbg.t6 sky130_asc_pfet_01v8_lvt_60_0/GATE.t227 VDD.t78 VDD.t77 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X496 VDD.t76 sky130_asc_pfet_01v8_lvt_60_0/GATE.t228 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t75 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X497 sky130_asc_pfet_01v8_lvt_60_0/GATE.t89 VDD.t12 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X498 sky130_asc_res_xhigh_po_2p85_1_6/Rout a_15392_17107.t0 VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X499 sky130_asc_pfet_01v8_lvt_60_0/GATE.t157 VDD.t11 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X500 sky130_asc_res_xhigh_po_2p85_1_2/Rin a_12648_13347# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X501 vbg.t5 sky130_asc_pfet_01v8_lvt_60_0/GATE.t229 VDD.t74 VDD.t73 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X502 VSS.t221 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X503 sky130_asc_pfet_01v8_lvt_60_0/GATE.t50 VDD.t72 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X504 VDD.t454 VDD.t452 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t453 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X505 VDD.t71 sky130_asc_pfet_01v8_lvt_60_0/GATE.t230 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t70 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X506 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t449 VDD.t451 VDD.t450 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X507 VSS VSS.t22 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X508 VDD.t448 VDD.t446 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t447 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X509 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t16 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t69 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X510 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t0 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.t16 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X511 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.t231 VDD.t43 VDD.t42 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X512 vbg.t4 sky130_asc_pfet_01v8_lvt_60_0/GATE.t232 VDD.t51 VDD.t50 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X513 sky130_asc_res_xhigh_po_2p85_1_4/Rin a_9904_13347# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X514 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t0 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t70 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t17 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X515 sky130_asc_pfet_01v8_lvt_60_0/GATE.t155 VDD.t58 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X516 sky130_asc_res_xhigh_po_2p85_1_28/Rout a_19606_5827# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X517 VDD.t69 sky130_asc_pfet_01v8_lvt_60_0/GATE.t233 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t68 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X518 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t1 sky130_asc_pfet_01v8_lvt_60_0/GATE.t234 VDD.t60 VDD.t59 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X519 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.t235 VDD.t65 VDD.t64 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X520 VSS.t223 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X521 vbg.t3 sky130_asc_pfet_01v8_lvt_60_0/GATE.t236 VDD.t67 VDD.t66 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X522 VSS.t224 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X523 sky130_asc_res_xhigh_po_2p85_1_9/Rout.t0 a_26159_9587# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=1.075e+07u
X524 sky130_asc_res_xhigh_po_2p85_1_22/Rin a_25584_13347# VSS sky130_fd_pr__res_xhigh_po w=2.85e+06u l=7.88e+06u
X525 VSS.t225 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X526 sky130_asc_pfet_01v8_lvt_60_0/GATE.t162 VDD.t63 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X527 VSS.t226 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X528 vbg.t2 sky130_asc_pfet_01v8_lvt_60_0/GATE.t237 VDD.t62 VDD.t61 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X529 sky130_asc_pfet_01v8_lvt_60_0/GATE.t97 VDD.t57 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X530 sky130_asc_pfet_01v8_lvt_60_0/GATE.t162 VDD.t56 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X531 VSS VSS.t20 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X532 VSS.t228 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X533 VDD.t55 sky130_asc_pfet_01v8_lvt_60_0/GATE.t238 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t54 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X534 VDD.t41 sky130_asc_pfet_01v8_lvt_60_0/GATE.t239 vbg.t1 VDD.t40 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X535 VSS.t229 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X536 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.t240 VDD.t39 VDD.t38 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X537 VSS VSS.t18 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
X538 sky130_asc_pfet_01v8_lvt_60_0/GATE.t72 VDD.t37 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X539 sky130_asc_pfet_01v8_lvt_60_0/GATE.t181 VDD.t36 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X540 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t0 sky130_asc_pfet_01v8_lvt_60_0/GATE.t241 VDD.t35 VDD.t34 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X541 sky130_asc_pfet_01v8_lvt_60_0/GATE.t81 VDD.t10 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X542 vbg.t0 sky130_asc_pfet_01v8_lvt_60_0/GATE.t242 VDD.t33 VDD.t32 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X543 VSS.t231 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X544 sky130_asc_pfet_01v8_lvt_60_0/GATE.t73 VDD.t9 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X545 VDD.t31 sky130_asc_pfet_01v8_lvt_60_0/GATE.t243 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VDD.t30 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X546 VSS.t232 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X547 VSS.t2 porst.t8 sky130_asc_pfet_01v8_lvt_60_0/GATE.t1 VSS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=2e+06u
X548 sky130_asc_pfet_01v8_lvt_60_0/GATE.t75 VDD.t8 sky130_fd_pr__cap_mim_m3_1 l=2e+06u w=2e+06u
X549 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.t244 VDD.t7 VDD.t6 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6.45e+06u l=2e+06u
X550 VSS VSS.t16 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_fd_pr__pnp_05v5_W3p40L3p40
R0 sky130_asc_pfet_01v8_lvt_60_0/GATE.n105 sky130_asc_pfet_01v8_lvt_60_0/GATE.t5 243.258
R1 sky130_asc_pfet_01v8_lvt_60_0/GATE.n173 sky130_asc_pfet_01v8_lvt_60_0/GATE.t107 222.22
R2 sky130_asc_pfet_01v8_lvt_60_0/GATE.n12 sky130_asc_pfet_01v8_lvt_60_0/GATE.n11 195.413
R3 sky130_asc_pfet_01v8_lvt_60_0/GATE.n13 sky130_asc_pfet_01v8_lvt_60_0/GATE.n12 195.413
R4 sky130_asc_pfet_01v8_lvt_60_0/GATE.n14 sky130_asc_pfet_01v8_lvt_60_0/GATE.n13 195.413
R5 sky130_asc_pfet_01v8_lvt_60_0/GATE.n108 sky130_asc_pfet_01v8_lvt_60_0/GATE.n107 195.413
R6 sky130_asc_pfet_01v8_lvt_60_0/GATE.n107 sky130_asc_pfet_01v8_lvt_60_0/GATE.n106 195.413
R7 sky130_asc_pfet_01v8_lvt_60_0/GATE.n106 sky130_asc_pfet_01v8_lvt_60_0/GATE.n105 195.413
R8 sky130_asc_pfet_01v8_lvt_60_0/GATE.n644 sky130_asc_pfet_01v8_lvt_60_0/GATE.n643 195.413
R9 sky130_asc_pfet_01v8_lvt_60_0/GATE.n643 sky130_asc_pfet_01v8_lvt_60_0/GATE.n642 195.413
R10 sky130_asc_pfet_01v8_lvt_60_0/GATE.n642 sky130_asc_pfet_01v8_lvt_60_0/GATE.n641 195.413
R11 sky130_asc_pfet_01v8_lvt_60_0/GATE.n159 sky130_asc_pfet_01v8_lvt_60_0/GATE.t47 166.1
R12 sky130_asc_pfet_01v8_lvt_60_0/GATE.n183 sky130_asc_pfet_01v8_lvt_60_0/GATE.t95 166.1
R13 sky130_asc_pfet_01v8_lvt_60_0/GATE.n563 sky130_asc_pfet_01v8_lvt_60_0/GATE.t224 166.1
R14 sky130_asc_pfet_01v8_lvt_60_0/GATE.n379 sky130_asc_pfet_01v8_lvt_60_0/GATE.t111 166.1
R15 sky130_asc_pfet_01v8_lvt_60_0/GATE.n156 sky130_asc_pfet_01v8_lvt_60_0/GATE.t87 166.1
R16 sky130_asc_pfet_01v8_lvt_60_0/GATE.n101 sky130_asc_pfet_01v8_lvt_60_0/GATE.t64 166.1
R17 sky130_asc_pfet_01v8_lvt_60_0/GATE.n180 sky130_asc_pfet_01v8_lvt_60_0/GATE.t244 166.1
R18 sky130_asc_pfet_01v8_lvt_60_0/GATE.n172 sky130_asc_pfet_01v8_lvt_60_0/GATE.t32 166.1
R19 sky130_asc_pfet_01v8_lvt_60_0/GATE.n568 sky130_asc_pfet_01v8_lvt_60_0/GATE.t197 166.1
R20 sky130_asc_pfet_01v8_lvt_60_0/GATE.n561 sky130_asc_pfet_01v8_lvt_60_0/GATE.t227 166.1
R21 sky130_asc_pfet_01v8_lvt_60_0/GATE.n384 sky130_asc_pfet_01v8_lvt_60_0/GATE.t209 166.1
R22 sky130_asc_pfet_01v8_lvt_60_0/GATE.n377 sky130_asc_pfet_01v8_lvt_60_0/GATE.t138 166.1
R23 sky130_asc_pfet_01v8_lvt_60_0/GATE.n153 sky130_asc_pfet_01v8_lvt_60_0/GATE.t37 166.1
R24 sky130_asc_pfet_01v8_lvt_60_0/GATE.n177 sky130_asc_pfet_01v8_lvt_60_0/GATE.t68 166.1
R25 sky130_asc_pfet_01v8_lvt_60_0/GATE.n171 sky130_asc_pfet_01v8_lvt_60_0/GATE.t56 166.1
R26 sky130_asc_pfet_01v8_lvt_60_0/GATE.n571 sky130_asc_pfet_01v8_lvt_60_0/GATE.t25 166.1
R27 sky130_asc_pfet_01v8_lvt_60_0/GATE.n559 sky130_asc_pfet_01v8_lvt_60_0/GATE.t163 166.1
R28 sky130_asc_pfet_01v8_lvt_60_0/GATE.n387 sky130_asc_pfet_01v8_lvt_60_0/GATE.t170 166.1
R29 sky130_asc_pfet_01v8_lvt_60_0/GATE.n375 sky130_asc_pfet_01v8_lvt_60_0/GATE.t144 166.1
R30 sky130_asc_pfet_01v8_lvt_60_0/GATE.n97 sky130_asc_pfet_01v8_lvt_60_0/GATE.t241 166.1
R31 sky130_asc_pfet_01v8_lvt_60_0/GATE.n150 sky130_asc_pfet_01v8_lvt_60_0/GATE.t234 166.1
R32 sky130_asc_pfet_01v8_lvt_60_0/GATE.n174 sky130_asc_pfet_01v8_lvt_60_0/GATE.t67 166.1
R33 sky130_asc_pfet_01v8_lvt_60_0/GATE.n188 sky130_asc_pfet_01v8_lvt_60_0/GATE.t57 166.1
R34 sky130_asc_pfet_01v8_lvt_60_0/GATE.n574 sky130_asc_pfet_01v8_lvt_60_0/GATE.t186 166.1
R35 sky130_asc_pfet_01v8_lvt_60_0/GATE.n556 sky130_asc_pfet_01v8_lvt_60_0/GATE.t232 166.1
R36 sky130_asc_pfet_01v8_lvt_60_0/GATE.n390 sky130_asc_pfet_01v8_lvt_60_0/GATE.t169 166.1
R37 sky130_asc_pfet_01v8_lvt_60_0/GATE.n372 sky130_asc_pfet_01v8_lvt_60_0/GATE.t145 166.1
R38 sky130_asc_pfet_01v8_lvt_60_0/GATE.n94 sky130_asc_pfet_01v8_lvt_60_0/GATE.t226 166.099
R39 sky130_asc_pfet_01v8_lvt_60_0/GATE.n146 sky130_asc_pfet_01v8_lvt_60_0/GATE.t45 166.099
R40 sky130_asc_pfet_01v8_lvt_60_0/GATE.n193 sky130_asc_pfet_01v8_lvt_60_0/GATE.t230 166.099
R41 sky130_asc_pfet_01v8_lvt_60_0/GATE.n577 sky130_asc_pfet_01v8_lvt_60_0/GATE.t239 166.099
R42 sky130_asc_pfet_01v8_lvt_60_0/GATE.n553 sky130_asc_pfet_01v8_lvt_60_0/GATE.t174 166.099
R43 sky130_asc_pfet_01v8_lvt_60_0/GATE.n393 sky130_asc_pfet_01v8_lvt_60_0/GATE.t160 166.099
R44 sky130_asc_pfet_01v8_lvt_60_0/GATE.n369 sky130_asc_pfet_01v8_lvt_60_0/GATE.t182 166.099
R45 sky130_asc_pfet_01v8_lvt_60_0/GATE.n91 sky130_asc_pfet_01v8_lvt_60_0/GATE.t28 166.098
R46 sky130_asc_pfet_01v8_lvt_60_0/GATE.n196 sky130_asc_pfet_01v8_lvt_60_0/GATE.t96 166.098
R47 sky130_asc_pfet_01v8_lvt_60_0/GATE.n550 sky130_asc_pfet_01v8_lvt_60_0/GATE.t176 166.098
R48 sky130_asc_pfet_01v8_lvt_60_0/GATE.n366 sky130_asc_pfet_01v8_lvt_60_0/GATE.t99 166.098
R49 sky130_asc_pfet_01v8_lvt_60_0/GATE.n88 sky130_asc_pfet_01v8_lvt_60_0/GATE.t30 166.098
R50 sky130_asc_pfet_01v8_lvt_60_0/GATE.n199 sky130_asc_pfet_01v8_lvt_60_0/GATE.t58 166.098
R51 sky130_asc_pfet_01v8_lvt_60_0/GATE.n547 sky130_asc_pfet_01v8_lvt_60_0/GATE.t212 166.098
R52 sky130_asc_pfet_01v8_lvt_60_0/GATE.n363 sky130_asc_pfet_01v8_lvt_60_0/GATE.t120 166.098
R53 sky130_asc_pfet_01v8_lvt_60_0/GATE.n84 sky130_asc_pfet_01v8_lvt_60_0/GATE.t202 166.097
R54 sky130_asc_pfet_01v8_lvt_60_0/GATE.n202 sky130_asc_pfet_01v8_lvt_60_0/GATE.t59 166.097
R55 sky130_asc_pfet_01v8_lvt_60_0/GATE.n542 sky130_asc_pfet_01v8_lvt_60_0/GATE.t229 166.097
R56 sky130_asc_pfet_01v8_lvt_60_0/GATE.n358 sky130_asc_pfet_01v8_lvt_60_0/GATE.t104 166.097
R57 sky130_asc_pfet_01v8_lvt_60_0/GATE.n170 sky130_asc_pfet_01v8_lvt_60_0/GATE.t78 166.095
R58 sky130_asc_pfet_01v8_lvt_60_0/GATE.n540 sky130_asc_pfet_01v8_lvt_60_0/GATE.t83 166.095
R59 sky130_asc_pfet_01v8_lvt_60_0/GATE.n356 sky130_asc_pfet_01v8_lvt_60_0/GATE.t126 166.095
R60 sky130_asc_pfet_01v8_lvt_60_0/GATE.n169 sky130_asc_pfet_01v8_lvt_60_0/GATE.t231 166.094
R61 sky130_asc_pfet_01v8_lvt_60_0/GATE.n538 sky130_asc_pfet_01v8_lvt_60_0/GATE.t236 166.094
R62 sky130_asc_pfet_01v8_lvt_60_0/GATE.n354 sky130_asc_pfet_01v8_lvt_60_0/GATE.t152 166.094
R63 sky130_asc_pfet_01v8_lvt_60_0/GATE.n208 sky130_asc_pfet_01v8_lvt_60_0/GATE.t84 166.093
R64 sky130_asc_pfet_01v8_lvt_60_0/GATE.n535 sky130_asc_pfet_01v8_lvt_60_0/GATE.t39 166.093
R65 sky130_asc_pfet_01v8_lvt_60_0/GATE.n351 sky130_asc_pfet_01v8_lvt_60_0/GATE.t187 166.093
R66 sky130_asc_pfet_01v8_lvt_60_0/GATE.n213 sky130_asc_pfet_01v8_lvt_60_0/GATE.t41 166.091
R67 sky130_asc_pfet_01v8_lvt_60_0/GATE.n532 sky130_asc_pfet_01v8_lvt_60_0/GATE.t214 166.091
R68 sky130_asc_pfet_01v8_lvt_60_0/GATE.n348 sky130_asc_pfet_01v8_lvt_60_0/GATE.t189 166.091
R69 sky130_asc_pfet_01v8_lvt_60_0/GATE.n580 sky130_asc_pfet_01v8_lvt_60_0/GATE.t42 166.089
R70 sky130_asc_pfet_01v8_lvt_60_0/GATE.n529 sky130_asc_pfet_01v8_lvt_60_0/GATE.t215 166.089
R71 sky130_asc_pfet_01v8_lvt_60_0/GATE.n345 sky130_asc_pfet_01v8_lvt_60_0/GATE.t198 166.089
R72 sky130_asc_pfet_01v8_lvt_60_0/GATE.n582 sky130_asc_pfet_01v8_lvt_60_0/GATE.t216 166.087
R73 sky130_asc_pfet_01v8_lvt_60_0/GATE.n526 sky130_asc_pfet_01v8_lvt_60_0/GATE.t65 166.087
R74 sky130_asc_pfet_01v8_lvt_60_0/GATE.n342 sky130_asc_pfet_01v8_lvt_60_0/GATE.t200 166.087
R75 sky130_asc_pfet_01v8_lvt_60_0/GATE.n585 sky130_asc_pfet_01v8_lvt_60_0/GATE.t217 166.085
R76 sky130_asc_pfet_01v8_lvt_60_0/GATE.n521 sky130_asc_pfet_01v8_lvt_60_0/GATE.t221 166.085
R77 sky130_asc_pfet_01v8_lvt_60_0/GATE.n337 sky130_asc_pfet_01v8_lvt_60_0/GATE.t129 166.085
R78 sky130_asc_pfet_01v8_lvt_60_0/GATE.n83 sky130_asc_pfet_01v8_lvt_60_0/GATE.t69 166.083
R79 sky130_asc_pfet_01v8_lvt_60_0/GATE.n519 sky130_asc_pfet_01v8_lvt_60_0/GATE.t242 166.083
R80 sky130_asc_pfet_01v8_lvt_60_0/GATE.n335 sky130_asc_pfet_01v8_lvt_60_0/GATE.t165 166.083
R81 sky130_asc_pfet_01v8_lvt_60_0/GATE.n82 sky130_asc_pfet_01v8_lvt_60_0/GATE.t222 166.08
R82 sky130_asc_pfet_01v8_lvt_60_0/GATE.n517 sky130_asc_pfet_01v8_lvt_60_0/GATE.t154 166.08
R83 sky130_asc_pfet_01v8_lvt_60_0/GATE.n333 sky130_asc_pfet_01v8_lvt_60_0/GATE.t166 166.08
R84 sky130_asc_pfet_01v8_lvt_60_0/GATE.n590 sky130_asc_pfet_01v8_lvt_60_0/GATE.t24 166.078
R85 sky130_asc_pfet_01v8_lvt_60_0/GATE.n514 sky130_asc_pfet_01v8_lvt_60_0/GATE.t192 166.078
R86 sky130_asc_pfet_01v8_lvt_60_0/GATE.n330 sky130_asc_pfet_01v8_lvt_60_0/GATE.t175 166.078
R87 sky130_asc_pfet_01v8_lvt_60_0/GATE.n595 sky130_asc_pfet_01v8_lvt_60_0/GATE.t158 166.075
R88 sky130_asc_pfet_01v8_lvt_60_0/GATE.n511 sky130_asc_pfet_01v8_lvt_60_0/GATE.t168 166.075
R89 sky130_asc_pfet_01v8_lvt_60_0/GATE.n327 sky130_asc_pfet_01v8_lvt_60_0/GATE.t178 166.075
R90 sky130_asc_pfet_01v8_lvt_60_0/GATE.n598 sky130_asc_pfet_01v8_lvt_60_0/GATE.t196 166.072
R91 sky130_asc_pfet_01v8_lvt_60_0/GATE.n508 sky130_asc_pfet_01v8_lvt_60_0/GATE.t204 166.072
R92 sky130_asc_pfet_01v8_lvt_60_0/GATE.n324 sky130_asc_pfet_01v8_lvt_60_0/GATE.t114 166.072
R93 sky130_asc_pfet_01v8_lvt_60_0/GATE.n601 sky130_asc_pfet_01v8_lvt_60_0/GATE.t171 166.068
R94 sky130_asc_pfet_01v8_lvt_60_0/GATE.n505 sky130_asc_pfet_01v8_lvt_60_0/GATE.t206 166.068
R95 sky130_asc_pfet_01v8_lvt_60_0/GATE.n321 sky130_asc_pfet_01v8_lvt_60_0/GATE.t116 166.068
R96 sky130_asc_pfet_01v8_lvt_60_0/GATE.n604 sky130_asc_pfet_01v8_lvt_60_0/GATE.t208 166.065
R97 sky130_asc_pfet_01v8_lvt_60_0/GATE.n500 sky130_asc_pfet_01v8_lvt_60_0/GATE.t133 166.065
R98 sky130_asc_pfet_01v8_lvt_60_0/GATE.n316 sky130_asc_pfet_01v8_lvt_60_0/GATE.t79 166.065
R99 sky130_asc_pfet_01v8_lvt_60_0/GATE.n81 sky130_asc_pfet_01v8_lvt_60_0/GATE.t211 166.061
R100 sky130_asc_pfet_01v8_lvt_60_0/GATE.n498 sky130_asc_pfet_01v8_lvt_60_0/GATE.t135 166.061
R101 sky130_asc_pfet_01v8_lvt_60_0/GATE.n314 sky130_asc_pfet_01v8_lvt_60_0/GATE.t121 166.061
R102 sky130_asc_pfet_01v8_lvt_60_0/GATE.n80 sky130_asc_pfet_01v8_lvt_60_0/GATE.t137 166.057
R103 sky130_asc_pfet_01v8_lvt_60_0/GATE.n312 sky130_asc_pfet_01v8_lvt_60_0/GATE.t150 166.057
R104 sky130_asc_pfet_01v8_lvt_60_0/GATE.n609 sky130_asc_pfet_01v8_lvt_60_0/GATE.t173 166.053
R105 sky130_asc_pfet_01v8_lvt_60_0/GATE.n487 sky130_asc_pfet_01v8_lvt_60_0/GATE.t179 166.053
R106 sky130_asc_pfet_01v8_lvt_60_0/GATE.n309 sky130_asc_pfet_01v8_lvt_60_0/GATE.t85 166.053
R107 sky130_asc_pfet_01v8_lvt_60_0/GATE.n614 sky130_asc_pfet_01v8_lvt_60_0/GATE.t146 166.048
R108 sky130_asc_pfet_01v8_lvt_60_0/GATE.n484 sky130_asc_pfet_01v8_lvt_60_0/GATE.t180 166.048
R109 sky130_asc_pfet_01v8_lvt_60_0/GATE.n306 sky130_asc_pfet_01v8_lvt_60_0/GATE.t102 166.048
R110 sky130_asc_pfet_01v8_lvt_60_0/GATE.n617 sky130_asc_pfet_01v8_lvt_60_0/GATE.t183 166.043
R111 sky130_asc_pfet_01v8_lvt_60_0/GATE.n481 sky130_asc_pfet_01v8_lvt_60_0/GATE.t117 166.043
R112 sky130_asc_pfet_01v8_lvt_60_0/GATE.n303 sky130_asc_pfet_01v8_lvt_60_0/GATE.t63 166.043
R113 sky130_asc_pfet_01v8_lvt_60_0/GATE.n620 sky130_asc_pfet_01v8_lvt_60_0/GATE.t60 166.038
R114 sky130_asc_pfet_01v8_lvt_60_0/GATE.n478 sky130_asc_pfet_01v8_lvt_60_0/GATE.t119 166.038
R115 sky130_asc_pfet_01v8_lvt_60_0/GATE.n300 sky130_asc_pfet_01v8_lvt_60_0/GATE.t108 166.038
R116 sky130_asc_pfet_01v8_lvt_60_0/GATE.n623 sky130_asc_pfet_01v8_lvt_60_0/GATE.t233 166.033
R117 sky130_asc_pfet_01v8_lvt_60_0/GATE.n473 sky130_asc_pfet_01v8_lvt_60_0/GATE.t123 166.033
R118 sky130_asc_pfet_01v8_lvt_60_0/GATE.n295 sky130_asc_pfet_01v8_lvt_60_0/GATE.t70 166.033
R119 sky130_asc_pfet_01v8_lvt_60_0/GATE.n79 sky130_asc_pfet_01v8_lvt_60_0/GATE.t235 166.027
R120 sky130_asc_pfet_01v8_lvt_60_0/GATE.n471 sky130_asc_pfet_01v8_lvt_60_0/GATE.t237 166.027
R121 sky130_asc_pfet_01v8_lvt_60_0/GATE.n293 sky130_asc_pfet_01v8_lvt_60_0/GATE.t71 166.027
R122 sky130_asc_pfet_01v8_lvt_60_0/GATE.n78 sky130_asc_pfet_01v8_lvt_60_0/GATE.t238 166.021
R123 sky130_asc_pfet_01v8_lvt_60_0/GATE.n469 sky130_asc_pfet_01v8_lvt_60_0/GATE.t184 166.021
R124 sky130_asc_pfet_01v8_lvt_60_0/GATE.n291 sky130_asc_pfet_01v8_lvt_60_0/GATE.t91 166.021
R125 sky130_asc_pfet_01v8_lvt_60_0/GATE.n77 sky130_asc_pfet_01v8_lvt_60_0/GATE.t240 166.014
R126 sky130_asc_pfet_01v8_lvt_60_0/GATE.n467 sky130_asc_pfet_01v8_lvt_60_0/GATE.t185 166.014
R127 sky130_asc_pfet_01v8_lvt_60_0/GATE.n289 sky130_asc_pfet_01v8_lvt_60_0/GATE.t105 166.014
R128 sky130_asc_pfet_01v8_lvt_60_0/GATE.n635 sky130_asc_pfet_01v8_lvt_60_0/GATE.t188 166.007
R129 sky130_asc_pfet_01v8_lvt_60_0/GATE.n464 sky130_asc_pfet_01v8_lvt_60_0/GATE.t218 166.007
R130 sky130_asc_pfet_01v8_lvt_60_0/GATE.n286 sky130_asc_pfet_01v8_lvt_60_0/GATE.t205 166.007
R131 sky130_asc_pfet_01v8_lvt_60_0/GATE.n637 sky130_asc_pfet_01v8_lvt_60_0/GATE.t190 165.999
R132 sky130_asc_pfet_01v8_lvt_60_0/GATE.n461 sky130_asc_pfet_01v8_lvt_60_0/GATE.t195 165.999
R133 sky130_asc_pfet_01v8_lvt_60_0/GATE.n283 sky130_asc_pfet_01v8_lvt_60_0/GATE.t110 165.999
R134 sky130_asc_pfet_01v8_lvt_60_0/GATE.n634 sky130_asc_pfet_01v8_lvt_60_0/GATE.t220 165.992
R135 sky130_asc_pfet_01v8_lvt_60_0/GATE.n458 sky130_asc_pfet_01v8_lvt_60_0/GATE.t223 165.992
R136 sky130_asc_pfet_01v8_lvt_60_0/GATE.n280 sky130_asc_pfet_01v8_lvt_60_0/GATE.t134 165.992
R137 sky130_asc_pfet_01v8_lvt_60_0/GATE.n632 sky130_asc_pfet_01v8_lvt_60_0/GATE.t225 165.983
R138 sky130_asc_pfet_01v8_lvt_60_0/GATE.n455 sky130_asc_pfet_01v8_lvt_60_0/GATE.t159 165.983
R139 sky130_asc_pfet_01v8_lvt_60_0/GATE.n277 sky130_asc_pfet_01v8_lvt_60_0/GATE.t136 165.983
R140 sky130_asc_pfet_01v8_lvt_60_0/GATE.n72 sky130_asc_pfet_01v8_lvt_60_0/GATE.t228 165.974
R141 sky130_asc_pfet_01v8_lvt_60_0/GATE.n451 sky130_asc_pfet_01v8_lvt_60_0/GATE.t161 165.974
R142 sky130_asc_pfet_01v8_lvt_60_0/GATE.n273 sky130_asc_pfet_01v8_lvt_60_0/GATE.t94 165.974
R143 sky130_asc_pfet_01v8_lvt_60_0/GATE.n70 sky130_asc_pfet_01v8_lvt_60_0/GATE.t164 165.965
R144 sky130_asc_pfet_01v8_lvt_60_0/GATE.n449 sky130_asc_pfet_01v8_lvt_60_0/GATE.t199 165.965
R145 sky130_asc_pfet_01v8_lvt_60_0/GATE.n271 sky130_asc_pfet_01v8_lvt_60_0/GATE.t143 165.965
R146 sky130_asc_pfet_01v8_lvt_60_0/GATE.n68 sky130_asc_pfet_01v8_lvt_60_0/GATE.t167 165.954
R147 sky130_asc_pfet_01v8_lvt_60_0/GATE.n447 sky130_asc_pfet_01v8_lvt_60_0/GATE.t172 165.954
R148 sky130_asc_pfet_01v8_lvt_60_0/GATE.n269 sky130_asc_pfet_01v8_lvt_60_0/GATE.t98 165.954
R149 sky130_asc_pfet_01v8_lvt_60_0/GATE.n65 sky130_asc_pfet_01v8_lvt_60_0/GATE.t203 165.943
R150 sky130_asc_pfet_01v8_lvt_60_0/GATE.n444 sky130_asc_pfet_01v8_lvt_60_0/GATE.t210 165.943
R151 sky130_asc_pfet_01v8_lvt_60_0/GATE.n266 sky130_asc_pfet_01v8_lvt_60_0/GATE.t118 165.943
R152 sky130_asc_pfet_01v8_lvt_60_0/GATE.n62 sky130_asc_pfet_01v8_lvt_60_0/GATE.t177 165.932
R153 sky130_asc_pfet_01v8_lvt_60_0/GATE.n441 sky130_asc_pfet_01v8_lvt_60_0/GATE.t112 165.932
R154 sky130_asc_pfet_01v8_lvt_60_0/GATE.n263 sky130_asc_pfet_01v8_lvt_60_0/GATE.t61 165.932
R155 sky130_asc_pfet_01v8_lvt_60_0/GATE.n59 sky130_asc_pfet_01v8_lvt_60_0/GATE.t213 165.919
R156 sky130_asc_pfet_01v8_lvt_60_0/GATE.n438 sky130_asc_pfet_01v8_lvt_60_0/GATE.t139 165.919
R157 sky130_asc_pfet_01v8_lvt_60_0/GATE.n260 sky130_asc_pfet_01v8_lvt_60_0/GATE.t82 165.919
R158 sky130_asc_pfet_01v8_lvt_60_0/GATE.n56 sky130_asc_pfet_01v8_lvt_60_0/GATE.t115 165.906
R159 sky130_asc_pfet_01v8_lvt_60_0/GATE.n435 sky130_asc_pfet_01v8_lvt_60_0/GATE.t76 165.906
R160 sky130_asc_pfet_01v8_lvt_60_0/GATE.n257 sky130_asc_pfet_01v8_lvt_60_0/GATE.t125 165.906
R161 sky130_asc_pfet_01v8_lvt_60_0/GATE.n51 sky130_asc_pfet_01v8_lvt_60_0/GATE.t141 165.891
R162 sky130_asc_pfet_01v8_lvt_60_0/GATE.n430 sky130_asc_pfet_01v8_lvt_60_0/GATE.t148 165.891
R163 sky130_asc_pfet_01v8_lvt_60_0/GATE.n252 sky130_asc_pfet_01v8_lvt_60_0/GATE.t86 165.891
R164 sky130_asc_pfet_01v8_lvt_60_0/GATE.n49 sky130_asc_pfet_01v8_lvt_60_0/GATE.t80 165.876
R165 sky130_asc_pfet_01v8_lvt_60_0/GATE.n428 sky130_asc_pfet_01v8_lvt_60_0/GATE.t149 165.876
R166 sky130_asc_pfet_01v8_lvt_60_0/GATE.n250 sky130_asc_pfet_01v8_lvt_60_0/GATE.t88 165.876
R167 sky130_asc_pfet_01v8_lvt_60_0/GATE.n47 sky130_asc_pfet_01v8_lvt_60_0/GATE.t151 165.859
R168 sky130_asc_pfet_01v8_lvt_60_0/GATE.n426 sky130_asc_pfet_01v8_lvt_60_0/GATE.t100 165.859
R169 sky130_asc_pfet_01v8_lvt_60_0/GATE.n248 sky130_asc_pfet_01v8_lvt_60_0/GATE.t48 165.859
R170 sky130_asc_pfet_01v8_lvt_60_0/GATE.n44 sky130_asc_pfet_01v8_lvt_60_0/GATE.t153 165.841
R171 sky130_asc_pfet_01v8_lvt_60_0/GATE.n423 sky130_asc_pfet_01v8_lvt_60_0/GATE.t101 165.841
R172 sky130_asc_pfet_01v8_lvt_60_0/GATE.n245 sky130_asc_pfet_01v8_lvt_60_0/GATE.t49 165.841
R173 sky130_asc_pfet_01v8_lvt_60_0/GATE.n41 sky130_asc_pfet_01v8_lvt_60_0/GATE.t103 165.822
R174 sky130_asc_pfet_01v8_lvt_60_0/GATE.n420 sky130_asc_pfet_01v8_lvt_60_0/GATE.t62 165.822
R175 sky130_asc_pfet_01v8_lvt_60_0/GATE.n242 sky130_asc_pfet_01v8_lvt_60_0/GATE.t52 165.822
R176 sky130_asc_pfet_01v8_lvt_60_0/GATE.n38 sky130_asc_pfet_01v8_lvt_60_0/GATE.t122 165.801
R177 sky130_asc_pfet_01v8_lvt_60_0/GATE.n417 sky130_asc_pfet_01v8_lvt_60_0/GATE.t128 165.801
R178 sky130_asc_pfet_01v8_lvt_60_0/GATE.n239 sky130_asc_pfet_01v8_lvt_60_0/GATE.t53 165.801
R179 sky130_asc_pfet_01v8_lvt_60_0/GATE.n35 sky130_asc_pfet_01v8_lvt_60_0/GATE.t147 165.777
R180 sky130_asc_pfet_01v8_lvt_60_0/GATE.n414 sky130_asc_pfet_01v8_lvt_60_0/GATE.t66 165.777
R181 sky130_asc_pfet_01v8_lvt_60_0/GATE.n236 sky130_asc_pfet_01v8_lvt_60_0/GATE.t74 165.777
R182 sky130_asc_pfet_01v8_lvt_60_0/GATE.n30 sky130_asc_pfet_01v8_lvt_60_0/GATE.t243 165.752
R183 sky130_asc_pfet_01v8_lvt_60_0/GATE.n409 sky130_asc_pfet_01v8_lvt_60_0/GATE.t90 165.752
R184 sky130_asc_pfet_01v8_lvt_60_0/GATE.n231 sky130_asc_pfet_01v8_lvt_60_0/GATE.t29 165.752
R185 sky130_asc_pfet_01v8_lvt_60_0/GATE.n28 sky130_asc_pfet_01v8_lvt_60_0/GATE.t156 165.725
R186 sky130_asc_pfet_01v8_lvt_60_0/GATE.n407 sky130_asc_pfet_01v8_lvt_60_0/GATE.t191 165.725
R187 sky130_asc_pfet_01v8_lvt_60_0/GATE.n229 sky130_asc_pfet_01v8_lvt_60_0/GATE.t31 165.725
R188 sky130_asc_pfet_01v8_lvt_60_0/GATE.n26 sky130_asc_pfet_01v8_lvt_60_0/GATE.t193 165.694
R189 sky130_asc_pfet_01v8_lvt_60_0/GATE.n405 sky130_asc_pfet_01v8_lvt_60_0/GATE.t124 165.694
R190 sky130_asc_pfet_01v8_lvt_60_0/GATE.n227 sky130_asc_pfet_01v8_lvt_60_0/GATE.t35 165.694
R191 sky130_asc_pfet_01v8_lvt_60_0/GATE.n23 sky130_asc_pfet_01v8_lvt_60_0/GATE.t194 165.661
R192 sky130_asc_pfet_01v8_lvt_60_0/GATE.n402 sky130_asc_pfet_01v8_lvt_60_0/GATE.t201 165.661
R193 sky130_asc_pfet_01v8_lvt_60_0/GATE.n224 sky130_asc_pfet_01v8_lvt_60_0/GATE.t113 165.661
R194 sky130_asc_pfet_01v8_lvt_60_0/GATE.n20 sky130_asc_pfet_01v8_lvt_60_0/GATE.t127 165.623
R195 sky130_asc_pfet_01v8_lvt_60_0/GATE.n399 sky130_asc_pfet_01v8_lvt_60_0/GATE.t131 165.623
R196 sky130_asc_pfet_01v8_lvt_60_0/GATE.n221 sky130_asc_pfet_01v8_lvt_60_0/GATE.t140 165.623
R197 sky130_asc_pfet_01v8_lvt_60_0/GATE.n17 sky130_asc_pfet_01v8_lvt_60_0/GATE.t207 165.582
R198 sky130_asc_pfet_01v8_lvt_60_0/GATE.n396 sky130_asc_pfet_01v8_lvt_60_0/GATE.t132 165.582
R199 sky130_asc_pfet_01v8_lvt_60_0/GATE.n218 sky130_asc_pfet_01v8_lvt_60_0/GATE.t77 165.582
R200 sky130_asc_pfet_01v8_lvt_60_0/GATE.n166 sky130_asc_pfet_01v8_lvt_60_0/GATE.t219 165.297
R201 sky130_asc_pfet_01v8_lvt_60_0/GATE.n492 sky130_asc_pfet_01v8_lvt_60_0/GATE.t142 163.403
R202 sky130_asc_pfet_01v8_lvt_60_0/GATE.n15 sky130_asc_pfet_01v8_lvt_60_0/GATE.t16 137.018
R203 sky130_asc_pfet_01v8_lvt_60_0/GATE.n176 sky130_asc_pfet_01v8_lvt_60_0/GATE.n173 122.204
R204 sky130_asc_pfet_01v8_lvt_60_0/GATE.n633 sky130_asc_pfet_01v8_lvt_60_0/GATE.n632 107.968
R205 sky130_asc_pfet_01v8_lvt_60_0/GATE.n636 sky130_asc_pfet_01v8_lvt_60_0/GATE.n635 107.968
R206 sky130_asc_pfet_01v8_lvt_60_0/GATE.n456 sky130_asc_pfet_01v8_lvt_60_0/GATE.n455 107.968
R207 sky130_asc_pfet_01v8_lvt_60_0/GATE.n278 sky130_asc_pfet_01v8_lvt_60_0/GATE.n277 107.968
R208 sky130_asc_pfet_01v8_lvt_60_0/GATE.n15 sky130_asc_pfet_01v8_lvt_60_0/GATE.n14 106.24
R209 sky130_asc_pfet_01v8_lvt_60_0/GATE.n57 sky130_asc_pfet_01v8_lvt_60_0/GATE.n56 104.112
R210 sky130_asc_pfet_01v8_lvt_60_0/GATE.n615 sky130_asc_pfet_01v8_lvt_60_0/GATE.n614 104.112
R211 sky130_asc_pfet_01v8_lvt_60_0/GATE.n436 sky130_asc_pfet_01v8_lvt_60_0/GATE.n435 104.112
R212 sky130_asc_pfet_01v8_lvt_60_0/GATE.n258 sky130_asc_pfet_01v8_lvt_60_0/GATE.n257 104.112
R213 sky130_asc_pfet_01v8_lvt_60_0/GATE.n36 sky130_asc_pfet_01v8_lvt_60_0/GATE.n35 100.256
R214 sky130_asc_pfet_01v8_lvt_60_0/GATE.n596 sky130_asc_pfet_01v8_lvt_60_0/GATE.n595 100.256
R215 sky130_asc_pfet_01v8_lvt_60_0/GATE.n569 sky130_asc_pfet_01v8_lvt_60_0/GATE.n568 100.256
R216 sky130_asc_pfet_01v8_lvt_60_0/GATE.n415 sky130_asc_pfet_01v8_lvt_60_0/GATE.n414 100.256
R217 sky130_asc_pfet_01v8_lvt_60_0/GATE.n385 sky130_asc_pfet_01v8_lvt_60_0/GATE.n384 100.256
R218 sky130_asc_pfet_01v8_lvt_60_0/GATE.n237 sky130_asc_pfet_01v8_lvt_60_0/GATE.n236 100.256
R219 sky130_asc_pfet_01v8_lvt_60_0/GATE.n89 sky130_asc_pfet_01v8_lvt_60_0/GATE.n88 96.4
R220 sky130_asc_pfet_01v8_lvt_60_0/GATE.n214 sky130_asc_pfet_01v8_lvt_60_0/GATE.n213 96.4
R221 sky130_asc_pfet_01v8_lvt_60_0/GATE.n548 sky130_asc_pfet_01v8_lvt_60_0/GATE.n547 96.4
R222 sky130_asc_pfet_01v8_lvt_60_0/GATE.n364 sky130_asc_pfet_01v8_lvt_60_0/GATE.n363 96.4
R223 sky130_asc_pfet_01v8_lvt_60_0/GATE.n147 sky130_asc_pfet_01v8_lvt_60_0/GATE.n146 95.28
R224 sky130_asc_pfet_01v8_lvt_60_0/GATE.n578 sky130_asc_pfet_01v8_lvt_60_0/GATE.n577 95.28
R225 sky130_asc_pfet_01v8_lvt_60_0/GATE.n394 sky130_asc_pfet_01v8_lvt_60_0/GATE.n393 95.28
R226 sky130_asc_pfet_01v8_lvt_60_0/GATE.n194 sky130_asc_pfet_01v8_lvt_60_0/GATE.n193 92.544
R227 sky130_asc_pfet_01v8_lvt_60_0/GATE.n582 sky130_asc_pfet_01v8_lvt_60_0/GATE.n581 92.544
R228 sky130_asc_pfet_01v8_lvt_60_0/GATE.n527 sky130_asc_pfet_01v8_lvt_60_0/GATE.n526 92.544
R229 sky130_asc_pfet_01v8_lvt_60_0/GATE.n343 sky130_asc_pfet_01v8_lvt_60_0/GATE.n342 92.544
R230 sky130_asc_pfet_01v8_lvt_60_0/GATE.n11 sky130_asc_nfet_01v8_lvt_9_1/DRAIN 91.306
R231 sky130_asc_pfet_01v8_lvt_60_0/GATE.n108 sky130_asc_nfet_01v8_lvt_9_0/DRAIN 91.306
R232 sky130_asc_pfet_01v8_lvt_60_0/GATE.n151 sky130_asc_pfet_01v8_lvt_60_0/GATE.n150 88.688
R233 sky130_asc_pfet_01v8_lvt_60_0/GATE.n175 sky130_asc_pfet_01v8_lvt_60_0/GATE.n174 88.688
R234 sky130_asc_pfet_01v8_lvt_60_0/GATE.n506 sky130_asc_pfet_01v8_lvt_60_0/GATE.n505 88.688
R235 sky130_asc_pfet_01v8_lvt_60_0/GATE.n322 sky130_asc_pfet_01v8_lvt_60_0/GATE.n321 88.688
R236 sky130_asc_pfet_01v8_lvt_60_0/GATE.n85 sky130_asc_pfet_01v8_lvt_60_0/GATE.n84 87.568
R237 sky130_asc_pfet_01v8_lvt_60_0/GATE.n87 sky130_asc_pfet_01v8_lvt_60_0/GATE.n85 85.333
R238 sky130_asc_pfet_01v8_lvt_60_0/GATE.n90 sky130_asc_pfet_01v8_lvt_60_0/GATE.n87 85.333
R239 sky130_asc_pfet_01v8_lvt_60_0/GATE.n93 sky130_asc_pfet_01v8_lvt_60_0/GATE.n90 85.333
R240 sky130_asc_pfet_01v8_lvt_60_0/GATE.n96 sky130_asc_pfet_01v8_lvt_60_0/GATE.n93 85.333
R241 sky130_asc_pfet_01v8_lvt_60_0/GATE.n99 sky130_asc_pfet_01v8_lvt_60_0/GATE.n96 85.333
R242 sky130_asc_pfet_01v8_lvt_60_0/GATE.n162 sky130_asc_pfet_01v8_lvt_60_0/GATE.n161 85.333
R243 sky130_asc_pfet_01v8_lvt_60_0/GATE.n161 sky130_asc_pfet_01v8_lvt_60_0/GATE.n158 85.333
R244 sky130_asc_pfet_01v8_lvt_60_0/GATE.n158 sky130_asc_pfet_01v8_lvt_60_0/GATE.n155 85.333
R245 sky130_asc_pfet_01v8_lvt_60_0/GATE.n155 sky130_asc_pfet_01v8_lvt_60_0/GATE.n152 85.333
R246 sky130_asc_pfet_01v8_lvt_60_0/GATE.n152 sky130_asc_pfet_01v8_lvt_60_0/GATE.n149 85.333
R247 sky130_asc_pfet_01v8_lvt_60_0/GATE.n149 sky130_asc_pfet_01v8_lvt_60_0/GATE.n147 85.333
R248 sky130_asc_pfet_01v8_lvt_60_0/GATE.n398 sky130_asc_pfet_01v8_lvt_60_0/GATE.n395 85.333
R249 sky130_asc_pfet_01v8_lvt_60_0/GATE.n401 sky130_asc_pfet_01v8_lvt_60_0/GATE.n398 85.333
R250 sky130_asc_pfet_01v8_lvt_60_0/GATE.n404 sky130_asc_pfet_01v8_lvt_60_0/GATE.n401 85.333
R251 sky130_asc_pfet_01v8_lvt_60_0/GATE.n406 sky130_asc_pfet_01v8_lvt_60_0/GATE.n404 85.333
R252 sky130_asc_pfet_01v8_lvt_60_0/GATE.n408 sky130_asc_pfet_01v8_lvt_60_0/GATE.n406 85.333
R253 sky130_asc_pfet_01v8_lvt_60_0/GATE.n411 sky130_asc_pfet_01v8_lvt_60_0/GATE.n408 85.333
R254 sky130_asc_pfet_01v8_lvt_60_0/GATE.n413 sky130_asc_pfet_01v8_lvt_60_0/GATE.n411 85.333
R255 sky130_asc_pfet_01v8_lvt_60_0/GATE.n416 sky130_asc_pfet_01v8_lvt_60_0/GATE.n413 85.333
R256 sky130_asc_pfet_01v8_lvt_60_0/GATE.n419 sky130_asc_pfet_01v8_lvt_60_0/GATE.n416 85.333
R257 sky130_asc_pfet_01v8_lvt_60_0/GATE.n422 sky130_asc_pfet_01v8_lvt_60_0/GATE.n419 85.333
R258 sky130_asc_pfet_01v8_lvt_60_0/GATE.n425 sky130_asc_pfet_01v8_lvt_60_0/GATE.n422 85.333
R259 sky130_asc_pfet_01v8_lvt_60_0/GATE.n427 sky130_asc_pfet_01v8_lvt_60_0/GATE.n425 85.333
R260 sky130_asc_pfet_01v8_lvt_60_0/GATE.n429 sky130_asc_pfet_01v8_lvt_60_0/GATE.n427 85.333
R261 sky130_asc_pfet_01v8_lvt_60_0/GATE.n432 sky130_asc_pfet_01v8_lvt_60_0/GATE.n429 85.333
R262 sky130_asc_pfet_01v8_lvt_60_0/GATE.n434 sky130_asc_pfet_01v8_lvt_60_0/GATE.n432 85.333
R263 sky130_asc_pfet_01v8_lvt_60_0/GATE.n437 sky130_asc_pfet_01v8_lvt_60_0/GATE.n434 85.333
R264 sky130_asc_pfet_01v8_lvt_60_0/GATE.n440 sky130_asc_pfet_01v8_lvt_60_0/GATE.n437 85.333
R265 sky130_asc_pfet_01v8_lvt_60_0/GATE.n443 sky130_asc_pfet_01v8_lvt_60_0/GATE.n440 85.333
R266 sky130_asc_pfet_01v8_lvt_60_0/GATE.n446 sky130_asc_pfet_01v8_lvt_60_0/GATE.n443 85.333
R267 sky130_asc_pfet_01v8_lvt_60_0/GATE.n448 sky130_asc_pfet_01v8_lvt_60_0/GATE.n446 85.333
R268 sky130_asc_pfet_01v8_lvt_60_0/GATE.n450 sky130_asc_pfet_01v8_lvt_60_0/GATE.n448 85.333
R269 sky130_asc_pfet_01v8_lvt_60_0/GATE.n452 sky130_asc_pfet_01v8_lvt_60_0/GATE.n450 85.333
R270 sky130_asc_pfet_01v8_lvt_60_0/GATE.n454 sky130_asc_pfet_01v8_lvt_60_0/GATE.n452 85.333
R271 sky130_asc_pfet_01v8_lvt_60_0/GATE.n457 sky130_asc_pfet_01v8_lvt_60_0/GATE.n454 85.333
R272 sky130_asc_pfet_01v8_lvt_60_0/GATE.n460 sky130_asc_pfet_01v8_lvt_60_0/GATE.n457 85.333
R273 sky130_asc_pfet_01v8_lvt_60_0/GATE.n463 sky130_asc_pfet_01v8_lvt_60_0/GATE.n460 85.333
R274 sky130_asc_pfet_01v8_lvt_60_0/GATE.n466 sky130_asc_pfet_01v8_lvt_60_0/GATE.n463 85.333
R275 sky130_asc_pfet_01v8_lvt_60_0/GATE.n468 sky130_asc_pfet_01v8_lvt_60_0/GATE.n466 85.333
R276 sky130_asc_pfet_01v8_lvt_60_0/GATE.n470 sky130_asc_pfet_01v8_lvt_60_0/GATE.n468 85.333
R277 sky130_asc_pfet_01v8_lvt_60_0/GATE.n472 sky130_asc_pfet_01v8_lvt_60_0/GATE.n470 85.333
R278 sky130_asc_pfet_01v8_lvt_60_0/GATE.n475 sky130_asc_pfet_01v8_lvt_60_0/GATE.n472 85.333
R279 sky130_asc_pfet_01v8_lvt_60_0/GATE.n477 sky130_asc_pfet_01v8_lvt_60_0/GATE.n475 85.333
R280 sky130_asc_pfet_01v8_lvt_60_0/GATE.n480 sky130_asc_pfet_01v8_lvt_60_0/GATE.n477 85.333
R281 sky130_asc_pfet_01v8_lvt_60_0/GATE.n483 sky130_asc_pfet_01v8_lvt_60_0/GATE.n480 85.333
R282 sky130_asc_pfet_01v8_lvt_60_0/GATE.n486 sky130_asc_pfet_01v8_lvt_60_0/GATE.n483 85.333
R283 sky130_asc_pfet_01v8_lvt_60_0/GATE.n489 sky130_asc_pfet_01v8_lvt_60_0/GATE.n486 85.333
R284 sky130_asc_pfet_01v8_lvt_60_0/GATE.n502 sky130_asc_pfet_01v8_lvt_60_0/GATE.n499 85.333
R285 sky130_asc_pfet_01v8_lvt_60_0/GATE.n504 sky130_asc_pfet_01v8_lvt_60_0/GATE.n502 85.333
R286 sky130_asc_pfet_01v8_lvt_60_0/GATE.n507 sky130_asc_pfet_01v8_lvt_60_0/GATE.n504 85.333
R287 sky130_asc_pfet_01v8_lvt_60_0/GATE.n510 sky130_asc_pfet_01v8_lvt_60_0/GATE.n507 85.333
R288 sky130_asc_pfet_01v8_lvt_60_0/GATE.n513 sky130_asc_pfet_01v8_lvt_60_0/GATE.n510 85.333
R289 sky130_asc_pfet_01v8_lvt_60_0/GATE.n516 sky130_asc_pfet_01v8_lvt_60_0/GATE.n513 85.333
R290 sky130_asc_pfet_01v8_lvt_60_0/GATE.n518 sky130_asc_pfet_01v8_lvt_60_0/GATE.n516 85.333
R291 sky130_asc_pfet_01v8_lvt_60_0/GATE.n520 sky130_asc_pfet_01v8_lvt_60_0/GATE.n518 85.333
R292 sky130_asc_pfet_01v8_lvt_60_0/GATE.n523 sky130_asc_pfet_01v8_lvt_60_0/GATE.n520 85.333
R293 sky130_asc_pfet_01v8_lvt_60_0/GATE.n525 sky130_asc_pfet_01v8_lvt_60_0/GATE.n523 85.333
R294 sky130_asc_pfet_01v8_lvt_60_0/GATE.n528 sky130_asc_pfet_01v8_lvt_60_0/GATE.n525 85.333
R295 sky130_asc_pfet_01v8_lvt_60_0/GATE.n531 sky130_asc_pfet_01v8_lvt_60_0/GATE.n528 85.333
R296 sky130_asc_pfet_01v8_lvt_60_0/GATE.n534 sky130_asc_pfet_01v8_lvt_60_0/GATE.n531 85.333
R297 sky130_asc_pfet_01v8_lvt_60_0/GATE.n537 sky130_asc_pfet_01v8_lvt_60_0/GATE.n534 85.333
R298 sky130_asc_pfet_01v8_lvt_60_0/GATE.n539 sky130_asc_pfet_01v8_lvt_60_0/GATE.n537 85.333
R299 sky130_asc_pfet_01v8_lvt_60_0/GATE.n541 sky130_asc_pfet_01v8_lvt_60_0/GATE.n539 85.333
R300 sky130_asc_pfet_01v8_lvt_60_0/GATE.n544 sky130_asc_pfet_01v8_lvt_60_0/GATE.n541 85.333
R301 sky130_asc_pfet_01v8_lvt_60_0/GATE.n546 sky130_asc_pfet_01v8_lvt_60_0/GATE.n544 85.333
R302 sky130_asc_pfet_01v8_lvt_60_0/GATE.n549 sky130_asc_pfet_01v8_lvt_60_0/GATE.n546 85.333
R303 sky130_asc_pfet_01v8_lvt_60_0/GATE.n552 sky130_asc_pfet_01v8_lvt_60_0/GATE.n549 85.333
R304 sky130_asc_pfet_01v8_lvt_60_0/GATE.n555 sky130_asc_pfet_01v8_lvt_60_0/GATE.n552 85.333
R305 sky130_asc_pfet_01v8_lvt_60_0/GATE.n558 sky130_asc_pfet_01v8_lvt_60_0/GATE.n555 85.333
R306 sky130_asc_pfet_01v8_lvt_60_0/GATE.n560 sky130_asc_pfet_01v8_lvt_60_0/GATE.n558 85.333
R307 sky130_asc_pfet_01v8_lvt_60_0/GATE.n562 sky130_asc_pfet_01v8_lvt_60_0/GATE.n560 85.333
R308 sky130_asc_pfet_01v8_lvt_60_0/GATE.n565 sky130_asc_pfet_01v8_lvt_60_0/GATE.n562 85.333
R309 sky130_asc_pfet_01v8_lvt_60_0/GATE.n567 sky130_asc_pfet_01v8_lvt_60_0/GATE.n565 85.333
R310 sky130_asc_pfet_01v8_lvt_60_0/GATE.n570 sky130_asc_pfet_01v8_lvt_60_0/GATE.n567 85.333
R311 sky130_asc_pfet_01v8_lvt_60_0/GATE.n573 sky130_asc_pfet_01v8_lvt_60_0/GATE.n570 85.333
R312 sky130_asc_pfet_01v8_lvt_60_0/GATE.n576 sky130_asc_pfet_01v8_lvt_60_0/GATE.n573 85.333
R313 sky130_asc_pfet_01v8_lvt_60_0/GATE.n578 sky130_asc_pfet_01v8_lvt_60_0/GATE.n576 85.333
R314 sky130_asc_pfet_01v8_lvt_60_0/GATE.n220 sky130_asc_pfet_01v8_lvt_60_0/GATE.n217 85.333
R315 sky130_asc_pfet_01v8_lvt_60_0/GATE.n223 sky130_asc_pfet_01v8_lvt_60_0/GATE.n220 85.333
R316 sky130_asc_pfet_01v8_lvt_60_0/GATE.n226 sky130_asc_pfet_01v8_lvt_60_0/GATE.n223 85.333
R317 sky130_asc_pfet_01v8_lvt_60_0/GATE.n228 sky130_asc_pfet_01v8_lvt_60_0/GATE.n226 85.333
R318 sky130_asc_pfet_01v8_lvt_60_0/GATE.n230 sky130_asc_pfet_01v8_lvt_60_0/GATE.n228 85.333
R319 sky130_asc_pfet_01v8_lvt_60_0/GATE.n233 sky130_asc_pfet_01v8_lvt_60_0/GATE.n230 85.333
R320 sky130_asc_pfet_01v8_lvt_60_0/GATE.n235 sky130_asc_pfet_01v8_lvt_60_0/GATE.n233 85.333
R321 sky130_asc_pfet_01v8_lvt_60_0/GATE.n238 sky130_asc_pfet_01v8_lvt_60_0/GATE.n235 85.333
R322 sky130_asc_pfet_01v8_lvt_60_0/GATE.n241 sky130_asc_pfet_01v8_lvt_60_0/GATE.n238 85.333
R323 sky130_asc_pfet_01v8_lvt_60_0/GATE.n244 sky130_asc_pfet_01v8_lvt_60_0/GATE.n241 85.333
R324 sky130_asc_pfet_01v8_lvt_60_0/GATE.n247 sky130_asc_pfet_01v8_lvt_60_0/GATE.n244 85.333
R325 sky130_asc_pfet_01v8_lvt_60_0/GATE.n249 sky130_asc_pfet_01v8_lvt_60_0/GATE.n247 85.333
R326 sky130_asc_pfet_01v8_lvt_60_0/GATE.n251 sky130_asc_pfet_01v8_lvt_60_0/GATE.n249 85.333
R327 sky130_asc_pfet_01v8_lvt_60_0/GATE.n254 sky130_asc_pfet_01v8_lvt_60_0/GATE.n251 85.333
R328 sky130_asc_pfet_01v8_lvt_60_0/GATE.n256 sky130_asc_pfet_01v8_lvt_60_0/GATE.n254 85.333
R329 sky130_asc_pfet_01v8_lvt_60_0/GATE.n259 sky130_asc_pfet_01v8_lvt_60_0/GATE.n256 85.333
R330 sky130_asc_pfet_01v8_lvt_60_0/GATE.n262 sky130_asc_pfet_01v8_lvt_60_0/GATE.n259 85.333
R331 sky130_asc_pfet_01v8_lvt_60_0/GATE.n265 sky130_asc_pfet_01v8_lvt_60_0/GATE.n262 85.333
R332 sky130_asc_pfet_01v8_lvt_60_0/GATE.n268 sky130_asc_pfet_01v8_lvt_60_0/GATE.n265 85.333
R333 sky130_asc_pfet_01v8_lvt_60_0/GATE.n270 sky130_asc_pfet_01v8_lvt_60_0/GATE.n268 85.333
R334 sky130_asc_pfet_01v8_lvt_60_0/GATE.n272 sky130_asc_pfet_01v8_lvt_60_0/GATE.n270 85.333
R335 sky130_asc_pfet_01v8_lvt_60_0/GATE.n274 sky130_asc_pfet_01v8_lvt_60_0/GATE.n272 85.333
R336 sky130_asc_pfet_01v8_lvt_60_0/GATE.n276 sky130_asc_pfet_01v8_lvt_60_0/GATE.n274 85.333
R337 sky130_asc_pfet_01v8_lvt_60_0/GATE.n279 sky130_asc_pfet_01v8_lvt_60_0/GATE.n276 85.333
R338 sky130_asc_pfet_01v8_lvt_60_0/GATE.n282 sky130_asc_pfet_01v8_lvt_60_0/GATE.n279 85.333
R339 sky130_asc_pfet_01v8_lvt_60_0/GATE.n285 sky130_asc_pfet_01v8_lvt_60_0/GATE.n282 85.333
R340 sky130_asc_pfet_01v8_lvt_60_0/GATE.n288 sky130_asc_pfet_01v8_lvt_60_0/GATE.n285 85.333
R341 sky130_asc_pfet_01v8_lvt_60_0/GATE.n290 sky130_asc_pfet_01v8_lvt_60_0/GATE.n288 85.333
R342 sky130_asc_pfet_01v8_lvt_60_0/GATE.n292 sky130_asc_pfet_01v8_lvt_60_0/GATE.n290 85.333
R343 sky130_asc_pfet_01v8_lvt_60_0/GATE.n294 sky130_asc_pfet_01v8_lvt_60_0/GATE.n292 85.333
R344 sky130_asc_pfet_01v8_lvt_60_0/GATE.n297 sky130_asc_pfet_01v8_lvt_60_0/GATE.n294 85.333
R345 sky130_asc_pfet_01v8_lvt_60_0/GATE.n299 sky130_asc_pfet_01v8_lvt_60_0/GATE.n297 85.333
R346 sky130_asc_pfet_01v8_lvt_60_0/GATE.n302 sky130_asc_pfet_01v8_lvt_60_0/GATE.n299 85.333
R347 sky130_asc_pfet_01v8_lvt_60_0/GATE.n305 sky130_asc_pfet_01v8_lvt_60_0/GATE.n302 85.333
R348 sky130_asc_pfet_01v8_lvt_60_0/GATE.n308 sky130_asc_pfet_01v8_lvt_60_0/GATE.n305 85.333
R349 sky130_asc_pfet_01v8_lvt_60_0/GATE.n311 sky130_asc_pfet_01v8_lvt_60_0/GATE.n308 85.333
R350 sky130_asc_pfet_01v8_lvt_60_0/GATE.n313 sky130_asc_pfet_01v8_lvt_60_0/GATE.n311 85.333
R351 sky130_asc_pfet_01v8_lvt_60_0/GATE.n315 sky130_asc_pfet_01v8_lvt_60_0/GATE.n313 85.333
R352 sky130_asc_pfet_01v8_lvt_60_0/GATE.n318 sky130_asc_pfet_01v8_lvt_60_0/GATE.n315 85.333
R353 sky130_asc_pfet_01v8_lvt_60_0/GATE.n320 sky130_asc_pfet_01v8_lvt_60_0/GATE.n318 85.333
R354 sky130_asc_pfet_01v8_lvt_60_0/GATE.n323 sky130_asc_pfet_01v8_lvt_60_0/GATE.n320 85.333
R355 sky130_asc_pfet_01v8_lvt_60_0/GATE.n326 sky130_asc_pfet_01v8_lvt_60_0/GATE.n323 85.333
R356 sky130_asc_pfet_01v8_lvt_60_0/GATE.n329 sky130_asc_pfet_01v8_lvt_60_0/GATE.n326 85.333
R357 sky130_asc_pfet_01v8_lvt_60_0/GATE.n332 sky130_asc_pfet_01v8_lvt_60_0/GATE.n329 85.333
R358 sky130_asc_pfet_01v8_lvt_60_0/GATE.n334 sky130_asc_pfet_01v8_lvt_60_0/GATE.n332 85.333
R359 sky130_asc_pfet_01v8_lvt_60_0/GATE.n336 sky130_asc_pfet_01v8_lvt_60_0/GATE.n334 85.333
R360 sky130_asc_pfet_01v8_lvt_60_0/GATE.n339 sky130_asc_pfet_01v8_lvt_60_0/GATE.n336 85.333
R361 sky130_asc_pfet_01v8_lvt_60_0/GATE.n341 sky130_asc_pfet_01v8_lvt_60_0/GATE.n339 85.333
R362 sky130_asc_pfet_01v8_lvt_60_0/GATE.n344 sky130_asc_pfet_01v8_lvt_60_0/GATE.n341 85.333
R363 sky130_asc_pfet_01v8_lvt_60_0/GATE.n347 sky130_asc_pfet_01v8_lvt_60_0/GATE.n344 85.333
R364 sky130_asc_pfet_01v8_lvt_60_0/GATE.n350 sky130_asc_pfet_01v8_lvt_60_0/GATE.n347 85.333
R365 sky130_asc_pfet_01v8_lvt_60_0/GATE.n353 sky130_asc_pfet_01v8_lvt_60_0/GATE.n350 85.333
R366 sky130_asc_pfet_01v8_lvt_60_0/GATE.n355 sky130_asc_pfet_01v8_lvt_60_0/GATE.n353 85.333
R367 sky130_asc_pfet_01v8_lvt_60_0/GATE.n357 sky130_asc_pfet_01v8_lvt_60_0/GATE.n355 85.333
R368 sky130_asc_pfet_01v8_lvt_60_0/GATE.n360 sky130_asc_pfet_01v8_lvt_60_0/GATE.n357 85.333
R369 sky130_asc_pfet_01v8_lvt_60_0/GATE.n362 sky130_asc_pfet_01v8_lvt_60_0/GATE.n360 85.333
R370 sky130_asc_pfet_01v8_lvt_60_0/GATE.n365 sky130_asc_pfet_01v8_lvt_60_0/GATE.n362 85.333
R371 sky130_asc_pfet_01v8_lvt_60_0/GATE.n368 sky130_asc_pfet_01v8_lvt_60_0/GATE.n365 85.333
R372 sky130_asc_pfet_01v8_lvt_60_0/GATE.n371 sky130_asc_pfet_01v8_lvt_60_0/GATE.n368 85.333
R373 sky130_asc_pfet_01v8_lvt_60_0/GATE.n374 sky130_asc_pfet_01v8_lvt_60_0/GATE.n371 85.333
R374 sky130_asc_pfet_01v8_lvt_60_0/GATE.n376 sky130_asc_pfet_01v8_lvt_60_0/GATE.n374 85.333
R375 sky130_asc_pfet_01v8_lvt_60_0/GATE.n378 sky130_asc_pfet_01v8_lvt_60_0/GATE.n376 85.333
R376 sky130_asc_pfet_01v8_lvt_60_0/GATE.n381 sky130_asc_pfet_01v8_lvt_60_0/GATE.n378 85.333
R377 sky130_asc_pfet_01v8_lvt_60_0/GATE.n383 sky130_asc_pfet_01v8_lvt_60_0/GATE.n381 85.333
R378 sky130_asc_pfet_01v8_lvt_60_0/GATE.n386 sky130_asc_pfet_01v8_lvt_60_0/GATE.n383 85.333
R379 sky130_asc_pfet_01v8_lvt_60_0/GATE.n389 sky130_asc_pfet_01v8_lvt_60_0/GATE.n386 85.333
R380 sky130_asc_pfet_01v8_lvt_60_0/GATE.n392 sky130_asc_pfet_01v8_lvt_60_0/GATE.n389 85.333
R381 sky130_asc_pfet_01v8_lvt_60_0/GATE.n394 sky130_asc_pfet_01v8_lvt_60_0/GATE.n392 85.333
R382 sky130_asc_pfet_01v8_lvt_60_0/GATE.n19 sky130_asc_pfet_01v8_lvt_60_0/GATE.n16 85.333
R383 sky130_asc_pfet_01v8_lvt_60_0/GATE.n22 sky130_asc_pfet_01v8_lvt_60_0/GATE.n19 85.333
R384 sky130_asc_pfet_01v8_lvt_60_0/GATE.n25 sky130_asc_pfet_01v8_lvt_60_0/GATE.n22 85.333
R385 sky130_asc_pfet_01v8_lvt_60_0/GATE.n27 sky130_asc_pfet_01v8_lvt_60_0/GATE.n25 85.333
R386 sky130_asc_pfet_01v8_lvt_60_0/GATE.n29 sky130_asc_pfet_01v8_lvt_60_0/GATE.n27 85.333
R387 sky130_asc_pfet_01v8_lvt_60_0/GATE.n32 sky130_asc_pfet_01v8_lvt_60_0/GATE.n29 85.333
R388 sky130_asc_pfet_01v8_lvt_60_0/GATE.n34 sky130_asc_pfet_01v8_lvt_60_0/GATE.n32 85.333
R389 sky130_asc_pfet_01v8_lvt_60_0/GATE.n37 sky130_asc_pfet_01v8_lvt_60_0/GATE.n34 85.333
R390 sky130_asc_pfet_01v8_lvt_60_0/GATE.n40 sky130_asc_pfet_01v8_lvt_60_0/GATE.n37 85.333
R391 sky130_asc_pfet_01v8_lvt_60_0/GATE.n43 sky130_asc_pfet_01v8_lvt_60_0/GATE.n40 85.333
R392 sky130_asc_pfet_01v8_lvt_60_0/GATE.n46 sky130_asc_pfet_01v8_lvt_60_0/GATE.n43 85.333
R393 sky130_asc_pfet_01v8_lvt_60_0/GATE.n48 sky130_asc_pfet_01v8_lvt_60_0/GATE.n46 85.333
R394 sky130_asc_pfet_01v8_lvt_60_0/GATE.n50 sky130_asc_pfet_01v8_lvt_60_0/GATE.n48 85.333
R395 sky130_asc_pfet_01v8_lvt_60_0/GATE.n53 sky130_asc_pfet_01v8_lvt_60_0/GATE.n50 85.333
R396 sky130_asc_pfet_01v8_lvt_60_0/GATE.n55 sky130_asc_pfet_01v8_lvt_60_0/GATE.n53 85.333
R397 sky130_asc_pfet_01v8_lvt_60_0/GATE.n58 sky130_asc_pfet_01v8_lvt_60_0/GATE.n55 85.333
R398 sky130_asc_pfet_01v8_lvt_60_0/GATE.n61 sky130_asc_pfet_01v8_lvt_60_0/GATE.n58 85.333
R399 sky130_asc_pfet_01v8_lvt_60_0/GATE.n64 sky130_asc_pfet_01v8_lvt_60_0/GATE.n61 85.333
R400 sky130_asc_pfet_01v8_lvt_60_0/GATE.n67 sky130_asc_pfet_01v8_lvt_60_0/GATE.n64 85.333
R401 sky130_asc_pfet_01v8_lvt_60_0/GATE.n69 sky130_asc_pfet_01v8_lvt_60_0/GATE.n67 85.333
R402 sky130_asc_pfet_01v8_lvt_60_0/GATE.n71 sky130_asc_pfet_01v8_lvt_60_0/GATE.n69 85.333
R403 sky130_asc_pfet_01v8_lvt_60_0/GATE.n73 sky130_asc_pfet_01v8_lvt_60_0/GATE.n71 85.333
R404 sky130_asc_pfet_01v8_lvt_60_0/GATE.n75 sky130_asc_pfet_01v8_lvt_60_0/GATE.n73 85.333
R405 sky130_asc_pfet_01v8_lvt_60_0/GATE.n76 sky130_asc_pfet_01v8_lvt_60_0/GATE.n75 85.333
R406 sky130_asc_pfet_01v8_lvt_60_0/GATE.n639 sky130_asc_pfet_01v8_lvt_60_0/GATE.n76 85.333
R407 sky130_asc_pfet_01v8_lvt_60_0/GATE.n639 sky130_asc_pfet_01v8_lvt_60_0/GATE.n631 85.333
R408 sky130_asc_pfet_01v8_lvt_60_0/GATE.n631 sky130_asc_pfet_01v8_lvt_60_0/GATE.n630 85.333
R409 sky130_asc_pfet_01v8_lvt_60_0/GATE.n630 sky130_asc_pfet_01v8_lvt_60_0/GATE.n628 85.333
R410 sky130_asc_pfet_01v8_lvt_60_0/GATE.n628 sky130_asc_pfet_01v8_lvt_60_0/GATE.n627 85.333
R411 sky130_asc_pfet_01v8_lvt_60_0/GATE.n627 sky130_asc_pfet_01v8_lvt_60_0/GATE.n626 85.333
R412 sky130_asc_pfet_01v8_lvt_60_0/GATE.n626 sky130_asc_pfet_01v8_lvt_60_0/GATE.n625 85.333
R413 sky130_asc_pfet_01v8_lvt_60_0/GATE.n625 sky130_asc_pfet_01v8_lvt_60_0/GATE.n622 85.333
R414 sky130_asc_pfet_01v8_lvt_60_0/GATE.n622 sky130_asc_pfet_01v8_lvt_60_0/GATE.n619 85.333
R415 sky130_asc_pfet_01v8_lvt_60_0/GATE.n619 sky130_asc_pfet_01v8_lvt_60_0/GATE.n616 85.333
R416 sky130_asc_pfet_01v8_lvt_60_0/GATE.n616 sky130_asc_pfet_01v8_lvt_60_0/GATE.n613 85.333
R417 sky130_asc_pfet_01v8_lvt_60_0/GATE.n613 sky130_asc_pfet_01v8_lvt_60_0/GATE.n611 85.333
R418 sky130_asc_pfet_01v8_lvt_60_0/GATE.n611 sky130_asc_pfet_01v8_lvt_60_0/GATE.n608 85.333
R419 sky130_asc_pfet_01v8_lvt_60_0/GATE.n608 sky130_asc_pfet_01v8_lvt_60_0/GATE.n607 85.333
R420 sky130_asc_pfet_01v8_lvt_60_0/GATE.n607 sky130_asc_pfet_01v8_lvt_60_0/GATE.n606 85.333
R421 sky130_asc_pfet_01v8_lvt_60_0/GATE.n606 sky130_asc_pfet_01v8_lvt_60_0/GATE.n603 85.333
R422 sky130_asc_pfet_01v8_lvt_60_0/GATE.n603 sky130_asc_pfet_01v8_lvt_60_0/GATE.n600 85.333
R423 sky130_asc_pfet_01v8_lvt_60_0/GATE.n600 sky130_asc_pfet_01v8_lvt_60_0/GATE.n597 85.333
R424 sky130_asc_pfet_01v8_lvt_60_0/GATE.n597 sky130_asc_pfet_01v8_lvt_60_0/GATE.n594 85.333
R425 sky130_asc_pfet_01v8_lvt_60_0/GATE.n594 sky130_asc_pfet_01v8_lvt_60_0/GATE.n592 85.333
R426 sky130_asc_pfet_01v8_lvt_60_0/GATE.n592 sky130_asc_pfet_01v8_lvt_60_0/GATE.n589 85.333
R427 sky130_asc_pfet_01v8_lvt_60_0/GATE.n589 sky130_asc_pfet_01v8_lvt_60_0/GATE.n588 85.333
R428 sky130_asc_pfet_01v8_lvt_60_0/GATE.n588 sky130_asc_pfet_01v8_lvt_60_0/GATE.n587 85.333
R429 sky130_asc_pfet_01v8_lvt_60_0/GATE.n587 sky130_asc_pfet_01v8_lvt_60_0/GATE.n584 85.333
R430 sky130_asc_pfet_01v8_lvt_60_0/GATE.n584 sky130_asc_pfet_01v8_lvt_60_0/GATE.n216 85.333
R431 sky130_asc_pfet_01v8_lvt_60_0/GATE.n216 sky130_asc_pfet_01v8_lvt_60_0/GATE.n215 85.333
R432 sky130_asc_pfet_01v8_lvt_60_0/GATE.n215 sky130_asc_pfet_01v8_lvt_60_0/GATE.n212 85.333
R433 sky130_asc_pfet_01v8_lvt_60_0/GATE.n212 sky130_asc_pfet_01v8_lvt_60_0/GATE.n210 85.333
R434 sky130_asc_pfet_01v8_lvt_60_0/GATE.n206 sky130_asc_pfet_01v8_lvt_60_0/GATE.n205 85.333
R435 sky130_asc_pfet_01v8_lvt_60_0/GATE.n205 sky130_asc_pfet_01v8_lvt_60_0/GATE.n204 85.333
R436 sky130_asc_pfet_01v8_lvt_60_0/GATE.n204 sky130_asc_pfet_01v8_lvt_60_0/GATE.n201 85.333
R437 sky130_asc_pfet_01v8_lvt_60_0/GATE.n201 sky130_asc_pfet_01v8_lvt_60_0/GATE.n198 85.333
R438 sky130_asc_pfet_01v8_lvt_60_0/GATE.n198 sky130_asc_pfet_01v8_lvt_60_0/GATE.n195 85.333
R439 sky130_asc_pfet_01v8_lvt_60_0/GATE.n195 sky130_asc_pfet_01v8_lvt_60_0/GATE.n192 85.333
R440 sky130_asc_pfet_01v8_lvt_60_0/GATE.n192 sky130_asc_pfet_01v8_lvt_60_0/GATE.n190 85.333
R441 sky130_asc_pfet_01v8_lvt_60_0/GATE.n190 sky130_asc_pfet_01v8_lvt_60_0/GATE.n187 85.333
R442 sky130_asc_pfet_01v8_lvt_60_0/GATE.n187 sky130_asc_pfet_01v8_lvt_60_0/GATE.n186 85.333
R443 sky130_asc_pfet_01v8_lvt_60_0/GATE.n186 sky130_asc_pfet_01v8_lvt_60_0/GATE.n185 85.333
R444 sky130_asc_pfet_01v8_lvt_60_0/GATE.n185 sky130_asc_pfet_01v8_lvt_60_0/GATE.n182 85.333
R445 sky130_asc_pfet_01v8_lvt_60_0/GATE.n182 sky130_asc_pfet_01v8_lvt_60_0/GATE.n179 85.333
R446 sky130_asc_pfet_01v8_lvt_60_0/GATE.n179 sky130_asc_pfet_01v8_lvt_60_0/GATE.n176 85.333
R447 sky130_asc_pfet_01v8_lvt_60_0/GATE.n479 sky130_asc_pfet_01v8_lvt_60_0/GATE.n478 84.832
R448 sky130_asc_pfet_01v8_lvt_60_0/GATE.n301 sky130_asc_pfet_01v8_lvt_60_0/GATE.n300 84.832
R449 sky130_asc_pfet_01v8_lvt_60_0/GATE.n163 sky130_asc_pfet_01v8_lvt_60_0/GATE.n162 83.413
R450 sky130_asc_pfet_01v8_lvt_60_0/GATE.n499 sky130_asc_pfet_01v8_lvt_60_0/GATE.n497 83.413
R451 sky130_asc_pfet_01v8_lvt_60_0/GATE.n638 sky130_asc_pfet_01v8_lvt_60_0/GATE.n634 80.976
R452 sky130_asc_pfet_01v8_lvt_60_0/GATE.n638 sky130_asc_pfet_01v8_lvt_60_0/GATE.n637 80.976
R453 sky130_asc_pfet_01v8_lvt_60_0/GATE.n459 sky130_asc_pfet_01v8_lvt_60_0/GATE.n458 80.976
R454 sky130_asc_pfet_01v8_lvt_60_0/GATE.n281 sky130_asc_pfet_01v8_lvt_60_0/GATE.n280 80.976
R455 sky130_asc_pfet_01v8_lvt_60_0/GATE.n100 sky130_asc_pfet_01v8_lvt_60_0/GATE.n99 80
R456 sky130_asc_pfet_01v8_lvt_60_0/GATE.n490 sky130_asc_pfet_01v8_lvt_60_0/GATE.n489 80
R457 sky130_asc_pfet_01v8_lvt_60_0/GATE.n60 sky130_asc_pfet_01v8_lvt_60_0/GATE.n59 77.12
R458 sky130_asc_pfet_01v8_lvt_60_0/GATE.n618 sky130_asc_pfet_01v8_lvt_60_0/GATE.n617 77.12
R459 sky130_asc_pfet_01v8_lvt_60_0/GATE.n439 sky130_asc_pfet_01v8_lvt_60_0/GATE.n438 77.12
R460 sky130_asc_pfet_01v8_lvt_60_0/GATE.n261 sky130_asc_pfet_01v8_lvt_60_0/GATE.n260 77.12
R461 sky130_asc_pfet_01v8_lvt_60_0/GATE.n162 sky130_asc_pfet_01v8_lvt_60_0/GATE.n101 76
R462 sky130_asc_pfet_01v8_lvt_60_0/GATE.n161 sky130_asc_pfet_01v8_lvt_60_0/GATE.n160 76
R463 sky130_asc_pfet_01v8_lvt_60_0/GATE.n158 sky130_asc_pfet_01v8_lvt_60_0/GATE.n157 76
R464 sky130_asc_pfet_01v8_lvt_60_0/GATE.n155 sky130_asc_pfet_01v8_lvt_60_0/GATE.n154 76
R465 sky130_asc_pfet_01v8_lvt_60_0/GATE.n152 sky130_asc_pfet_01v8_lvt_60_0/GATE.n151 76
R466 sky130_asc_pfet_01v8_lvt_60_0/GATE.n149 sky130_asc_pfet_01v8_lvt_60_0/GATE.n148 76
R467 sky130_asc_pfet_01v8_lvt_60_0/GATE.n87 sky130_asc_pfet_01v8_lvt_60_0/GATE.n86 76
R468 sky130_asc_pfet_01v8_lvt_60_0/GATE.n90 sky130_asc_pfet_01v8_lvt_60_0/GATE.n89 76
R469 sky130_asc_pfet_01v8_lvt_60_0/GATE.n93 sky130_asc_pfet_01v8_lvt_60_0/GATE.n92 76
R470 sky130_asc_pfet_01v8_lvt_60_0/GATE.n96 sky130_asc_pfet_01v8_lvt_60_0/GATE.n95 76
R471 sky130_asc_pfet_01v8_lvt_60_0/GATE.n99 sky130_asc_pfet_01v8_lvt_60_0/GATE.n98 76
R472 sky130_asc_pfet_01v8_lvt_60_0/GATE.n398 sky130_asc_pfet_01v8_lvt_60_0/GATE.n397 76
R473 sky130_asc_pfet_01v8_lvt_60_0/GATE.n401 sky130_asc_pfet_01v8_lvt_60_0/GATE.n400 76
R474 sky130_asc_pfet_01v8_lvt_60_0/GATE.n404 sky130_asc_pfet_01v8_lvt_60_0/GATE.n403 76
R475 sky130_asc_pfet_01v8_lvt_60_0/GATE.n406 sky130_asc_pfet_01v8_lvt_60_0/GATE.n405 76
R476 sky130_asc_pfet_01v8_lvt_60_0/GATE.n408 sky130_asc_pfet_01v8_lvt_60_0/GATE.n407 76
R477 sky130_asc_pfet_01v8_lvt_60_0/GATE.n411 sky130_asc_pfet_01v8_lvt_60_0/GATE.n410 76
R478 sky130_asc_pfet_01v8_lvt_60_0/GATE.n413 sky130_asc_pfet_01v8_lvt_60_0/GATE.n412 76
R479 sky130_asc_pfet_01v8_lvt_60_0/GATE.n416 sky130_asc_pfet_01v8_lvt_60_0/GATE.n415 76
R480 sky130_asc_pfet_01v8_lvt_60_0/GATE.n419 sky130_asc_pfet_01v8_lvt_60_0/GATE.n418 76
R481 sky130_asc_pfet_01v8_lvt_60_0/GATE.n422 sky130_asc_pfet_01v8_lvt_60_0/GATE.n421 76
R482 sky130_asc_pfet_01v8_lvt_60_0/GATE.n425 sky130_asc_pfet_01v8_lvt_60_0/GATE.n424 76
R483 sky130_asc_pfet_01v8_lvt_60_0/GATE.n427 sky130_asc_pfet_01v8_lvt_60_0/GATE.n426 76
R484 sky130_asc_pfet_01v8_lvt_60_0/GATE.n429 sky130_asc_pfet_01v8_lvt_60_0/GATE.n428 76
R485 sky130_asc_pfet_01v8_lvt_60_0/GATE.n432 sky130_asc_pfet_01v8_lvt_60_0/GATE.n431 76
R486 sky130_asc_pfet_01v8_lvt_60_0/GATE.n434 sky130_asc_pfet_01v8_lvt_60_0/GATE.n433 76
R487 sky130_asc_pfet_01v8_lvt_60_0/GATE.n437 sky130_asc_pfet_01v8_lvt_60_0/GATE.n436 76
R488 sky130_asc_pfet_01v8_lvt_60_0/GATE.n440 sky130_asc_pfet_01v8_lvt_60_0/GATE.n439 76
R489 sky130_asc_pfet_01v8_lvt_60_0/GATE.n443 sky130_asc_pfet_01v8_lvt_60_0/GATE.n442 76
R490 sky130_asc_pfet_01v8_lvt_60_0/GATE.n446 sky130_asc_pfet_01v8_lvt_60_0/GATE.n445 76
R491 sky130_asc_pfet_01v8_lvt_60_0/GATE.n448 sky130_asc_pfet_01v8_lvt_60_0/GATE.n447 76
R492 sky130_asc_pfet_01v8_lvt_60_0/GATE.n450 sky130_asc_pfet_01v8_lvt_60_0/GATE.n449 76
R493 sky130_asc_pfet_01v8_lvt_60_0/GATE.n452 sky130_asc_pfet_01v8_lvt_60_0/GATE.n451 76
R494 sky130_asc_pfet_01v8_lvt_60_0/GATE.n454 sky130_asc_pfet_01v8_lvt_60_0/GATE.n453 76
R495 sky130_asc_pfet_01v8_lvt_60_0/GATE.n457 sky130_asc_pfet_01v8_lvt_60_0/GATE.n456 76
R496 sky130_asc_pfet_01v8_lvt_60_0/GATE.n460 sky130_asc_pfet_01v8_lvt_60_0/GATE.n459 76
R497 sky130_asc_pfet_01v8_lvt_60_0/GATE.n463 sky130_asc_pfet_01v8_lvt_60_0/GATE.n462 76
R498 sky130_asc_pfet_01v8_lvt_60_0/GATE.n466 sky130_asc_pfet_01v8_lvt_60_0/GATE.n465 76
R499 sky130_asc_pfet_01v8_lvt_60_0/GATE.n468 sky130_asc_pfet_01v8_lvt_60_0/GATE.n467 76
R500 sky130_asc_pfet_01v8_lvt_60_0/GATE.n470 sky130_asc_pfet_01v8_lvt_60_0/GATE.n469 76
R501 sky130_asc_pfet_01v8_lvt_60_0/GATE.n472 sky130_asc_pfet_01v8_lvt_60_0/GATE.n471 76
R502 sky130_asc_pfet_01v8_lvt_60_0/GATE.n475 sky130_asc_pfet_01v8_lvt_60_0/GATE.n474 76
R503 sky130_asc_pfet_01v8_lvt_60_0/GATE.n477 sky130_asc_pfet_01v8_lvt_60_0/GATE.n476 76
R504 sky130_asc_pfet_01v8_lvt_60_0/GATE.n480 sky130_asc_pfet_01v8_lvt_60_0/GATE.n479 76
R505 sky130_asc_pfet_01v8_lvt_60_0/GATE.n483 sky130_asc_pfet_01v8_lvt_60_0/GATE.n482 76
R506 sky130_asc_pfet_01v8_lvt_60_0/GATE.n486 sky130_asc_pfet_01v8_lvt_60_0/GATE.n485 76
R507 sky130_asc_pfet_01v8_lvt_60_0/GATE.n489 sky130_asc_pfet_01v8_lvt_60_0/GATE.n488 76
R508 sky130_asc_pfet_01v8_lvt_60_0/GATE.n499 sky130_asc_pfet_01v8_lvt_60_0/GATE.n498 76
R509 sky130_asc_pfet_01v8_lvt_60_0/GATE.n502 sky130_asc_pfet_01v8_lvt_60_0/GATE.n501 76
R510 sky130_asc_pfet_01v8_lvt_60_0/GATE.n504 sky130_asc_pfet_01v8_lvt_60_0/GATE.n503 76
R511 sky130_asc_pfet_01v8_lvt_60_0/GATE.n507 sky130_asc_pfet_01v8_lvt_60_0/GATE.n506 76
R512 sky130_asc_pfet_01v8_lvt_60_0/GATE.n510 sky130_asc_pfet_01v8_lvt_60_0/GATE.n509 76
R513 sky130_asc_pfet_01v8_lvt_60_0/GATE.n513 sky130_asc_pfet_01v8_lvt_60_0/GATE.n512 76
R514 sky130_asc_pfet_01v8_lvt_60_0/GATE.n516 sky130_asc_pfet_01v8_lvt_60_0/GATE.n515 76
R515 sky130_asc_pfet_01v8_lvt_60_0/GATE.n518 sky130_asc_pfet_01v8_lvt_60_0/GATE.n517 76
R516 sky130_asc_pfet_01v8_lvt_60_0/GATE.n520 sky130_asc_pfet_01v8_lvt_60_0/GATE.n519 76
R517 sky130_asc_pfet_01v8_lvt_60_0/GATE.n523 sky130_asc_pfet_01v8_lvt_60_0/GATE.n522 76
R518 sky130_asc_pfet_01v8_lvt_60_0/GATE.n525 sky130_asc_pfet_01v8_lvt_60_0/GATE.n524 76
R519 sky130_asc_pfet_01v8_lvt_60_0/GATE.n528 sky130_asc_pfet_01v8_lvt_60_0/GATE.n527 76
R520 sky130_asc_pfet_01v8_lvt_60_0/GATE.n531 sky130_asc_pfet_01v8_lvt_60_0/GATE.n530 76
R521 sky130_asc_pfet_01v8_lvt_60_0/GATE.n534 sky130_asc_pfet_01v8_lvt_60_0/GATE.n533 76
R522 sky130_asc_pfet_01v8_lvt_60_0/GATE.n537 sky130_asc_pfet_01v8_lvt_60_0/GATE.n536 76
R523 sky130_asc_pfet_01v8_lvt_60_0/GATE.n539 sky130_asc_pfet_01v8_lvt_60_0/GATE.n538 76
R524 sky130_asc_pfet_01v8_lvt_60_0/GATE.n541 sky130_asc_pfet_01v8_lvt_60_0/GATE.n540 76
R525 sky130_asc_pfet_01v8_lvt_60_0/GATE.n544 sky130_asc_pfet_01v8_lvt_60_0/GATE.n543 76
R526 sky130_asc_pfet_01v8_lvt_60_0/GATE.n546 sky130_asc_pfet_01v8_lvt_60_0/GATE.n545 76
R527 sky130_asc_pfet_01v8_lvt_60_0/GATE.n549 sky130_asc_pfet_01v8_lvt_60_0/GATE.n548 76
R528 sky130_asc_pfet_01v8_lvt_60_0/GATE.n552 sky130_asc_pfet_01v8_lvt_60_0/GATE.n551 76
R529 sky130_asc_pfet_01v8_lvt_60_0/GATE.n555 sky130_asc_pfet_01v8_lvt_60_0/GATE.n554 76
R530 sky130_asc_pfet_01v8_lvt_60_0/GATE.n558 sky130_asc_pfet_01v8_lvt_60_0/GATE.n557 76
R531 sky130_asc_pfet_01v8_lvt_60_0/GATE.n560 sky130_asc_pfet_01v8_lvt_60_0/GATE.n559 76
R532 sky130_asc_pfet_01v8_lvt_60_0/GATE.n562 sky130_asc_pfet_01v8_lvt_60_0/GATE.n561 76
R533 sky130_asc_pfet_01v8_lvt_60_0/GATE.n565 sky130_asc_pfet_01v8_lvt_60_0/GATE.n564 76
R534 sky130_asc_pfet_01v8_lvt_60_0/GATE.n567 sky130_asc_pfet_01v8_lvt_60_0/GATE.n566 76
R535 sky130_asc_pfet_01v8_lvt_60_0/GATE.n570 sky130_asc_pfet_01v8_lvt_60_0/GATE.n569 76
R536 sky130_asc_pfet_01v8_lvt_60_0/GATE.n573 sky130_asc_pfet_01v8_lvt_60_0/GATE.n572 76
R537 sky130_asc_pfet_01v8_lvt_60_0/GATE.n576 sky130_asc_pfet_01v8_lvt_60_0/GATE.n575 76
R538 sky130_asc_pfet_01v8_lvt_60_0/GATE.n228 sky130_asc_pfet_01v8_lvt_60_0/GATE.n227 76
R539 sky130_asc_pfet_01v8_lvt_60_0/GATE.n230 sky130_asc_pfet_01v8_lvt_60_0/GATE.n229 76
R540 sky130_asc_pfet_01v8_lvt_60_0/GATE.n249 sky130_asc_pfet_01v8_lvt_60_0/GATE.n248 76
R541 sky130_asc_pfet_01v8_lvt_60_0/GATE.n251 sky130_asc_pfet_01v8_lvt_60_0/GATE.n250 76
R542 sky130_asc_pfet_01v8_lvt_60_0/GATE.n270 sky130_asc_pfet_01v8_lvt_60_0/GATE.n269 76
R543 sky130_asc_pfet_01v8_lvt_60_0/GATE.n272 sky130_asc_pfet_01v8_lvt_60_0/GATE.n271 76
R544 sky130_asc_pfet_01v8_lvt_60_0/GATE.n274 sky130_asc_pfet_01v8_lvt_60_0/GATE.n273 76
R545 sky130_asc_pfet_01v8_lvt_60_0/GATE.n276 sky130_asc_pfet_01v8_lvt_60_0/GATE.n275 76
R546 sky130_asc_pfet_01v8_lvt_60_0/GATE.n290 sky130_asc_pfet_01v8_lvt_60_0/GATE.n289 76
R547 sky130_asc_pfet_01v8_lvt_60_0/GATE.n292 sky130_asc_pfet_01v8_lvt_60_0/GATE.n291 76
R548 sky130_asc_pfet_01v8_lvt_60_0/GATE.n294 sky130_asc_pfet_01v8_lvt_60_0/GATE.n293 76
R549 sky130_asc_pfet_01v8_lvt_60_0/GATE.n313 sky130_asc_pfet_01v8_lvt_60_0/GATE.n312 76
R550 sky130_asc_pfet_01v8_lvt_60_0/GATE.n315 sky130_asc_pfet_01v8_lvt_60_0/GATE.n314 76
R551 sky130_asc_pfet_01v8_lvt_60_0/GATE.n334 sky130_asc_pfet_01v8_lvt_60_0/GATE.n333 76
R552 sky130_asc_pfet_01v8_lvt_60_0/GATE.n336 sky130_asc_pfet_01v8_lvt_60_0/GATE.n335 76
R553 sky130_asc_pfet_01v8_lvt_60_0/GATE.n355 sky130_asc_pfet_01v8_lvt_60_0/GATE.n354 76
R554 sky130_asc_pfet_01v8_lvt_60_0/GATE.n357 sky130_asc_pfet_01v8_lvt_60_0/GATE.n356 76
R555 sky130_asc_pfet_01v8_lvt_60_0/GATE.n376 sky130_asc_pfet_01v8_lvt_60_0/GATE.n375 76
R556 sky130_asc_pfet_01v8_lvt_60_0/GATE.n378 sky130_asc_pfet_01v8_lvt_60_0/GATE.n377 76
R557 sky130_asc_pfet_01v8_lvt_60_0/GATE.n220 sky130_asc_pfet_01v8_lvt_60_0/GATE.n219 76
R558 sky130_asc_pfet_01v8_lvt_60_0/GATE.n223 sky130_asc_pfet_01v8_lvt_60_0/GATE.n222 76
R559 sky130_asc_pfet_01v8_lvt_60_0/GATE.n226 sky130_asc_pfet_01v8_lvt_60_0/GATE.n225 76
R560 sky130_asc_pfet_01v8_lvt_60_0/GATE.n233 sky130_asc_pfet_01v8_lvt_60_0/GATE.n232 76
R561 sky130_asc_pfet_01v8_lvt_60_0/GATE.n235 sky130_asc_pfet_01v8_lvt_60_0/GATE.n234 76
R562 sky130_asc_pfet_01v8_lvt_60_0/GATE.n238 sky130_asc_pfet_01v8_lvt_60_0/GATE.n237 76
R563 sky130_asc_pfet_01v8_lvt_60_0/GATE.n241 sky130_asc_pfet_01v8_lvt_60_0/GATE.n240 76
R564 sky130_asc_pfet_01v8_lvt_60_0/GATE.n244 sky130_asc_pfet_01v8_lvt_60_0/GATE.n243 76
R565 sky130_asc_pfet_01v8_lvt_60_0/GATE.n247 sky130_asc_pfet_01v8_lvt_60_0/GATE.n246 76
R566 sky130_asc_pfet_01v8_lvt_60_0/GATE.n254 sky130_asc_pfet_01v8_lvt_60_0/GATE.n253 76
R567 sky130_asc_pfet_01v8_lvt_60_0/GATE.n256 sky130_asc_pfet_01v8_lvt_60_0/GATE.n255 76
R568 sky130_asc_pfet_01v8_lvt_60_0/GATE.n259 sky130_asc_pfet_01v8_lvt_60_0/GATE.n258 76
R569 sky130_asc_pfet_01v8_lvt_60_0/GATE.n262 sky130_asc_pfet_01v8_lvt_60_0/GATE.n261 76
R570 sky130_asc_pfet_01v8_lvt_60_0/GATE.n265 sky130_asc_pfet_01v8_lvt_60_0/GATE.n264 76
R571 sky130_asc_pfet_01v8_lvt_60_0/GATE.n268 sky130_asc_pfet_01v8_lvt_60_0/GATE.n267 76
R572 sky130_asc_pfet_01v8_lvt_60_0/GATE.n279 sky130_asc_pfet_01v8_lvt_60_0/GATE.n278 76
R573 sky130_asc_pfet_01v8_lvt_60_0/GATE.n282 sky130_asc_pfet_01v8_lvt_60_0/GATE.n281 76
R574 sky130_asc_pfet_01v8_lvt_60_0/GATE.n285 sky130_asc_pfet_01v8_lvt_60_0/GATE.n284 76
R575 sky130_asc_pfet_01v8_lvt_60_0/GATE.n288 sky130_asc_pfet_01v8_lvt_60_0/GATE.n287 76
R576 sky130_asc_pfet_01v8_lvt_60_0/GATE.n297 sky130_asc_pfet_01v8_lvt_60_0/GATE.n296 76
R577 sky130_asc_pfet_01v8_lvt_60_0/GATE.n299 sky130_asc_pfet_01v8_lvt_60_0/GATE.n298 76
R578 sky130_asc_pfet_01v8_lvt_60_0/GATE.n302 sky130_asc_pfet_01v8_lvt_60_0/GATE.n301 76
R579 sky130_asc_pfet_01v8_lvt_60_0/GATE.n305 sky130_asc_pfet_01v8_lvt_60_0/GATE.n304 76
R580 sky130_asc_pfet_01v8_lvt_60_0/GATE.n308 sky130_asc_pfet_01v8_lvt_60_0/GATE.n307 76
R581 sky130_asc_pfet_01v8_lvt_60_0/GATE.n311 sky130_asc_pfet_01v8_lvt_60_0/GATE.n310 76
R582 sky130_asc_pfet_01v8_lvt_60_0/GATE.n318 sky130_asc_pfet_01v8_lvt_60_0/GATE.n317 76
R583 sky130_asc_pfet_01v8_lvt_60_0/GATE.n320 sky130_asc_pfet_01v8_lvt_60_0/GATE.n319 76
R584 sky130_asc_pfet_01v8_lvt_60_0/GATE.n323 sky130_asc_pfet_01v8_lvt_60_0/GATE.n322 76
R585 sky130_asc_pfet_01v8_lvt_60_0/GATE.n326 sky130_asc_pfet_01v8_lvt_60_0/GATE.n325 76
R586 sky130_asc_pfet_01v8_lvt_60_0/GATE.n329 sky130_asc_pfet_01v8_lvt_60_0/GATE.n328 76
R587 sky130_asc_pfet_01v8_lvt_60_0/GATE.n332 sky130_asc_pfet_01v8_lvt_60_0/GATE.n331 76
R588 sky130_asc_pfet_01v8_lvt_60_0/GATE.n339 sky130_asc_pfet_01v8_lvt_60_0/GATE.n338 76
R589 sky130_asc_pfet_01v8_lvt_60_0/GATE.n341 sky130_asc_pfet_01v8_lvt_60_0/GATE.n340 76
R590 sky130_asc_pfet_01v8_lvt_60_0/GATE.n344 sky130_asc_pfet_01v8_lvt_60_0/GATE.n343 76
R591 sky130_asc_pfet_01v8_lvt_60_0/GATE.n347 sky130_asc_pfet_01v8_lvt_60_0/GATE.n346 76
R592 sky130_asc_pfet_01v8_lvt_60_0/GATE.n350 sky130_asc_pfet_01v8_lvt_60_0/GATE.n349 76
R593 sky130_asc_pfet_01v8_lvt_60_0/GATE.n353 sky130_asc_pfet_01v8_lvt_60_0/GATE.n352 76
R594 sky130_asc_pfet_01v8_lvt_60_0/GATE.n360 sky130_asc_pfet_01v8_lvt_60_0/GATE.n359 76
R595 sky130_asc_pfet_01v8_lvt_60_0/GATE.n362 sky130_asc_pfet_01v8_lvt_60_0/GATE.n361 76
R596 sky130_asc_pfet_01v8_lvt_60_0/GATE.n365 sky130_asc_pfet_01v8_lvt_60_0/GATE.n364 76
R597 sky130_asc_pfet_01v8_lvt_60_0/GATE.n368 sky130_asc_pfet_01v8_lvt_60_0/GATE.n367 76
R598 sky130_asc_pfet_01v8_lvt_60_0/GATE.n371 sky130_asc_pfet_01v8_lvt_60_0/GATE.n370 76
R599 sky130_asc_pfet_01v8_lvt_60_0/GATE.n374 sky130_asc_pfet_01v8_lvt_60_0/GATE.n373 76
R600 sky130_asc_pfet_01v8_lvt_60_0/GATE.n381 sky130_asc_pfet_01v8_lvt_60_0/GATE.n380 76
R601 sky130_asc_pfet_01v8_lvt_60_0/GATE.n383 sky130_asc_pfet_01v8_lvt_60_0/GATE.n382 76
R602 sky130_asc_pfet_01v8_lvt_60_0/GATE.n386 sky130_asc_pfet_01v8_lvt_60_0/GATE.n385 76
R603 sky130_asc_pfet_01v8_lvt_60_0/GATE.n389 sky130_asc_pfet_01v8_lvt_60_0/GATE.n388 76
R604 sky130_asc_pfet_01v8_lvt_60_0/GATE.n392 sky130_asc_pfet_01v8_lvt_60_0/GATE.n391 76
R605 sky130_asc_pfet_01v8_lvt_60_0/GATE.n628 sky130_asc_pfet_01v8_lvt_60_0/GATE.n77 76
R606 sky130_asc_pfet_01v8_lvt_60_0/GATE.n627 sky130_asc_pfet_01v8_lvt_60_0/GATE.n78 76
R607 sky130_asc_pfet_01v8_lvt_60_0/GATE.n626 sky130_asc_pfet_01v8_lvt_60_0/GATE.n79 76
R608 sky130_asc_pfet_01v8_lvt_60_0/GATE.n608 sky130_asc_pfet_01v8_lvt_60_0/GATE.n80 76
R609 sky130_asc_pfet_01v8_lvt_60_0/GATE.n607 sky130_asc_pfet_01v8_lvt_60_0/GATE.n81 76
R610 sky130_asc_pfet_01v8_lvt_60_0/GATE.n589 sky130_asc_pfet_01v8_lvt_60_0/GATE.n82 76
R611 sky130_asc_pfet_01v8_lvt_60_0/GATE.n588 sky130_asc_pfet_01v8_lvt_60_0/GATE.n83 76
R612 sky130_asc_pfet_01v8_lvt_60_0/GATE.n27 sky130_asc_pfet_01v8_lvt_60_0/GATE.n26 76
R613 sky130_asc_pfet_01v8_lvt_60_0/GATE.n29 sky130_asc_pfet_01v8_lvt_60_0/GATE.n28 76
R614 sky130_asc_pfet_01v8_lvt_60_0/GATE.n48 sky130_asc_pfet_01v8_lvt_60_0/GATE.n47 76
R615 sky130_asc_pfet_01v8_lvt_60_0/GATE.n50 sky130_asc_pfet_01v8_lvt_60_0/GATE.n49 76
R616 sky130_asc_pfet_01v8_lvt_60_0/GATE.n69 sky130_asc_pfet_01v8_lvt_60_0/GATE.n68 76
R617 sky130_asc_pfet_01v8_lvt_60_0/GATE.n71 sky130_asc_pfet_01v8_lvt_60_0/GATE.n70 76
R618 sky130_asc_pfet_01v8_lvt_60_0/GATE.n73 sky130_asc_pfet_01v8_lvt_60_0/GATE.n72 76
R619 sky130_asc_pfet_01v8_lvt_60_0/GATE.n630 sky130_asc_pfet_01v8_lvt_60_0/GATE.n629 76
R620 sky130_asc_pfet_01v8_lvt_60_0/GATE.n625 sky130_asc_pfet_01v8_lvt_60_0/GATE.n624 76
R621 sky130_asc_pfet_01v8_lvt_60_0/GATE.n622 sky130_asc_pfet_01v8_lvt_60_0/GATE.n621 76
R622 sky130_asc_pfet_01v8_lvt_60_0/GATE.n619 sky130_asc_pfet_01v8_lvt_60_0/GATE.n618 76
R623 sky130_asc_pfet_01v8_lvt_60_0/GATE.n616 sky130_asc_pfet_01v8_lvt_60_0/GATE.n615 76
R624 sky130_asc_pfet_01v8_lvt_60_0/GATE.n613 sky130_asc_pfet_01v8_lvt_60_0/GATE.n612 76
R625 sky130_asc_pfet_01v8_lvt_60_0/GATE.n611 sky130_asc_pfet_01v8_lvt_60_0/GATE.n610 76
R626 sky130_asc_pfet_01v8_lvt_60_0/GATE.n606 sky130_asc_pfet_01v8_lvt_60_0/GATE.n605 76
R627 sky130_asc_pfet_01v8_lvt_60_0/GATE.n603 sky130_asc_pfet_01v8_lvt_60_0/GATE.n602 76
R628 sky130_asc_pfet_01v8_lvt_60_0/GATE.n600 sky130_asc_pfet_01v8_lvt_60_0/GATE.n599 76
R629 sky130_asc_pfet_01v8_lvt_60_0/GATE.n597 sky130_asc_pfet_01v8_lvt_60_0/GATE.n596 76
R630 sky130_asc_pfet_01v8_lvt_60_0/GATE.n594 sky130_asc_pfet_01v8_lvt_60_0/GATE.n593 76
R631 sky130_asc_pfet_01v8_lvt_60_0/GATE.n592 sky130_asc_pfet_01v8_lvt_60_0/GATE.n591 76
R632 sky130_asc_pfet_01v8_lvt_60_0/GATE.n587 sky130_asc_pfet_01v8_lvt_60_0/GATE.n586 76
R633 sky130_asc_pfet_01v8_lvt_60_0/GATE.n206 sky130_asc_pfet_01v8_lvt_60_0/GATE.n169 76
R634 sky130_asc_pfet_01v8_lvt_60_0/GATE.n205 sky130_asc_pfet_01v8_lvt_60_0/GATE.n170 76
R635 sky130_asc_pfet_01v8_lvt_60_0/GATE.n187 sky130_asc_pfet_01v8_lvt_60_0/GATE.n171 76
R636 sky130_asc_pfet_01v8_lvt_60_0/GATE.n186 sky130_asc_pfet_01v8_lvt_60_0/GATE.n172 76
R637 sky130_asc_pfet_01v8_lvt_60_0/GATE.n215 sky130_asc_pfet_01v8_lvt_60_0/GATE.n214 76
R638 sky130_asc_pfet_01v8_lvt_60_0/GATE.n212 sky130_asc_pfet_01v8_lvt_60_0/GATE.n211 76
R639 sky130_asc_pfet_01v8_lvt_60_0/GATE.n210 sky130_asc_pfet_01v8_lvt_60_0/GATE.n209 76
R640 sky130_asc_pfet_01v8_lvt_60_0/GATE.n204 sky130_asc_pfet_01v8_lvt_60_0/GATE.n203 76
R641 sky130_asc_pfet_01v8_lvt_60_0/GATE.n201 sky130_asc_pfet_01v8_lvt_60_0/GATE.n200 76
R642 sky130_asc_pfet_01v8_lvt_60_0/GATE.n198 sky130_asc_pfet_01v8_lvt_60_0/GATE.n197 76
R643 sky130_asc_pfet_01v8_lvt_60_0/GATE.n195 sky130_asc_pfet_01v8_lvt_60_0/GATE.n194 76
R644 sky130_asc_pfet_01v8_lvt_60_0/GATE.n192 sky130_asc_pfet_01v8_lvt_60_0/GATE.n191 76
R645 sky130_asc_pfet_01v8_lvt_60_0/GATE.n190 sky130_asc_pfet_01v8_lvt_60_0/GATE.n189 76
R646 sky130_asc_pfet_01v8_lvt_60_0/GATE.n185 sky130_asc_pfet_01v8_lvt_60_0/GATE.n184 76
R647 sky130_asc_pfet_01v8_lvt_60_0/GATE.n182 sky130_asc_pfet_01v8_lvt_60_0/GATE.n181 76
R648 sky130_asc_pfet_01v8_lvt_60_0/GATE.n179 sky130_asc_pfet_01v8_lvt_60_0/GATE.n178 76
R649 sky130_asc_pfet_01v8_lvt_60_0/GATE.n176 sky130_asc_pfet_01v8_lvt_60_0/GATE.n175 76
R650 sky130_asc_pfet_01v8_lvt_60_0/GATE.n19 sky130_asc_pfet_01v8_lvt_60_0/GATE.n18 76
R651 sky130_asc_pfet_01v8_lvt_60_0/GATE.n22 sky130_asc_pfet_01v8_lvt_60_0/GATE.n21 76
R652 sky130_asc_pfet_01v8_lvt_60_0/GATE.n25 sky130_asc_pfet_01v8_lvt_60_0/GATE.n24 76
R653 sky130_asc_pfet_01v8_lvt_60_0/GATE.n32 sky130_asc_pfet_01v8_lvt_60_0/GATE.n31 76
R654 sky130_asc_pfet_01v8_lvt_60_0/GATE.n34 sky130_asc_pfet_01v8_lvt_60_0/GATE.n33 76
R655 sky130_asc_pfet_01v8_lvt_60_0/GATE.n37 sky130_asc_pfet_01v8_lvt_60_0/GATE.n36 76
R656 sky130_asc_pfet_01v8_lvt_60_0/GATE.n40 sky130_asc_pfet_01v8_lvt_60_0/GATE.n39 76
R657 sky130_asc_pfet_01v8_lvt_60_0/GATE.n43 sky130_asc_pfet_01v8_lvt_60_0/GATE.n42 76
R658 sky130_asc_pfet_01v8_lvt_60_0/GATE.n46 sky130_asc_pfet_01v8_lvt_60_0/GATE.n45 76
R659 sky130_asc_pfet_01v8_lvt_60_0/GATE.n53 sky130_asc_pfet_01v8_lvt_60_0/GATE.n52 76
R660 sky130_asc_pfet_01v8_lvt_60_0/GATE.n55 sky130_asc_pfet_01v8_lvt_60_0/GATE.n54 76
R661 sky130_asc_pfet_01v8_lvt_60_0/GATE.n58 sky130_asc_pfet_01v8_lvt_60_0/GATE.n57 76
R662 sky130_asc_pfet_01v8_lvt_60_0/GATE.n61 sky130_asc_pfet_01v8_lvt_60_0/GATE.n60 76
R663 sky130_asc_pfet_01v8_lvt_60_0/GATE.n64 sky130_asc_pfet_01v8_lvt_60_0/GATE.n63 76
R664 sky130_asc_pfet_01v8_lvt_60_0/GATE.n67 sky130_asc_pfet_01v8_lvt_60_0/GATE.n66 76
R665 sky130_asc_pfet_01v8_lvt_60_0/GATE.n75 sky130_asc_pfet_01v8_lvt_60_0/GATE.n74 76
R666 sky130_asc_pfet_01v8_lvt_60_0/GATE.n207 sky130_asc_pfet_01v8_lvt_60_0/GATE.n206 73.386
R667 sky130_asc_pfet_01v8_lvt_60_0/GATE.n39 sky130_asc_pfet_01v8_lvt_60_0/GATE.n38 73.264
R668 sky130_asc_pfet_01v8_lvt_60_0/GATE.n599 sky130_asc_pfet_01v8_lvt_60_0/GATE.n598 73.264
R669 sky130_asc_pfet_01v8_lvt_60_0/GATE.n572 sky130_asc_pfet_01v8_lvt_60_0/GATE.n571 73.264
R670 sky130_asc_pfet_01v8_lvt_60_0/GATE.n418 sky130_asc_pfet_01v8_lvt_60_0/GATE.n417 73.264
R671 sky130_asc_pfet_01v8_lvt_60_0/GATE.n388 sky130_asc_pfet_01v8_lvt_60_0/GATE.n387 73.264
R672 sky130_asc_pfet_01v8_lvt_60_0/GATE.n240 sky130_asc_pfet_01v8_lvt_60_0/GATE.n239 73.264
R673 sky130_asc_pfet_01v8_lvt_60_0/GATE.n92 sky130_asc_pfet_01v8_lvt_60_0/GATE.n91 69.408
R674 sky130_asc_pfet_01v8_lvt_60_0/GATE.n581 sky130_asc_pfet_01v8_lvt_60_0/GATE.n580 69.408
R675 sky130_asc_pfet_01v8_lvt_60_0/GATE.n18 sky130_asc_pfet_01v8_lvt_60_0/GATE.n17 69.408
R676 sky130_asc_pfet_01v8_lvt_60_0/GATE.n551 sky130_asc_pfet_01v8_lvt_60_0/GATE.n550 69.408
R677 sky130_asc_pfet_01v8_lvt_60_0/GATE.n397 sky130_asc_pfet_01v8_lvt_60_0/GATE.n396 69.408
R678 sky130_asc_pfet_01v8_lvt_60_0/GATE.n367 sky130_asc_pfet_01v8_lvt_60_0/GATE.n366 69.408
R679 sky130_asc_pfet_01v8_lvt_60_0/GATE.n219 sky130_asc_pfet_01v8_lvt_60_0/GATE.n218 69.408
R680 sky130_asc_pfet_01v8_lvt_60_0/GATE.n197 sky130_asc_pfet_01v8_lvt_60_0/GATE.n196 65.552
R681 sky130_asc_pfet_01v8_lvt_60_0/GATE.n530 sky130_asc_pfet_01v8_lvt_60_0/GATE.n529 65.552
R682 sky130_asc_pfet_01v8_lvt_60_0/GATE.n346 sky130_asc_pfet_01v8_lvt_60_0/GATE.n345 65.552
R683 sky130_asc_pfet_01v8_lvt_60_0/GATE.n154 sky130_asc_pfet_01v8_lvt_60_0/GATE.n153 61.696
R684 sky130_asc_pfet_01v8_lvt_60_0/GATE.n178 sky130_asc_pfet_01v8_lvt_60_0/GATE.n177 61.696
R685 sky130_asc_pfet_01v8_lvt_60_0/GATE.n509 sky130_asc_pfet_01v8_lvt_60_0/GATE.n508 61.696
R686 sky130_asc_pfet_01v8_lvt_60_0/GATE.n325 sky130_asc_pfet_01v8_lvt_60_0/GATE.n324 61.696
R687 sky130_asc_pfet_01v8_lvt_60_0/GATE.n482 sky130_asc_pfet_01v8_lvt_60_0/GATE.n481 57.84
R688 sky130_asc_pfet_01v8_lvt_60_0/GATE.n304 sky130_asc_pfet_01v8_lvt_60_0/GATE.n303 57.84
R689 sky130_asc_pfet_01v8_lvt_60_0/GATE.n634 sky130_asc_pfet_01v8_lvt_60_0/GATE.n633 53.984
R690 sky130_asc_pfet_01v8_lvt_60_0/GATE.n637 sky130_asc_pfet_01v8_lvt_60_0/GATE.n636 53.984
R691 sky130_asc_pfet_01v8_lvt_60_0/GATE.n462 sky130_asc_pfet_01v8_lvt_60_0/GATE.n461 53.984
R692 sky130_asc_pfet_01v8_lvt_60_0/GATE.n284 sky130_asc_pfet_01v8_lvt_60_0/GATE.n283 53.984
R693 sky130_asc_pfet_01v8_lvt_60_0/GATE.n641 sky130_asc_pfet_01v8_lvt_60_0/GATE.n640 53.471
R694 sky130_asc_pfet_01v8_lvt_60_0/GATE.n644 sky130_asc_pfet_01v8_lvt_60_0/GATE.t21 52.312
R695 sky130_asc_pfet_01v8_lvt_60_0/GATE.n641 sky130_asc_pfet_01v8_lvt_60_0/GATE.t6 52.311
R696 sky130_asc_pfet_01v8_lvt_60_0/GATE.n63 sky130_asc_pfet_01v8_lvt_60_0/GATE.n62 50.128
R697 sky130_asc_pfet_01v8_lvt_60_0/GATE.n621 sky130_asc_pfet_01v8_lvt_60_0/GATE.n620 50.128
R698 sky130_asc_pfet_01v8_lvt_60_0/GATE.n442 sky130_asc_pfet_01v8_lvt_60_0/GATE.n441 50.128
R699 sky130_asc_pfet_01v8_lvt_60_0/GATE.n264 sky130_asc_pfet_01v8_lvt_60_0/GATE.n263 50.128
R700 sky130_asc_pfet_01v8_lvt_60_0/GATE.n643 sky130_asc_pfet_01v8_lvt_60_0/GATE.n5 47.884
R701 sky130_asc_pfet_01v8_lvt_60_0/GATE.n642 sky130_asc_pfet_01v8_lvt_60_0/GATE.n6 47.884
R702 sky130_asc_pfet_01v8_lvt_60_0/GATE.t75 sky130_asc_pfet_01v8_lvt_60_0/GATE.n578 47.192
R703 sky130_asc_pfet_01v8_lvt_60_0/GATE.n42 sky130_asc_pfet_01v8_lvt_60_0/GATE.n41 46.272
R704 sky130_asc_pfet_01v8_lvt_60_0/GATE.n602 sky130_asc_pfet_01v8_lvt_60_0/GATE.n601 46.272
R705 sky130_asc_pfet_01v8_lvt_60_0/GATE.n575 sky130_asc_pfet_01v8_lvt_60_0/GATE.n574 46.272
R706 sky130_asc_pfet_01v8_lvt_60_0/GATE.n421 sky130_asc_pfet_01v8_lvt_60_0/GATE.n420 46.272
R707 sky130_asc_pfet_01v8_lvt_60_0/GATE.n391 sky130_asc_pfet_01v8_lvt_60_0/GATE.n390 46.272
R708 sky130_asc_pfet_01v8_lvt_60_0/GATE.n243 sky130_asc_pfet_01v8_lvt_60_0/GATE.n242 46.272
R709 sky130_asc_pfet_01v8_lvt_60_0/GATE.n11 sky130_asc_pfet_01v8_lvt_60_0/GATE.n10 43.495
R710 sky130_asc_pfet_01v8_lvt_60_0/GATE.n12 sky130_asc_pfet_01v8_lvt_60_0/GATE.n9 43.495
R711 sky130_asc_pfet_01v8_lvt_60_0/GATE.n13 sky130_asc_pfet_01v8_lvt_60_0/GATE.n8 43.495
R712 sky130_asc_pfet_01v8_lvt_60_0/GATE.n14 sky130_asc_pfet_01v8_lvt_60_0/GATE.n7 43.495
R713 sky130_asc_pfet_01v8_lvt_60_0/GATE.n107 sky130_asc_pfet_01v8_lvt_60_0/GATE.n102 43.495
R714 sky130_asc_pfet_01v8_lvt_60_0/GATE.n106 sky130_asc_pfet_01v8_lvt_60_0/GATE.n103 43.495
R715 sky130_asc_pfet_01v8_lvt_60_0/GATE.n105 sky130_asc_pfet_01v8_lvt_60_0/GATE.n104 43.495
R716 sky130_asc_pfet_01v8_lvt_60_0/GATE.n95 sky130_asc_pfet_01v8_lvt_60_0/GATE.n94 42.416
R717 sky130_asc_pfet_01v8_lvt_60_0/GATE.n21 sky130_asc_pfet_01v8_lvt_60_0/GATE.n20 42.416
R718 sky130_asc_pfet_01v8_lvt_60_0/GATE.n583 sky130_asc_pfet_01v8_lvt_60_0/GATE.n582 42.416
R719 sky130_asc_pfet_01v8_lvt_60_0/GATE.n554 sky130_asc_pfet_01v8_lvt_60_0/GATE.n553 42.416
R720 sky130_asc_pfet_01v8_lvt_60_0/GATE.n400 sky130_asc_pfet_01v8_lvt_60_0/GATE.n399 42.416
R721 sky130_asc_pfet_01v8_lvt_60_0/GATE.n370 sky130_asc_pfet_01v8_lvt_60_0/GATE.n369 42.416
R722 sky130_asc_pfet_01v8_lvt_60_0/GATE.n222 sky130_asc_pfet_01v8_lvt_60_0/GATE.n221 42.416
R723 sky130_asc_pfet_01v8_lvt_60_0/GATE.n110 sky130_asc_pfet_01v8_lvt_60_0/GATE.n108 40.588
R724 sky130_asc_pfet_01v8_lvt_60_0/GATE.n147 sky130_asc_pfet_01v8_lvt_60_0/GATE.n4 40.368
R725 sky130_asc_pfet_01v8_lvt_60_0/GATE.n200 sky130_asc_pfet_01v8_lvt_60_0/GATE.n199 38.56
R726 sky130_asc_pfet_01v8_lvt_60_0/GATE.n533 sky130_asc_pfet_01v8_lvt_60_0/GATE.n532 38.56
R727 sky130_asc_pfet_01v8_lvt_60_0/GATE.n349 sky130_asc_pfet_01v8_lvt_60_0/GATE.n348 38.56
R728 sky130_asc_pfet_01v8_lvt_60_0/GATE.n85 sky130_asc_pfet_01v8_lvt_12_1/GATE 34.986
R729 sky130_asc_pfet_01v8_lvt_60_0/GATE.n157 sky130_asc_pfet_01v8_lvt_60_0/GATE.n156 34.704
R730 sky130_asc_pfet_01v8_lvt_60_0/GATE.n181 sky130_asc_pfet_01v8_lvt_60_0/GATE.n180 34.704
R731 sky130_asc_pfet_01v8_lvt_60_0/GATE.n512 sky130_asc_pfet_01v8_lvt_60_0/GATE.n511 34.704
R732 sky130_asc_pfet_01v8_lvt_60_0/GATE.n328 sky130_asc_pfet_01v8_lvt_60_0/GATE.n327 34.704
R733 sky130_asc_pfet_01v8_lvt_60_0/GATE.n579 sky130_asc_pfet_01v8_lvt_60_0/GATE.n394 31.596
R734 sky130_asc_pfet_01v8_lvt_60_0/GATE.n395 sky130_asc_pfet_01v8_lvt_60_0/GATE 31.573
R735 sky130_asc_pfet_01v8_lvt_60_0/GATE.n217 sky130_asc_pfet_01v8_lvt_60_1/GATE 31.573
R736 sky130_asc_pfet_01v8_lvt_60_0/GATE.n16 sky130_asc_pfet_01v8_lvt_60_2/GATE 31.573
R737 sky130_asc_pfet_01v8_lvt_60_0/GATE.n485 sky130_asc_pfet_01v8_lvt_60_0/GATE.n484 30.848
R738 sky130_asc_pfet_01v8_lvt_60_0/GATE.n307 sky130_asc_pfet_01v8_lvt_60_0/GATE.n306 30.848
R739 sky130_asc_pfet_01v8_lvt_60_0/GATE.n465 sky130_asc_pfet_01v8_lvt_60_0/GATE.n464 26.992
R740 sky130_asc_pfet_01v8_lvt_60_0/GATE.n287 sky130_asc_pfet_01v8_lvt_60_0/GATE.n286 26.992
R741 sky130_asc_pfet_01v8_lvt_60_0/GATE.n207 sky130_asc_pfet_01v8_lvt_60_0/GATE.n168 24.874
R742 sky130_asc_pfet_01v8_lvt_60_0/GATE.n66 sky130_asc_pfet_01v8_lvt_60_0/GATE.n65 23.136
R743 sky130_asc_pfet_01v8_lvt_60_0/GATE.n624 sky130_asc_pfet_01v8_lvt_60_0/GATE.n623 23.136
R744 sky130_asc_pfet_01v8_lvt_60_0/GATE.n474 sky130_asc_pfet_01v8_lvt_60_0/GATE.n473 23.136
R745 sky130_asc_pfet_01v8_lvt_60_0/GATE.n445 sky130_asc_pfet_01v8_lvt_60_0/GATE.n444 23.136
R746 sky130_asc_pfet_01v8_lvt_60_0/GATE.n296 sky130_asc_pfet_01v8_lvt_60_0/GATE.n295 23.136
R747 sky130_asc_pfet_01v8_lvt_60_0/GATE.n267 sky130_asc_pfet_01v8_lvt_60_0/GATE.n266 23.136
R748 sky130_asc_pfet_01v8_lvt_60_0/GATE.n584 sky130_asc_pfet_01v8_lvt_60_0/GATE.n579 19.816
R749 sky130_asc_pfet_01v8_lvt_60_0/GATE.n45 sky130_asc_pfet_01v8_lvt_60_0/GATE.n44 19.28
R750 sky130_asc_pfet_01v8_lvt_60_0/GATE.n605 sky130_asc_pfet_01v8_lvt_60_0/GATE.n604 19.28
R751 sky130_asc_pfet_01v8_lvt_60_0/GATE.n501 sky130_asc_pfet_01v8_lvt_60_0/GATE.n500 19.28
R752 sky130_asc_pfet_01v8_lvt_60_0/GATE.n424 sky130_asc_pfet_01v8_lvt_60_0/GATE.n423 19.28
R753 sky130_asc_pfet_01v8_lvt_60_0/GATE.n317 sky130_asc_pfet_01v8_lvt_60_0/GATE.n316 19.28
R754 sky130_asc_pfet_01v8_lvt_60_0/GATE.n246 sky130_asc_pfet_01v8_lvt_60_0/GATE.n245 19.28
R755 sky130_asc_pfet_01v8_lvt_60_0/GATE.n640 sky130_asc_pfet_01v8_lvt_60_0/GATE.n639 18.072
R756 sky130_asc_pfet_01v8_lvt_60_0/GATE.n98 sky130_asc_pfet_01v8_lvt_60_0/GATE.n97 15.424
R757 sky130_asc_pfet_01v8_lvt_60_0/GATE.n189 sky130_asc_pfet_01v8_lvt_60_0/GATE.n188 15.424
R758 sky130_asc_pfet_01v8_lvt_60_0/GATE.n24 sky130_asc_pfet_01v8_lvt_60_0/GATE.n23 15.424
R759 sky130_asc_pfet_01v8_lvt_60_0/GATE.n586 sky130_asc_pfet_01v8_lvt_60_0/GATE.n585 15.424
R760 sky130_asc_pfet_01v8_lvt_60_0/GATE.n557 sky130_asc_pfet_01v8_lvt_60_0/GATE.n556 15.424
R761 sky130_asc_pfet_01v8_lvt_60_0/GATE.n522 sky130_asc_pfet_01v8_lvt_60_0/GATE.n521 15.424
R762 sky130_asc_pfet_01v8_lvt_60_0/GATE.n403 sky130_asc_pfet_01v8_lvt_60_0/GATE.n402 15.424
R763 sky130_asc_pfet_01v8_lvt_60_0/GATE.n373 sky130_asc_pfet_01v8_lvt_60_0/GATE.n372 15.424
R764 sky130_asc_pfet_01v8_lvt_60_0/GATE.n338 sky130_asc_pfet_01v8_lvt_60_0/GATE.n337 15.424
R765 sky130_asc_pfet_01v8_lvt_60_0/GATE.n225 sky130_asc_pfet_01v8_lvt_60_0/GATE.n224 15.424
R766 sky130_asc_pfet_01v8_lvt_60_0/GATE.n210 sky130_asc_pfet_01v8_lvt_60_0/GATE.n207 11.946
R767 sky130_asc_pfet_01v8_lvt_60_0/GATE.n203 sky130_asc_pfet_01v8_lvt_60_0/GATE.n202 11.568
R768 sky130_asc_pfet_01v8_lvt_60_0/GATE.n209 sky130_asc_pfet_01v8_lvt_60_0/GATE.n208 11.568
R769 sky130_asc_pfet_01v8_lvt_60_0/GATE.n543 sky130_asc_pfet_01v8_lvt_60_0/GATE.n542 11.568
R770 sky130_asc_pfet_01v8_lvt_60_0/GATE.n536 sky130_asc_pfet_01v8_lvt_60_0/GATE.n535 11.568
R771 sky130_asc_pfet_01v8_lvt_60_0/GATE.n359 sky130_asc_pfet_01v8_lvt_60_0/GATE.n358 11.568
R772 sky130_asc_pfet_01v8_lvt_60_0/GATE.n352 sky130_asc_pfet_01v8_lvt_60_0/GATE.n351 11.568
R773 sky130_asc_pfet_01v8_lvt_60_0/GATE.n4 sky130_asc_pfet_01v8_lvt_60_0/GATE.n142 9.3
R774 sky130_asc_pfet_01v8_lvt_60_0/GATE.n3 sky130_asc_pfet_01v8_lvt_60_0/GATE.n138 9.3
R775 sky130_asc_pfet_01v8_lvt_60_0/GATE.n2 sky130_asc_pfet_01v8_lvt_60_0/GATE.n134 9.3
R776 sky130_asc_pfet_01v8_lvt_60_0/GATE.n2 sky130_asc_pfet_01v8_lvt_60_0/GATE.n130 9.3
R777 sky130_asc_pfet_01v8_lvt_60_0/GATE.n0 sky130_asc_pfet_01v8_lvt_60_0/GATE.n124 9.3
R778 sky130_asc_pfet_01v8_lvt_60_0/GATE.n0 sky130_asc_pfet_01v8_lvt_60_0/GATE.n120 9.3
R779 sky130_asc_pfet_01v8_lvt_60_0/GATE.n0 sky130_asc_pfet_01v8_lvt_60_0/GATE.n116 9.3
R780 sky130_asc_pfet_01v8_lvt_60_0/GATE.n1 sky130_asc_pfet_01v8_lvt_60_0/GATE.n112 9.3
R781 sky130_asc_pfet_01v8_lvt_60_0/GATE.n1 sky130_asc_pfet_01v8_lvt_60_0/GATE.n111 9.3
R782 sky130_asc_pfet_01v8_lvt_60_0/GATE.n1 sky130_asc_pfet_01v8_lvt_60_0/GATE.n114 9.3
R783 sky130_asc_pfet_01v8_lvt_60_0/GATE.n0 sky130_asc_pfet_01v8_lvt_60_0/GATE.n115 9.3
R784 sky130_asc_pfet_01v8_lvt_60_0/GATE.n0 sky130_asc_pfet_01v8_lvt_60_0/GATE.n118 9.3
R785 sky130_asc_pfet_01v8_lvt_60_0/GATE.n0 sky130_asc_pfet_01v8_lvt_60_0/GATE.n119 9.3
R786 sky130_asc_pfet_01v8_lvt_60_0/GATE.n0 sky130_asc_pfet_01v8_lvt_60_0/GATE.n122 9.3
R787 sky130_asc_pfet_01v8_lvt_60_0/GATE.n0 sky130_asc_pfet_01v8_lvt_60_0/GATE.n123 9.3
R788 sky130_asc_pfet_01v8_lvt_60_0/GATE.n0 sky130_asc_pfet_01v8_lvt_60_0/GATE.n126 9.3
R789 sky130_asc_pfet_01v8_lvt_60_0/GATE.n2 sky130_asc_pfet_01v8_lvt_60_0/GATE.n129 9.3
R790 sky130_asc_pfet_01v8_lvt_60_0/GATE.n2 sky130_asc_pfet_01v8_lvt_60_0/GATE.n131 9.3
R791 sky130_asc_pfet_01v8_lvt_60_0/GATE.n2 sky130_asc_pfet_01v8_lvt_60_0/GATE.n133 9.3
R792 sky130_asc_pfet_01v8_lvt_60_0/GATE.n2 sky130_asc_pfet_01v8_lvt_60_0/GATE.n135 9.3
R793 sky130_asc_pfet_01v8_lvt_60_0/GATE.n3 sky130_asc_pfet_01v8_lvt_60_0/GATE.n137 9.3
R794 sky130_asc_pfet_01v8_lvt_60_0/GATE.n3 sky130_asc_pfet_01v8_lvt_60_0/GATE.n139 9.3
R795 sky130_asc_pfet_01v8_lvt_60_0/GATE.n4 sky130_asc_pfet_01v8_lvt_60_0/GATE.n141 9.3
R796 sky130_asc_pfet_01v8_lvt_60_0/GATE.n4 sky130_asc_pfet_01v8_lvt_60_0/GATE.n143 9.3
R797 sky130_asc_pfet_01v8_lvt_60_0/GATE.n167 sky130_asc_pfet_01v8_lvt_60_0/GATE.n166 9.3
R798 sky130_asc_pfet_01v8_lvt_60_0/GATE.n495 sky130_asc_pfet_01v8_lvt_60_0/GATE.n494 9.3
R799 sky130_asc_pfet_01v8_lvt_60_0/GATE.n584 sky130_asc_pfet_01v8_lvt_60_0/GATE.n583 8.286
R800 sky130_asc_pfet_01v8_lvt_60_0/GATE.n639 sky130_asc_pfet_01v8_lvt_60_0/GATE.n638 8.286
R801 sky130_asc_pfet_01v8_lvt_60_0/GATE.n145 sky130_asc_pfet_01v8_lvt_60_0/GATE.n144 8.043
R802 sky130_asc_pfet_01v8_lvt_60_0/GATE.n160 sky130_asc_pfet_01v8_lvt_60_0/GATE.n159 7.712
R803 sky130_asc_pfet_01v8_lvt_60_0/GATE.n184 sky130_asc_pfet_01v8_lvt_60_0/GATE.n183 7.712
R804 sky130_asc_pfet_01v8_lvt_60_0/GATE.n31 sky130_asc_pfet_01v8_lvt_60_0/GATE.n30 7.712
R805 sky130_asc_pfet_01v8_lvt_60_0/GATE.n591 sky130_asc_pfet_01v8_lvt_60_0/GATE.n590 7.712
R806 sky130_asc_pfet_01v8_lvt_60_0/GATE.n564 sky130_asc_pfet_01v8_lvt_60_0/GATE.n563 7.712
R807 sky130_asc_pfet_01v8_lvt_60_0/GATE.n515 sky130_asc_pfet_01v8_lvt_60_0/GATE.n514 7.712
R808 sky130_asc_pfet_01v8_lvt_60_0/GATE.n410 sky130_asc_pfet_01v8_lvt_60_0/GATE.n409 7.712
R809 sky130_asc_pfet_01v8_lvt_60_0/GATE.n380 sky130_asc_pfet_01v8_lvt_60_0/GATE.n379 7.712
R810 sky130_asc_pfet_01v8_lvt_60_0/GATE.n331 sky130_asc_pfet_01v8_lvt_60_0/GATE.n330 7.712
R811 sky130_asc_pfet_01v8_lvt_60_0/GATE.n232 sky130_asc_pfet_01v8_lvt_60_0/GATE.n231 7.712
R812 sky130_asc_pfet_01v8_lvt_60_0/GATE.n491 sky130_asc_pfet_01v8_lvt_60_0/GATE.t181 9.123
R813 sky130_asc_pfet_01v8_lvt_60_0/GATE.n128 sky130_asc_pfet_01v8_lvt_60_0/GATE.n127 5.341
R814 sky130_asc_pfet_01v8_lvt_60_0/GATE.n0 sky130_asc_pfet_01v8_lvt_60_0/GATE.n128 4.65
R815 sky130_asc_pfet_01v8_lvt_60_0/GATE.n5 sky130_asc_pfet_01v8_lvt_60_0/GATE.t20 4.428
R816 sky130_asc_pfet_01v8_lvt_60_0/GATE.n5 sky130_asc_pfet_01v8_lvt_60_0/GATE.t19 4.428
R817 sky130_asc_pfet_01v8_lvt_60_0/GATE.n6 sky130_asc_pfet_01v8_lvt_60_0/GATE.t18 4.428
R818 sky130_asc_pfet_01v8_lvt_60_0/GATE.n6 sky130_asc_pfet_01v8_lvt_60_0/GATE.t7 4.428
R819 sky130_asc_pfet_01v8_lvt_60_0/GATE.n10 sky130_asc_pfet_01v8_lvt_60_0/GATE.t17 4.35
R820 sky130_asc_pfet_01v8_lvt_60_0/GATE.n10 sky130_asc_pfet_01v8_lvt_60_0/GATE.t12 4.35
R821 sky130_asc_pfet_01v8_lvt_60_0/GATE.n9 sky130_asc_pfet_01v8_lvt_60_0/GATE.t9 4.35
R822 sky130_asc_pfet_01v8_lvt_60_0/GATE.n9 sky130_asc_pfet_01v8_lvt_60_0/GATE.t14 4.35
R823 sky130_asc_pfet_01v8_lvt_60_0/GATE.n8 sky130_asc_pfet_01v8_lvt_60_0/GATE.t10 4.35
R824 sky130_asc_pfet_01v8_lvt_60_0/GATE.n8 sky130_asc_pfet_01v8_lvt_60_0/GATE.t13 4.35
R825 sky130_asc_pfet_01v8_lvt_60_0/GATE.n7 sky130_asc_pfet_01v8_lvt_60_0/GATE.t11 4.35
R826 sky130_asc_pfet_01v8_lvt_60_0/GATE.n7 sky130_asc_pfet_01v8_lvt_60_0/GATE.t15 4.35
R827 sky130_asc_pfet_01v8_lvt_60_0/GATE.n144 sky130_asc_pfet_01v8_lvt_60_0/GATE.t0 4.35
R828 sky130_asc_pfet_01v8_lvt_60_0/GATE.n144 sky130_asc_pfet_01v8_lvt_60_0/GATE.t22 4.35
R829 sky130_asc_pfet_01v8_lvt_60_0/GATE.n102 sky130_asc_pfet_01v8_lvt_60_0/GATE.t8 4.35
R830 sky130_asc_pfet_01v8_lvt_60_0/GATE.n102 sky130_asc_pfet_01v8_lvt_60_0/GATE.t23 4.35
R831 sky130_asc_pfet_01v8_lvt_60_0/GATE.n103 sky130_asc_pfet_01v8_lvt_60_0/GATE.t1 4.35
R832 sky130_asc_pfet_01v8_lvt_60_0/GATE.n103 sky130_asc_pfet_01v8_lvt_60_0/GATE.t3 4.35
R833 sky130_asc_pfet_01v8_lvt_60_0/GATE.n104 sky130_asc_pfet_01v8_lvt_60_0/GATE.t4 4.35
R834 sky130_asc_pfet_01v8_lvt_60_0/GATE.n104 sky130_asc_pfet_01v8_lvt_60_0/GATE.t2 4.35
R835 sky130_asc_pfet_01v8_lvt_60_0/GATE.n52 sky130_asc_pfet_01v8_lvt_60_0/GATE.n51 3.856
R836 sky130_asc_pfet_01v8_lvt_60_0/GATE.n610 sky130_asc_pfet_01v8_lvt_60_0/GATE.n609 3.856
R837 sky130_asc_pfet_01v8_lvt_60_0/GATE.n488 sky130_asc_pfet_01v8_lvt_60_0/GATE.n487 3.856
R838 sky130_asc_pfet_01v8_lvt_60_0/GATE.n431 sky130_asc_pfet_01v8_lvt_60_0/GATE.n430 3.856
R839 sky130_asc_pfet_01v8_lvt_60_0/GATE.n310 sky130_asc_pfet_01v8_lvt_60_0/GATE.n309 3.856
R840 sky130_asc_pfet_01v8_lvt_60_0/GATE.n253 sky130_asc_pfet_01v8_lvt_60_0/GATE.n252 3.856
R841 sky130_asc_pfet_01v8_lvt_60_0/GATE.n640 sky130_asc_pfet_01v8_lvt_60_0/GATE.n15 3.772
R842 sky130_asc_pfet_01v8_lvt_60_0/GATE.n4 sky130_asc_pfet_01v8_lvt_60_0/GATE.n145 3.033
R843 sky130_asc_pfet_01v8_lvt_60_0/GATE.n579 sky130_asc_pfet_01v8_lvt_60_0/GATE.t155 2.914
R844 sky130_asc_pfet_01v8_lvt_60_0/GATE.n110 sky130_asc_pfet_01v8_lvt_60_0/GATE.n109 2.885
R845 sky130_asc_pfet_01v8_lvt_60_0/GATE.n493 sky130_asc_pfet_01v8_lvt_60_0/GATE.n492 2.567
R846 sky130_asc_pfet_01v8_lvt_60_0/GATE.n1 sky130_asc_pfet_01v8_lvt_60_0/GATE.n110 2.249
R847 sky130_asc_pfet_01v8_lvt_60_0/GATE.t155 sky130_asc_cap_mim_m3_1_3/Cout 1.994
R848 sky130_asc_cap_mim_m3_1_3/Cout sky130_asc_pfet_01v8_lvt_60_0/GATE.t75 1.962
R849 sky130_asc_pfet_01v8_lvt_60_0/GATE.n168 sky130_asc_pfet_01v8_lvt_60_0/GATE.n100 1.92
R850 sky130_asc_pfet_01v8_lvt_60_0/GATE.n164 sky130_asc_pfet_01v8_lvt_60_0/GATE.n163 1.92
R851 sky130_asc_pfet_01v8_lvt_60_0/GATE.n491 sky130_asc_pfet_01v8_lvt_60_0/GATE.n490 1.92
R852 sky130_asc_pfet_01v8_lvt_60_0/GATE.n497 sky130_asc_pfet_01v8_lvt_60_0/GATE.n496 1.92
R853 sky130_asc_pfet_01v8_lvt_60_0/GATE.n168 sky130_asc_pfet_01v8_lvt_60_0/GATE.n167 1.706
R854 sky130_asc_pfet_01v8_lvt_60_0/GATE.n167 sky130_asc_pfet_01v8_lvt_60_0/GATE.n164 1.706
R855 sky130_asc_pfet_01v8_lvt_60_0/GATE.n495 sky130_asc_pfet_01v8_lvt_60_0/GATE.n491 1.706
R856 sky130_asc_pfet_01v8_lvt_60_0/GATE.n496 sky130_asc_pfet_01v8_lvt_60_0/GATE.n495 1.706
R857 sky130_asc_pfet_01v8_lvt_60_0/GATE.n494 sky130_asc_pfet_01v8_lvt_60_0/GATE.n493 1.606
R858 sky130_asc_pfet_01v8_lvt_6_0/DRAIN sky130_asc_pfet_01v8_lvt_60_0/GATE.n644 0.853
R859 sky130_asc_pfet_01v8_lvt_60_0/GATE.n166 sky130_asc_pfet_01v8_lvt_60_0/GATE.n165 0.803
R860 sky130_asc_pfet_01v8_lvt_60_0/GATE.n0 sky130_asc_pfet_01v8_lvt_60_0/GATE.n1 0.612
R861 sky130_asc_cap_mim_m3_1_3/Cout sky130_asc_pfet_01v8_lvt_60_0/GATE.t46 0.525
R862 sky130_asc_pfet_01v8_lvt_60_0/GATE.t155 sky130_asc_pfet_01v8_lvt_60_0/GATE.t81 0.516
R863 sky130_asc_pfet_01v8_lvt_60_0/GATE.t181 sky130_asc_pfet_01v8_lvt_60_0/GATE.t40 0.516
R864 sky130_asc_pfet_01v8_lvt_60_0/GATE.n141 sky130_asc_pfet_01v8_lvt_60_0/GATE.n140 0.414
R865 sky130_asc_pfet_01v8_lvt_60_0/GATE.n114 sky130_asc_pfet_01v8_lvt_60_0/GATE.n113 0.414
R866 sky130_asc_pfet_01v8_lvt_60_0/GATE.t162 sky130_asc_pfet_01v8_lvt_60_0/GATE.t38 0.392
R867 sky130_asc_pfet_01v8_lvt_60_0/GATE.t44 sky130_asc_pfet_01v8_lvt_60_0/GATE.t162 0.392
R868 sky130_asc_pfet_01v8_lvt_60_0/GATE.t81 sky130_asc_pfet_01v8_lvt_60_0/GATE.t44 0.392
R869 sky130_asc_pfet_01v8_lvt_60_0/GATE.t109 sky130_asc_pfet_01v8_lvt_60_0/GATE.t54 0.392
R870 sky130_asc_pfet_01v8_lvt_60_0/GATE.t50 sky130_asc_pfet_01v8_lvt_60_0/GATE.t109 0.392
R871 sky130_asc_pfet_01v8_lvt_60_0/GATE.t26 sky130_asc_pfet_01v8_lvt_60_0/GATE.t50 0.392
R872 sky130_asc_pfet_01v8_lvt_60_0/GATE.t46 sky130_asc_pfet_01v8_lvt_60_0/GATE.t26 0.392
R873 sky130_asc_pfet_01v8_lvt_60_0/GATE.t55 sky130_asc_pfet_01v8_lvt_60_0/GATE.t106 0.392
R874 sky130_asc_pfet_01v8_lvt_60_0/GATE.t73 sky130_asc_pfet_01v8_lvt_60_0/GATE.t55 0.392
R875 sky130_asc_pfet_01v8_lvt_60_0/GATE.t89 sky130_asc_pfet_01v8_lvt_60_0/GATE.t73 0.392
R876 sky130_asc_cap_mim_m3_1_3/Cout sky130_asc_pfet_01v8_lvt_60_0/GATE.t89 0.392
R877 sky130_asc_pfet_01v8_lvt_60_0/GATE.t34 sky130_asc_pfet_01v8_lvt_60_0/GATE.t97 0.392
R878 sky130_asc_pfet_01v8_lvt_60_0/GATE.t43 sky130_asc_pfet_01v8_lvt_60_0/GATE.t34 0.392
R879 sky130_asc_pfet_01v8_lvt_60_0/GATE.t40 sky130_asc_pfet_01v8_lvt_60_0/GATE.t43 0.392
R880 sky130_asc_pfet_01v8_lvt_60_0/GATE.t93 sky130_asc_pfet_01v8_lvt_60_0/GATE.t33 0.392
R881 sky130_asc_pfet_01v8_lvt_60_0/GATE.t27 sky130_asc_pfet_01v8_lvt_60_0/GATE.t93 0.392
R882 sky130_asc_pfet_01v8_lvt_60_0/GATE.t157 sky130_asc_pfet_01v8_lvt_60_0/GATE.t27 0.392
R883 sky130_asc_pfet_01v8_lvt_60_0/GATE.n137 sky130_asc_pfet_01v8_lvt_60_0/GATE.n136 0.382
R884 sky130_asc_pfet_01v8_lvt_60_0/GATE.n118 sky130_asc_pfet_01v8_lvt_60_0/GATE.n117 0.382
R885 sky130_asc_pfet_01v8_lvt_60_0/GATE.n2 sky130_asc_pfet_01v8_lvt_60_0/GATE.n0 0.38
R886 sky130_asc_pfet_01v8_lvt_60_0/GATE.n3 sky130_asc_pfet_01v8_lvt_60_0/GATE.n2 0.378
R887 sky130_asc_pfet_01v8_lvt_60_0/GATE.t75 sky130_asc_pfet_01v8_lvt_60_0/GATE.t157 0.372
R888 sky130_asc_pfet_01v8_lvt_60_0/GATE.n133 sky130_asc_pfet_01v8_lvt_60_0/GATE.n132 0.35
R889 sky130_asc_pfet_01v8_lvt_60_0/GATE.n122 sky130_asc_pfet_01v8_lvt_60_0/GATE.n121 0.35
R890 sky130_asc_pfet_01v8_lvt_60_0/GATE.n4 sky130_asc_pfet_01v8_lvt_60_0/GATE.n3 0.33
R891 sky130_asc_pfet_01v8_lvt_60_0/GATE.t106 sky130_asc_pfet_01v8_lvt_60_0/GATE.t92 0.32
R892 sky130_asc_pfet_01v8_lvt_60_0/GATE.t38 sky130_asc_pfet_01v8_lvt_60_0/GATE.t51 0.32
R893 sky130_asc_pfet_01v8_lvt_60_0/GATE.t54 sky130_asc_pfet_01v8_lvt_60_0/GATE.t72 0.32
R894 sky130_asc_pfet_01v8_lvt_60_0/GATE.t97 sky130_asc_pfet_01v8_lvt_60_0/GATE.t36 0.32
R895 sky130_asc_pfet_01v8_lvt_60_0/GATE.t33 sky130_asc_pfet_01v8_lvt_60_0/GATE.t130 0.32
R896 sky130_asc_pfet_01v8_lvt_60_0/GATE.n126 sky130_asc_pfet_01v8_lvt_60_0/GATE.n125 0.317
R897 VDD.n725 VDD.t440 6271.13
R898 VDD.n560 VDD.t416 6271.13
R899 VDD.n725 sky130_asc_pfet_01v8_lvt_6_0/VPWR 1077.32
R900 VDD.n1 sky130_asc_pfet_01v8_lvt_12_0/VPWR 1077.32
R901 VDD.n560 sky130_asc_pfet_01v8_lvt_12_1/VPWR 1077.32
R902 VDD.n4 sky130_asc_pfet_01v8_lvt_60_2/VPWR 1077.32
R903 VDD.n513 sky130_asc_pfet_01v8_lvt_6_1/VPWR 1077.32
R904 VDD.n81 sky130_asc_pfet_01v8_lvt_60_1/VPWR 1077.32
R905 VDD.n991 VDD 1077.32
R906 VDD.n720 VDD.n719 325.944
R907 VDD.n333 VDD.n332 325.944
R908 VDD.n283 VDD.n282 325.944
R909 VDD.n976 VDD.n975 325.944
R910 VDD.n572 VDD.n570 324.987
R911 VDD.n72 VDD.n70 324.921
R912 VDD.n625 VDD.n624 293.12
R913 VDD.n626 VDD.n625 293.12
R914 VDD.n627 VDD.n626 293.12
R915 VDD.n628 VDD.n627 293.12
R916 VDD.n567 VDD.n566 293.12
R917 VDD.n568 VDD.n567 293.12
R918 VDD.n569 VDD.n568 293.12
R919 VDD.n570 VDD.n569 293.12
R920 VDD.n305 VDD.n304 293.12
R921 VDD.n306 VDD.n305 293.12
R922 VDD.n307 VDD.n306 293.12
R923 VDD.n308 VDD.n307 293.12
R924 VDD.n309 VDD.n308 293.12
R925 VDD.n310 VDD.n309 293.12
R926 VDD.n311 VDD.n310 293.12
R927 VDD.n312 VDD.n311 293.12
R928 VDD.n313 VDD.n312 293.12
R929 VDD.n314 VDD.n313 293.12
R930 VDD.n315 VDD.n314 293.12
R931 VDD.n316 VDD.n315 293.12
R932 VDD.n317 VDD.n316 293.12
R933 VDD.n318 VDD.n317 293.12
R934 VDD.n319 VDD.n318 293.12
R935 VDD.n320 VDD.n319 293.12
R936 VDD.n344 VDD.n320 293.12
R937 VDD.n344 VDD.n343 293.12
R938 VDD.n343 VDD.n342 293.12
R939 VDD.n342 VDD.n341 293.12
R940 VDD.n341 VDD.n340 293.12
R941 VDD.n340 VDD.n339 293.12
R942 VDD.n339 VDD.n338 293.12
R943 VDD.n338 VDD.n337 293.12
R944 VDD.n337 VDD.n336 293.12
R945 VDD.n336 VDD.n335 293.12
R946 VDD.n335 VDD.n334 293.12
R947 VDD.n334 VDD.n333 293.12
R948 VDD.n283 VDD.n281 293.12
R949 VDD.n43 VDD.n42 293.12
R950 VDD.n44 VDD.n43 293.12
R951 VDD.n45 VDD.n44 293.12
R952 VDD.n46 VDD.n45 293.12
R953 VDD.n47 VDD.n46 293.12
R954 VDD.n48 VDD.n47 293.12
R955 VDD.n49 VDD.n48 293.12
R956 VDD.n50 VDD.n49 293.12
R957 VDD.n51 VDD.n50 293.12
R958 VDD.n52 VDD.n51 293.12
R959 VDD.n53 VDD.n52 293.12
R960 VDD.n54 VDD.n53 293.12
R961 VDD.n55 VDD.n54 293.12
R962 VDD.n56 VDD.n55 293.12
R963 VDD.n57 VDD.n56 293.12
R964 VDD.n58 VDD.n57 293.12
R965 VDD.n59 VDD.n58 293.12
R966 VDD.n60 VDD.n59 293.12
R967 VDD.n61 VDD.n60 293.12
R968 VDD.n62 VDD.n61 293.12
R969 VDD.n63 VDD.n62 293.12
R970 VDD.n64 VDD.n63 293.12
R971 VDD.n65 VDD.n64 293.12
R972 VDD.n66 VDD.n65 293.12
R973 VDD.n67 VDD.n66 293.12
R974 VDD.n68 VDD.n67 293.12
R975 VDD.n69 VDD.n68 293.12
R976 VDD.n70 VDD.n69 293.12
R977 VDD.n948 VDD.n947 293.12
R978 VDD.n949 VDD.n948 293.12
R979 VDD.n950 VDD.n949 293.12
R980 VDD.n951 VDD.n950 293.12
R981 VDD.n952 VDD.n951 293.12
R982 VDD.n953 VDD.n952 293.12
R983 VDD.n954 VDD.n953 293.12
R984 VDD.n955 VDD.n954 293.12
R985 VDD.n956 VDD.n955 293.12
R986 VDD.n957 VDD.n956 293.12
R987 VDD.n958 VDD.n957 293.12
R988 VDD.n959 VDD.n958 293.12
R989 VDD.n960 VDD.n959 293.12
R990 VDD.n961 VDD.n960 293.12
R991 VDD.n962 VDD.n961 293.12
R992 VDD.n963 VDD.n962 293.12
R993 VDD.n964 VDD.n963 293.12
R994 VDD.n986 VDD.n964 293.12
R995 VDD.n986 VDD.n985 293.12
R996 VDD.n985 VDD.n984 293.12
R997 VDD.n984 VDD.n983 293.12
R998 VDD.n983 VDD.n982 293.12
R999 VDD.n982 VDD.n981 293.12
R1000 VDD.n981 VDD.n980 293.12
R1001 VDD.n980 VDD.n979 293.12
R1002 VDD.n979 VDD.n978 293.12
R1003 VDD.n978 VDD.n977 293.12
R1004 VDD.n977 VDD.n976 293.12
R1005 VDD.t488 VDD.t490 264.177
R1006 VDD.t484 VDD.t488 264.177
R1007 VDD.t482 VDD.t484 264.177
R1008 VDD.t440 VDD.t442 264.177
R1009 VDD.t477 VDD.t459 264.177
R1010 VDD.t480 VDD.t477 264.177
R1011 VDD.t447 VDD.t480 264.177
R1012 VDD.t450 VDD.t456 264.177
R1013 VDD.t465 VDD.t462 264.177
R1014 VDD.t471 VDD.t474 264.177
R1015 VDD.t430 VDD.t134 264.177
R1016 VDD.t434 VDD.t430 264.177
R1017 VDD.t79 VDD.t434 264.177
R1018 VDD.t96 VDD.t34 264.177
R1019 VDD.t386 VDD.t96 264.177
R1020 VDD.t346 VDD.t412 264.177
R1021 VDD.t422 VDD.t346 264.177
R1022 VDD.t416 VDD.t59 264.177
R1023 VDD.t274 VDD.t122 264.177
R1024 VDD.t168 VDD.t274 264.177
R1025 VDD.t172 VDD.t168 264.177
R1026 VDD.t238 VDD.t30 264.177
R1027 VDD.t232 VDD.t317 264.177
R1028 VDD.t248 VDD.t296 264.177
R1029 VDD.t190 VDD.t132 264.177
R1030 VDD.t207 VDD.t75 264.177
R1031 VDD.t178 VDD.t174 264.177
R1032 VDD.t64 VDD.t54 264.177
R1033 VDD.t188 VDD.t240 264.177
R1034 VDD.t46 VDD.t114 264.177
R1035 VDD.t203 VDD.t163 264.177
R1036 VDD.t376 VDD.t89 264.177
R1037 VDD.t396 VDD.t103 264.177
R1038 VDD.t42 VDD.t364 264.177
R1039 VDD.t400 VDD.t332 264.177
R1040 VDD.t402 VDD.t404 264.177
R1041 VDD.t378 VDD.t6 264.177
R1042 VDD.t380 VDD.t313 264.177
R1043 VDD.t2 VDD.t486 264.177
R1044 VDD.t444 VDD.t2 264.177
R1045 VDD.t492 VDD.t444 264.177
R1046 VDD.t4 VDD.t0 264.177
R1047 VDD.t250 VDD.t366 264.177
R1048 VDD.t300 VDD.t250 264.177
R1049 VDD.t424 VDD.t300 264.177
R1050 VDD.t370 VDD.t432 264.177
R1051 VDD.t410 VDD.t408 264.177
R1052 VDD.t352 VDD.t280 264.177
R1053 VDD.t392 VDD.t290 264.177
R1054 VDD.t244 VDD.t336 264.177
R1055 VDD.t128 VDD.t307 264.177
R1056 VDD.t372 VDD.t338 264.177
R1057 VDD.t388 VDD.t321 264.177
R1058 VDD.t26 VDD.t286 264.177
R1059 VDD.t294 VDD.t298 264.177
R1060 VDD.t209 VDD.t217 264.177
R1061 VDD.t159 VDD.t138 264.177
R1062 VDD.t52 VDD.t276 264.177
R1063 VDD.t284 VDD.t328 264.177
R1064 VDD.t242 VDD.t28 264.177
R1065 VDD.t205 VDD.t118 264.177
R1066 VDD.t211 VDD.t221 264.177
R1067 VDD.t268 VDD.t266 264.177
R1068 VDD.t136 VDD.t268 264.177
R1069 VDD.t278 VDD.t136 264.177
R1070 VDD.t382 VDD.t341 264.177
R1071 VDD.t323 VDD.t390 264.177
R1072 VDD.t236 VDD.t368 264.177
R1073 VDD.t302 VDD.t116 264.177
R1074 VDD.t157 VDD.t219 264.177
R1075 VDD.t99 VDD.t165 264.177
R1076 VDD.t61 VDD.t186 264.177
R1077 VDD.t292 VDD.t192 264.177
R1078 VDD.t246 VDD.t258 264.177
R1079 VDD.t130 VDD.t126 264.177
R1080 VDD.t32 VDD.t230 264.177
R1081 VDD.t105 VDD.t384 264.177
R1082 VDD.t66 VDD.t356 264.177
R1083 VDD.t112 VDD.t153 264.177
R1084 VDD.t50 VDD.t145 264.177
R1085 VDD.t436 VDD.t161 264.177
R1086 VDD.t182 VDD.t40 264.177
R1087 VDD.n726 VDD.n725 259.666
R1088 VDD.n2 VDD.n1 259.666
R1089 VDD.n575 VDD.n560 259.666
R1090 VDD.n5 VDD.n4 259.666
R1091 VDD.n514 VDD.n513 259.666
R1092 VDD.n82 VDD.n81 259.666
R1093 VDD.n992 VDD.n991 259.666
R1094 VDD.n383 VDD.t350 256.678
R1095 VDD.n121 VDD.t180 256.678
R1096 VDD.n1030 VDD.t420 256.678
R1097 VDD.n630 VDD.n628 253.44
R1098 VDD.n721 VDD.n720 252.16
R1099 VDD.n436 VDD.t394 248.603
R1100 VDD.n173 VDD.t310 248.603
R1101 VDD.n1083 VDD.t288 248.603
R1102 VDD.n494 VDD.t44 245.142
R1103 VDD.n231 VDD.t414 245.142
R1104 VDD.n1141 VDD.t326 245.142
R1105 VDD.n486 VDD.t360 240.528
R1106 VDD.n223 VDD.t344 240.528
R1107 VDD.n1133 VDD.t234 240.528
R1108 VDD.n444 VDD.t68 237.067
R1109 VDD.n181 VDD.t374 237.067
R1110 VDD.n1091 VDD.t24 237.067
R1111 VDD.n391 VDD.t418 228.992
R1112 VDD.n129 VDD.t176 228.992
R1113 VDD.n1038 VDD.t108 228.992
R1114 VDD.n663 VDD.t473 222.22
R1115 VDD.n375 VDD.t398 213.995
R1116 VDD.n113 VDD.t319 213.995
R1117 VDD.n1022 VDD.t73 213.995
R1118 VDD.n426 VDD.t200 205.919
R1119 VDD.n163 VDD.t354 205.919
R1120 VDD.n1073 VDD.t194 205.919
R1121 VDD.n504 VDD.t282 202.459
R1122 VDD.n241 VDD.t406 202.459
R1123 VDD.n1151 VDD.t272 202.459
R1124 VDD.n478 VDD.t110 197.844
R1125 VDD.n215 VDD.t358 197.844
R1126 VDD.n1125 VDD.t252 197.844
R1127 VDD.n452 VDD.t38 194.383
R1128 VDD.n189 VDD.t315 194.383
R1129 VDD.n1099 VDD.t184 194.383
R1130 VDD.n401 VDD.t101 186.308
R1131 VDD.n139 VDD.t270 186.308
R1132 VDD.n1048 VDD.t92 186.308
R1133 VDD.n731 VDD.n723 185
R1134 VDD.n670 VDD.n669 185
R1135 VDD.n678 VDD.n677 185
R1136 VDD.n618 VDD.n617 185
R1137 VDD.n559 VDD.n555 185
R1138 VDD.n558 VDD.n553 185
R1139 VDD.n557 VDD.n551 185
R1140 VDD.n350 VDD.n349 185
R1141 VDD.n358 VDD.n357 185
R1142 VDD.n368 VDD.n367 185
R1143 VDD.n376 VDD.n375 185
R1144 VDD.n384 VDD.n383 185
R1145 VDD.n392 VDD.n391 185
R1146 VDD.n402 VDD.n401 185
R1147 VDD.n410 VDD.n409 185
R1148 VDD.n418 VDD.n417 185
R1149 VDD.n427 VDD.n426 185
R1150 VDD.n437 VDD.n436 185
R1151 VDD.n445 VDD.n444 185
R1152 VDD.n453 VDD.n452 185
R1153 VDD.n461 VDD.n460 185
R1154 VDD.n471 VDD.n470 185
R1155 VDD.n479 VDD.n478 185
R1156 VDD.n487 VDD.n486 185
R1157 VDD.n495 VDD.n494 185
R1158 VDD.n505 VDD.n504 185
R1159 VDD.n286 VDD.n285 185
R1160 VDD.n519 VDD.n518 185
R1161 VDD.n88 VDD.n87 185
R1162 VDD.n96 VDD.n95 185
R1163 VDD.n106 VDD.n105 185
R1164 VDD.n114 VDD.n113 185
R1165 VDD.n122 VDD.n121 185
R1166 VDD.n130 VDD.n129 185
R1167 VDD.n140 VDD.n139 185
R1168 VDD.n148 VDD.n147 185
R1169 VDD.n156 VDD.n155 185
R1170 VDD.n164 VDD.n163 185
R1171 VDD.n174 VDD.n173 185
R1172 VDD.n182 VDD.n181 185
R1173 VDD.n190 VDD.n189 185
R1174 VDD.n198 VDD.n197 185
R1175 VDD.n208 VDD.n207 185
R1176 VDD.n216 VDD.n215 185
R1177 VDD.n224 VDD.n223 185
R1178 VDD.n232 VDD.n231 185
R1179 VDD.n242 VDD.n241 185
R1180 VDD.n250 VDD.n249 185
R1181 VDD.n997 VDD.n996 185
R1182 VDD.n1005 VDD.n1004 185
R1183 VDD.n1015 VDD.n1014 185
R1184 VDD.n1023 VDD.n1022 185
R1185 VDD.n1031 VDD.n1030 185
R1186 VDD.n1039 VDD.n1038 185
R1187 VDD.n1049 VDD.n1048 185
R1188 VDD.n1057 VDD.n1056 185
R1189 VDD.n1066 VDD.n1065 185
R1190 VDD.n1074 VDD.n1073 185
R1191 VDD.n1084 VDD.n1083 185
R1192 VDD.n1092 VDD.n1091 185
R1193 VDD.n1100 VDD.n1099 185
R1194 VDD.n1108 VDD.n1107 185
R1195 VDD.n1118 VDD.n1117 185
R1196 VDD.n1126 VDD.n1125 185
R1197 VDD.n1134 VDD.n1133 185
R1198 VDD.n1142 VDD.n1141 185
R1199 VDD.n1152 VDD.n1151 185
R1200 VDD.n928 VDD.n927 185
R1201 VDD.t442 VDD.n723 178.233
R1202 VDD.n669 VDD.t471 178.233
R1203 VDD.t59 VDD.n559 178.233
R1204 VDD.n349 VDD.t380 178.233
R1205 VDD.n518 VDD.t4 178.233
R1206 VDD.n87 VDD.t211 178.233
R1207 VDD.n996 VDD.t182 178.233
R1208 VDD.n617 VDD.t447 171.311
R1209 VDD.n557 VDD.t79 171.311
R1210 VDD.n367 VDD.t70 171.311
R1211 VDD.n105 VDD.t147 171.311
R1212 VDD.n1014 VDD.t198 171.311
R1213 VDD.n651 VDD.t452 166.1
R1214 VDD.n649 VDD.t467 166.1
R1215 VDD.n656 VDD.t461 166.1
R1216 VDD.n647 VDD.t455 166.1
R1217 VDD.n659 VDD.t464 166.1
R1218 VDD.n644 VDD.t449 166.1
R1219 VDD.n662 VDD.t470 166.1
R1220 VDD.n641 VDD.t446 166.099
R1221 VDD.n638 VDD.t479 166.098
R1222 VDD.n635 VDD.t476 166.098
R1223 VDD.n631 VDD.t458 166.097
R1224 VDD.n417 VDD.t120 163.236
R1225 VDD.n155 VDD.t362 163.236
R1226 VDD.n1065 VDD.t262 163.236
R1227 VDD.n285 VDD.t227 159.775
R1228 VDD.n249 VDD.t428 159.775
R1229 VDD.n927 VDD.t151 159.775
R1230 VDD.n470 VDD.t215 155.16
R1231 VDD.n207 VDD.t330 155.16
R1232 VDD.n1117 VDD.t155 155.16
R1233 VDD.n460 VDD.t94 151.7
R1234 VDD.n197 VDD.t260 151.7
R1235 VDD.n1107 VDD.t85 151.7
R1236 VDD.n717 sky130_asc_pfet_01v8_lvt_6_0/SOURCE 147.84
R1237 VDD.n624 sky130_asc_pfet_01v8_lvt_12_0/SOURCE 147.84
R1238 VDD.n566 sky130_asc_pfet_01v8_lvt_12_1/SOURCE 147.84
R1239 VDD.n304 sky130_asc_pfet_01v8_lvt_60_2/SOURCE 147.84
R1240 VDD.n281 sky130_asc_pfet_01v8_lvt_6_1/SOURCE 147.84
R1241 VDD.n42 sky130_asc_pfet_01v8_lvt_60_1/SOURCE 147.84
R1242 VDD.n947 sky130_asc_pfet_01v8_lvt_60_0/SOURCE 147.84
R1243 VDD.n409 VDD.t438 143.624
R1244 VDD.n147 VDD.t149 143.624
R1245 VDD.n1056 VDD.t170 143.624
R1246 VDD.n677 VDD.t453 135.549
R1247 VDD.t412 VDD.n558 135.549
R1248 VDD.n357 VDD.t48 135.549
R1249 VDD.n95 VDD.t305 135.549
R1250 VDD.n1004 VDD.t83 135.549
R1251 VDD.n677 VDD.t468 128.627
R1252 VDD.n558 VDD.t386 128.627
R1253 VDD.n357 VDD.t426 128.627
R1254 VDD.n95 VDD.t254 128.627
R1255 VDD.n1004 VDD.t77 128.627
R1256 VDD.n409 VDD.t225 120.552
R1257 VDD.n147 VDD.t196 120.552
R1258 VDD.n1056 VDD.t213 120.552
R1259 VDD.n460 VDD.t81 112.477
R1260 VDD.n197 VDD.t256 112.477
R1261 VDD.n1107 VDD.t223 112.477
R1262 VDD.n470 VDD.t207 109.016
R1263 VDD.n207 VDD.t244 109.016
R1264 VDD.n1117 VDD.t157 109.016
R1265 VDD.n285 VDD.t172 104.401
R1266 VDD.n249 VDD.t424 104.401
R1267 VDD.n927 VDD.t278 104.401
R1268 VDD.n417 VDD.t203 100.941
R1269 VDD.n155 VDD.t294 100.941
R1270 VDD.n1065 VDD.t130 100.941
R1271 VDD.n657 VDD.n656 100.256
R1272 VDD.n636 VDD.n635 96.4
R1273 VDD.n617 VDD.t450 92.865
R1274 VDD.t34 VDD.n557 92.865
R1275 VDD.n367 VDD.t402 92.865
R1276 VDD.n105 VDD.t242 92.865
R1277 VDD.n1014 VDD.t50 92.865
R1278 VDD.n737 VDD.n715 89.983
R1279 VDD.n632 VDD.n631 87.568
R1280 VDD.n723 VDD.t482 85.944
R1281 VDD.n669 VDD.t465 85.944
R1282 VDD.n559 VDD.t422 85.944
R1283 VDD.n349 VDD.t378 85.944
R1284 VDD.n518 VDD.t492 85.944
R1285 VDD.n87 VDD.t205 85.944
R1286 VDD.n996 VDD.t436 85.944
R1287 VDD.n726 VDD.n724 85.333
R1288 VDD.n733 VDD.n715 85.333
R1289 VDD.n733 VDD.n732 85.333
R1290 VDD.n634 VDD.n632 85.333
R1291 VDD.n637 VDD.n634 85.333
R1292 VDD.n640 VDD.n637 85.333
R1293 VDD.n643 VDD.n640 85.333
R1294 VDD.n646 VDD.n643 85.333
R1295 VDD.n648 VDD.n646 85.333
R1296 VDD.n650 VDD.n648 85.333
R1297 VDD.n653 VDD.n650 85.333
R1298 VDD.n655 VDD.n653 85.333
R1299 VDD.n658 VDD.n655 85.333
R1300 VDD.n661 VDD.n658 85.333
R1301 VDD.n576 VDD.n575 85.333
R1302 VDD.n582 VDD.n581 85.333
R1303 VDD.n581 VDD.n580 85.333
R1304 VDD.n587 VDD.n586 85.333
R1305 VDD.n586 VDD.n585 85.333
R1306 VDD.n730 VDD.n724 82.651
R1307 VDD.n577 VDD.n576 82.651
R1308 VDD.n401 VDD.t376 77.868
R1309 VDD.n139 VDD.t209 77.868
R1310 VDD.n1048 VDD.t32 77.868
R1311 VDD.n634 VDD.n633 76
R1312 VDD.n637 VDD.n636 76
R1313 VDD.n640 VDD.n639 76
R1314 VDD.n643 VDD.n642 76
R1315 VDD.n646 VDD.n645 76
R1316 VDD.n648 VDD.n647 76
R1317 VDD.n650 VDD.n649 76
R1318 VDD.n653 VDD.n652 76
R1319 VDD.n655 VDD.n654 76
R1320 VDD.n658 VDD.n657 76
R1321 VDD.n661 VDD.n660 76
R1322 VDD.n664 VDD.n661 75.52
R1323 VDD.n660 VDD.n659 73.264
R1324 VDD.n630 VDD.n629 72.504
R1325 VDD.n663 VDD.n662 69.888
R1326 VDD.n452 VDD.t178 69.793
R1327 VDD.n189 VDD.t128 69.793
R1328 VDD.n1099 VDD.t99 69.793
R1329 VDD.n639 VDD.n638 69.408
R1330 VDD.n478 VDD.t190 66.332
R1331 VDD.n215 VDD.t392 66.332
R1332 VDD.n1125 VDD.t302 66.332
R1333 VDD.n732 VDD.n731 63.024
R1334 VDD.n580 VDD.n555 63.024
R1335 VDD.n504 VDD.t238 61.718
R1336 VDD.n241 VDD.t370 61.718
R1337 VDD.n1151 VDD.t382 61.718
R1338 VDD.n426 VDD.t46 58.257
R1339 VDD.n163 VDD.t26 58.257
R1340 VDD.n1073 VDD.t246 58.257
R1341 VDD.n375 VDD.t400 50.182
R1342 VDD.n113 VDD.t284 50.182
R1343 VDD.n1022 VDD.t112 50.182
R1344 VDD.n664 VDD.n663 46.684
R1345 VDD.n587 VDD.n551 45.47
R1346 VDD.n642 VDD.n641 42.416
R1347 VDD.n585 VDD.n553 41.691
R1348 VDD.n721 VDD.n717 40.96
R1349 VDD.n391 VDD.t396 35.185
R1350 VDD.n129 VDD.t159 35.185
R1351 VDD.n1038 VDD.t105 35.185
R1352 VDD.n632 sky130_asc_pfet_01v8_lvt_12_0/GATE 34.986
R1353 VDD.n720 VDD.n718 32.824
R1354 VDD.n717 VDD.n716 32.824
R1355 VDD.n628 VDD.n619 32.824
R1356 VDD.n627 VDD.n620 32.824
R1357 VDD.n626 VDD.n621 32.824
R1358 VDD.n625 VDD.n622 32.824
R1359 VDD.n624 VDD.n623 32.824
R1360 VDD.n570 VDD.n561 32.824
R1361 VDD.n569 VDD.n562 32.824
R1362 VDD.n568 VDD.n563 32.824
R1363 VDD.n567 VDD.n564 32.824
R1364 VDD.n566 VDD.n565 32.824
R1365 VDD.n333 VDD.n331 32.824
R1366 VDD.n334 VDD.n330 32.824
R1367 VDD.n335 VDD.n329 32.824
R1368 VDD.n336 VDD.n328 32.824
R1369 VDD.n337 VDD.n327 32.824
R1370 VDD.n338 VDD.n326 32.824
R1371 VDD.n339 VDD.n325 32.824
R1372 VDD.n340 VDD.n324 32.824
R1373 VDD.n341 VDD.n323 32.824
R1374 VDD.n342 VDD.n322 32.824
R1375 VDD.n343 VDD.n321 32.824
R1376 VDD.n320 VDD.n287 32.824
R1377 VDD.n319 VDD.n288 32.824
R1378 VDD.n318 VDD.n289 32.824
R1379 VDD.n317 VDD.n290 32.824
R1380 VDD.n316 VDD.n291 32.824
R1381 VDD.n315 VDD.n292 32.824
R1382 VDD.n314 VDD.n293 32.824
R1383 VDD.n313 VDD.n294 32.824
R1384 VDD.n312 VDD.n295 32.824
R1385 VDD.n311 VDD.n296 32.824
R1386 VDD.n310 VDD.n297 32.824
R1387 VDD.n309 VDD.n298 32.824
R1388 VDD.n308 VDD.n299 32.824
R1389 VDD.n307 VDD.n300 32.824
R1390 VDD.n306 VDD.n301 32.824
R1391 VDD.n305 VDD.n302 32.824
R1392 VDD.n304 VDD.n303 32.824
R1393 VDD.n281 VDD.n280 32.824
R1394 VDD.n70 VDD.n13 32.824
R1395 VDD.n69 VDD.n14 32.824
R1396 VDD.n68 VDD.n15 32.824
R1397 VDD.n67 VDD.n16 32.824
R1398 VDD.n66 VDD.n17 32.824
R1399 VDD.n65 VDD.n18 32.824
R1400 VDD.n64 VDD.n19 32.824
R1401 VDD.n63 VDD.n20 32.824
R1402 VDD.n62 VDD.n21 32.824
R1403 VDD.n61 VDD.n22 32.824
R1404 VDD.n60 VDD.n23 32.824
R1405 VDD.n59 VDD.n24 32.824
R1406 VDD.n58 VDD.n25 32.824
R1407 VDD.n57 VDD.n26 32.824
R1408 VDD.n56 VDD.n27 32.824
R1409 VDD.n55 VDD.n28 32.824
R1410 VDD.n54 VDD.n29 32.824
R1411 VDD.n53 VDD.n30 32.824
R1412 VDD.n52 VDD.n31 32.824
R1413 VDD.n51 VDD.n32 32.824
R1414 VDD.n50 VDD.n33 32.824
R1415 VDD.n49 VDD.n34 32.824
R1416 VDD.n48 VDD.n35 32.824
R1417 VDD.n47 VDD.n36 32.824
R1418 VDD.n46 VDD.n37 32.824
R1419 VDD.n45 VDD.n38 32.824
R1420 VDD.n44 VDD.n39 32.824
R1421 VDD.n43 VDD.n40 32.824
R1422 VDD.n42 VDD.n41 32.824
R1423 VDD.n976 VDD.n974 32.824
R1424 VDD.n977 VDD.n973 32.824
R1425 VDD.n978 VDD.n972 32.824
R1426 VDD.n979 VDD.n971 32.824
R1427 VDD.n980 VDD.n970 32.824
R1428 VDD.n981 VDD.n969 32.824
R1429 VDD.n982 VDD.n968 32.824
R1430 VDD.n983 VDD.n967 32.824
R1431 VDD.n984 VDD.n966 32.824
R1432 VDD.n985 VDD.n965 32.824
R1433 VDD.n964 VDD.n929 32.824
R1434 VDD.n963 VDD.n930 32.824
R1435 VDD.n962 VDD.n931 32.824
R1436 VDD.n961 VDD.n932 32.824
R1437 VDD.n960 VDD.n933 32.824
R1438 VDD.n959 VDD.n934 32.824
R1439 VDD.n958 VDD.n935 32.824
R1440 VDD.n957 VDD.n936 32.824
R1441 VDD.n956 VDD.n937 32.824
R1442 VDD.n955 VDD.n938 32.824
R1443 VDD.n954 VDD.n939 32.824
R1444 VDD.n953 VDD.n940 32.824
R1445 VDD.n952 VDD.n941 32.824
R1446 VDD.n951 VDD.n942 32.824
R1447 VDD.n950 VDD.n943 32.824
R1448 VDD.n949 VDD.n944 32.824
R1449 VDD.n948 VDD.n945 32.824
R1450 VDD.n947 VDD.n946 32.824
R1451 VDD.n284 VDD.n283 31.801
R1452 VDD.n346 VDD.n344 31.801
R1453 VDD.n988 VDD.n986 31.801
R1454 VDD.n444 VDD.t64 27.109
R1455 VDD.n181 VDD.t372 27.109
R1456 VDD.n1091 VDD.t61 27.109
R1457 VDD.n687 VDD.n618 24.758
R1458 VDD.n589 VDD.n551 24.758
R1459 VDD.n679 VDD.n678 24.137
R1460 VDD.n582 VDD.n553 24.137
R1461 VDD.n359 VDD.n358 24.137
R1462 VDD.n393 VDD.n392 24.137
R1463 VDD.n428 VDD.n427 24.137
R1464 VDD.n462 VDD.n461 24.137
R1465 VDD.n496 VDD.n495 24.137
R1466 VDD.n97 VDD.n96 24.137
R1467 VDD.n131 VDD.n130 24.137
R1468 VDD.n165 VDD.n164 24.137
R1469 VDD.n199 VDD.n198 24.137
R1470 VDD.n233 VDD.n232 24.137
R1471 VDD.n1006 VDD.n1005 24.137
R1472 VDD.n1040 VDD.n1039 24.137
R1473 VDD.n1075 VDD.n1074 24.137
R1474 VDD.n1109 VDD.n1108 24.137
R1475 VDD.n1143 VDD.n1142 24.137
R1476 VDD.n486 VDD.t248 23.649
R1477 VDD.n223 VDD.t352 23.649
R1478 VDD.n1133 VDD.t236 23.649
R1479 VDD.n369 VDD.n368 20.357
R1480 VDD.n403 VDD.n402 20.357
R1481 VDD.n438 VDD.n437 20.357
R1482 VDD.n472 VDD.n471 20.357
R1483 VDD.n506 VDD.n505 20.357
R1484 VDD.n107 VDD.n106 20.357
R1485 VDD.n141 VDD.n140 20.357
R1486 VDD.n175 VDD.n174 20.357
R1487 VDD.n209 VDD.n208 20.357
R1488 VDD.n243 VDD.n242 20.357
R1489 VDD.n1016 VDD.n1015 20.357
R1490 VDD.n1050 VDD.n1049 20.357
R1491 VDD.n1085 VDD.n1084 20.357
R1492 VDD.n1119 VDD.n1118 20.357
R1493 VDD.n1153 VDD.n1152 20.357
R1494 VDD.n494 VDD.t232 19.034
R1495 VDD.n231 VDD.t410 19.034
R1496 VDD.n1141 VDD.t323 19.034
R1497 VDD.n436 VDD.t188 15.573
R1498 VDD.n173 VDD.t388 15.573
R1499 VDD.n1083 VDD.t292 15.573
R1500 VDD.n645 VDD.n644 15.424
R1501 sky130_asc_res_xhigh_po_2p85_1_8/VPWR sky130_asc_pnp_05v5_W3p40L3p40_8_1/VPWR 11.947
R1502 sky130_asc_res_xhigh_po_2p85_1_0/VPWR sky130_asc_pnp_05v5_W3p40L3p40_8_2/VPWR 11.947
R1503 sky130_asc_res_xhigh_po_2p85_1_16/VPWR sky130_asc_pnp_05v5_W3p40L3p40_8_3/VPWR 11.437
R1504 sky130_asc_res_xhigh_po_2p85_1_17/VPWR sky130_asc_pnp_05v5_W3p40L3p40_8_0/VPWR 11.437
R1505 VDD.n665 VDD.n664 11.352
R1506 sky130_asc_pnp_05v5_W3p40L3p40_7_0/VPWR sky130_asc_res_xhigh_po_2p85_1_19/VPWR 10.111
R1507 VDD.n727 sky130_asc_cap_mim_m3_1_7/VPWR 8.345
R1508 VDD.n512 VDD.n286 8.045
R1509 VDD.n251 VDD.n250 8.045
R1510 VDD.n1159 VDD.n928 8.045
R1511 sky130_asc_nfet_01v8_lvt_9_1/VPWR sky130_asc_cap_mim_m3_1_9/VPWR 7.83
R1512 sky130_asc_res_xhigh_po_2p85_2_0/VPWR sky130_asc_cap_mim_m3_1_8/VPWR 7.751
R1513 sky130_asc_res_xhigh_po_2p85_1_22/VPWR sky130_asc_cap_mim_m3_1_6/VPWR 7.749
R1514 sky130_asc_pnp_05v5_W3p40L3p40_1_0/VPWR sky130_asc_cap_mim_m3_1_5/VPWR 7.728
R1515 VDD.n652 VDD.n651 7.712
R1516 VDD.n383 VDD.t42 7.498
R1517 VDD.n121 VDD.t52 7.498
R1518 VDD.n1030 VDD.t66 7.498
R1519 sky130_asc_cap_mim_m3_1_0/VPWR VDD.n870 7.376
R1520 sky130_asc_cap_mim_m3_1_1/VPWR VDD.n885 7.368
R1521 sky130_asc_res_xhigh_po_2p85_1_1/VPWR sky130_asc_res_xhigh_po_2p85_2_1/VPWR 6.634
R1522 VDD.n816 sky130_asc_res_xhigh_po_2p85_1_15/VPWR 6.167
R1523 VDD.n792 sky130_asc_res_xhigh_po_2p85_1_12/VPWR 6.068
R1524 VDD.n990 sky130_asc_cap_mim_m3_1_4/VPWR 5.879
R1525 sky130_asc_pnp_05v5_W3p40L3p40_8_1/VPWR sky130_asc_nfet_01v8_lvt_9_2/VPWR 5.498
R1526 sky130_asc_pnp_05v5_W3p40L3p40_8_2/VPWR sky130_asc_nfet_01v8_lvt_9_1/VPWR 5.498
R1527 VDD.n731 VDD.n730 5.485
R1528 VDD.n671 VDD.n670 5.485
R1529 VDD.n577 VDD.n555 5.485
R1530 VDD.n351 VDD.n350 5.485
R1531 VDD.n385 VDD.n384 5.485
R1532 VDD.n419 VDD.n418 5.485
R1533 VDD.n454 VDD.n453 5.485
R1534 VDD.n488 VDD.n487 5.485
R1535 VDD.n520 VDD.n519 5.485
R1536 VDD.n89 VDD.n88 5.485
R1537 VDD.n123 VDD.n122 5.485
R1538 VDD.n157 VDD.n156 5.485
R1539 VDD.n191 VDD.n190 5.485
R1540 VDD.n225 VDD.n224 5.485
R1541 VDD.n998 VDD.n997 5.485
R1542 VDD.n1032 VDD.n1031 5.485
R1543 VDD.n1067 VDD.n1066 5.485
R1544 VDD.n1101 VDD.n1100 5.485
R1545 VDD.n1135 VDD.n1134 5.485
R1546 VDD.n990 VDD.n989 5.164
R1547 VDD.n736 VDD.n721 5.096
R1548 sky130_asc_pnp_05v5_W3p40L3p40_8_3/VPWR sky130_asc_res_xhigh_po_2p85_1_22/VPWR 4.876
R1549 sky130_asc_res_xhigh_po_2p85_1_5/VPWR sky130_asc_nfet_01v8_lvt_9_0/VPWR 4.804
R1550 VDD.n735 VDD.n715 4.65
R1551 VDD.n734 VDD.n733 4.65
R1552 VDD.n732 VDD.n722 4.65
R1553 VDD.n730 VDD.n729 4.65
R1554 VDD.n728 VDD.n724 4.65
R1555 VDD.n727 VDD.n726 4.65
R1556 VDD.n686 VDD.n685 4.65
R1557 VDD.n684 VDD.n683 4.65
R1558 VDD.n682 VDD.n681 4.65
R1559 VDD.n680 VDD.n679 4.65
R1560 VDD.n676 VDD.n675 4.65
R1561 VDD.n674 VDD.n673 4.65
R1562 VDD.n672 VDD.n671 4.65
R1563 VDD.n667 VDD.n666 4.65
R1564 VDD.n3 VDD.n2 4.65
R1565 VDD.n588 VDD.n587 4.65
R1566 VDD.n586 VDD.n552 4.65
R1567 VDD.n585 VDD.n584 4.65
R1568 VDD.n583 VDD.n582 4.65
R1569 VDD.n581 VDD.n554 4.65
R1570 VDD.n580 VDD.n579 4.65
R1571 VDD.n578 VDD.n577 4.65
R1572 VDD.n576 VDD.n556 4.65
R1573 VDD.n575 VDD.n574 4.65
R1574 VDD.n521 VDD.n520 4.65
R1575 VDD.n517 VDD.n516 4.65
R1576 VDD.n515 VDD.n514 4.65
R1577 VDD.n511 VDD.n510 4.65
R1578 VDD.n509 VDD.n508 4.65
R1579 VDD.n507 VDD.n506 4.65
R1580 VDD.n503 VDD.n502 4.65
R1581 VDD.n501 VDD.n500 4.65
R1582 VDD.n499 VDD.n498 4.65
R1583 VDD.n497 VDD.n496 4.65
R1584 VDD.n493 VDD.n492 4.65
R1585 VDD.n491 VDD.n490 4.65
R1586 VDD.n489 VDD.n488 4.65
R1587 VDD.n485 VDD.n484 4.65
R1588 VDD.n483 VDD.n482 4.65
R1589 VDD.n481 VDD.n480 4.65
R1590 VDD.n477 VDD.n476 4.65
R1591 VDD.n475 VDD.n474 4.65
R1592 VDD.n473 VDD.n472 4.65
R1593 VDD.n469 VDD.n468 4.65
R1594 VDD.n467 VDD.n466 4.65
R1595 VDD.n465 VDD.n464 4.65
R1596 VDD.n463 VDD.n462 4.65
R1597 VDD.n459 VDD.n458 4.65
R1598 VDD.n457 VDD.n456 4.65
R1599 VDD.n455 VDD.n454 4.65
R1600 VDD.n451 VDD.n450 4.65
R1601 VDD.n449 VDD.n448 4.65
R1602 VDD.n447 VDD.n446 4.65
R1603 VDD.n443 VDD.n442 4.65
R1604 VDD.n441 VDD.n440 4.65
R1605 VDD.n439 VDD.n438 4.65
R1606 VDD.n435 VDD.n434 4.65
R1607 VDD.n433 VDD.n432 4.65
R1608 VDD.n431 VDD.n430 4.65
R1609 VDD.n429 VDD.n428 4.65
R1610 VDD.n425 VDD.n424 4.65
R1611 VDD.n423 VDD.n422 4.65
R1612 VDD.n420 VDD.n419 4.65
R1613 VDD.n416 VDD.n415 4.65
R1614 VDD.n414 VDD.n413 4.65
R1615 VDD.n412 VDD.n411 4.65
R1616 VDD.n408 VDD.n407 4.65
R1617 VDD.n406 VDD.n405 4.65
R1618 VDD.n404 VDD.n403 4.65
R1619 VDD.n400 VDD.n399 4.65
R1620 VDD.n398 VDD.n397 4.65
R1621 VDD.n396 VDD.n395 4.65
R1622 VDD.n394 VDD.n393 4.65
R1623 VDD.n390 VDD.n389 4.65
R1624 VDD.n388 VDD.n387 4.65
R1625 VDD.n386 VDD.n385 4.65
R1626 VDD.n382 VDD.n381 4.65
R1627 VDD.n380 VDD.n379 4.65
R1628 VDD.n378 VDD.n377 4.65
R1629 VDD.n374 VDD.n373 4.65
R1630 VDD.n372 VDD.n371 4.65
R1631 VDD.n370 VDD.n369 4.65
R1632 VDD.n366 VDD.n365 4.65
R1633 VDD.n364 VDD.n363 4.65
R1634 VDD.n362 VDD.n361 4.65
R1635 VDD.n360 VDD.n359 4.65
R1636 VDD.n356 VDD.n355 4.65
R1637 VDD.n354 VDD.n353 4.65
R1638 VDD.n352 VDD.n351 4.65
R1639 VDD.n348 VDD.n347 4.65
R1640 VDD.n6 VDD.n5 4.65
R1641 VDD.n248 VDD.n247 4.65
R1642 VDD.n246 VDD.n245 4.65
R1643 VDD.n244 VDD.n243 4.65
R1644 VDD.n240 VDD.n239 4.65
R1645 VDD.n238 VDD.n237 4.65
R1646 VDD.n236 VDD.n235 4.65
R1647 VDD.n234 VDD.n233 4.65
R1648 VDD.n230 VDD.n229 4.65
R1649 VDD.n228 VDD.n227 4.65
R1650 VDD.n226 VDD.n225 4.65
R1651 VDD.n222 VDD.n221 4.65
R1652 VDD.n220 VDD.n219 4.65
R1653 VDD.n218 VDD.n217 4.65
R1654 VDD.n214 VDD.n213 4.65
R1655 VDD.n212 VDD.n211 4.65
R1656 VDD.n210 VDD.n209 4.65
R1657 VDD.n206 VDD.n205 4.65
R1658 VDD.n204 VDD.n203 4.65
R1659 VDD.n202 VDD.n201 4.65
R1660 VDD.n200 VDD.n199 4.65
R1661 VDD.n196 VDD.n195 4.65
R1662 VDD.n194 VDD.n193 4.65
R1663 VDD.n192 VDD.n191 4.65
R1664 VDD.n188 VDD.n187 4.65
R1665 VDD.n186 VDD.n185 4.65
R1666 VDD.n184 VDD.n183 4.65
R1667 VDD.n180 VDD.n179 4.65
R1668 VDD.n178 VDD.n177 4.65
R1669 VDD.n176 VDD.n175 4.65
R1670 VDD.n172 VDD.n171 4.65
R1671 VDD.n170 VDD.n169 4.65
R1672 VDD.n168 VDD.n167 4.65
R1673 VDD.n166 VDD.n165 4.65
R1674 VDD.n162 VDD.n161 4.65
R1675 VDD.n160 VDD.n159 4.65
R1676 VDD.n158 VDD.n157 4.65
R1677 VDD.n154 VDD.n153 4.65
R1678 VDD.n152 VDD.n151 4.65
R1679 VDD.n150 VDD.n149 4.65
R1680 VDD.n146 VDD.n145 4.65
R1681 VDD.n144 VDD.n143 4.65
R1682 VDD.n142 VDD.n141 4.65
R1683 VDD.n138 VDD.n137 4.65
R1684 VDD.n136 VDD.n135 4.65
R1685 VDD.n134 VDD.n133 4.65
R1686 VDD.n132 VDD.n131 4.65
R1687 VDD.n128 VDD.n127 4.65
R1688 VDD.n126 VDD.n125 4.65
R1689 VDD.n124 VDD.n123 4.65
R1690 VDD.n120 VDD.n119 4.65
R1691 VDD.n118 VDD.n117 4.65
R1692 VDD.n116 VDD.n115 4.65
R1693 VDD.n112 VDD.n111 4.65
R1694 VDD.n110 VDD.n109 4.65
R1695 VDD.n108 VDD.n107 4.65
R1696 VDD.n104 VDD.n103 4.65
R1697 VDD.n102 VDD.n101 4.65
R1698 VDD.n100 VDD.n99 4.65
R1699 VDD.n98 VDD.n97 4.65
R1700 VDD.n94 VDD.n93 4.65
R1701 VDD.n92 VDD.n91 4.65
R1702 VDD.n90 VDD.n89 4.65
R1703 VDD.n86 VDD.n85 4.65
R1704 VDD.n83 VDD.n82 4.65
R1705 VDD.n1158 VDD.n1157 4.65
R1706 VDD.n1156 VDD.n1155 4.65
R1707 VDD.n1154 VDD.n1153 4.65
R1708 VDD.n1150 VDD.n1149 4.65
R1709 VDD.n1148 VDD.n1147 4.65
R1710 VDD.n1146 VDD.n1145 4.65
R1711 VDD.n1144 VDD.n1143 4.65
R1712 VDD.n1140 VDD.n1139 4.65
R1713 VDD.n1138 VDD.n1137 4.65
R1714 VDD.n1136 VDD.n1135 4.65
R1715 VDD.n1132 VDD.n1131 4.65
R1716 VDD.n1130 VDD.n1129 4.65
R1717 VDD.n1128 VDD.n1127 4.65
R1718 VDD.n1124 VDD.n1123 4.65
R1719 VDD.n1122 VDD.n1121 4.65
R1720 VDD.n1120 VDD.n1119 4.65
R1721 VDD.n1116 VDD.n1115 4.65
R1722 VDD.n1114 VDD.n1113 4.65
R1723 VDD.n1112 VDD.n1111 4.65
R1724 VDD.n1110 VDD.n1109 4.65
R1725 VDD.n1106 VDD.n1105 4.65
R1726 VDD.n1104 VDD.n1103 4.65
R1727 VDD.n1102 VDD.n1101 4.65
R1728 VDD.n1098 VDD.n1097 4.65
R1729 VDD.n1096 VDD.n1095 4.65
R1730 VDD.n1094 VDD.n1093 4.65
R1731 VDD.n1090 VDD.n1089 4.65
R1732 VDD.n1088 VDD.n1087 4.65
R1733 VDD.n1086 VDD.n1085 4.65
R1734 VDD.n1082 VDD.n1081 4.65
R1735 VDD.n1080 VDD.n1079 4.65
R1736 VDD.n1078 VDD.n1077 4.65
R1737 VDD.n1076 VDD.n1075 4.65
R1738 VDD.n1072 VDD.n1071 4.65
R1739 VDD.n1070 VDD.n1069 4.65
R1740 VDD.n1068 VDD.n1067 4.65
R1741 VDD.n1064 VDD.n1063 4.65
R1742 VDD.n1062 VDD.n1061 4.65
R1743 VDD.n1059 VDD.n1058 4.65
R1744 VDD.n1055 VDD.n1054 4.65
R1745 VDD.n1053 VDD.n1052 4.65
R1746 VDD.n1051 VDD.n1050 4.65
R1747 VDD.n1047 VDD.n1046 4.65
R1748 VDD.n1045 VDD.n1044 4.65
R1749 VDD.n1043 VDD.n1042 4.65
R1750 VDD.n1041 VDD.n1040 4.65
R1751 VDD.n1037 VDD.n1036 4.65
R1752 VDD.n1035 VDD.n1034 4.65
R1753 VDD.n1033 VDD.n1032 4.65
R1754 VDD.n1029 VDD.n1028 4.65
R1755 VDD.n1027 VDD.n1026 4.65
R1756 VDD.n1025 VDD.n1024 4.65
R1757 VDD.n1021 VDD.n1020 4.65
R1758 VDD.n1019 VDD.n1018 4.65
R1759 VDD.n1017 VDD.n1016 4.65
R1760 VDD.n1013 VDD.n1012 4.65
R1761 VDD.n1011 VDD.n1010 4.65
R1762 VDD.n1009 VDD.n1008 4.65
R1763 VDD.n1007 VDD.n1006 4.65
R1764 VDD.n1003 VDD.n1002 4.65
R1765 VDD.n1001 VDD.n1000 4.65
R1766 VDD.n999 VDD.n998 4.65
R1767 VDD.n995 VDD.n994 4.65
R1768 VDD.n993 VDD.n992 4.65
R1769 VDD.n765 sky130_asc_res_xhigh_po_2p85_1_16/VPWR 4.639
R1770 VDD.n738 sky130_asc_res_xhigh_po_2p85_1_17/VPWR 4.639
R1771 VDD.n83 VDD.n80 4.507
R1772 VDD.n719 VDD.t443 4.428
R1773 VDD.n719 VDD.t441 4.428
R1774 VDD.n718 VDD.t485 4.428
R1775 VDD.n718 VDD.t483 4.428
R1776 VDD.n716 VDD.t491 4.428
R1777 VDD.n716 VDD.t489 4.428
R1778 VDD.n629 VDD.t472 4.428
R1779 VDD.n629 VDD.t475 4.428
R1780 VDD.n619 VDD.t463 4.428
R1781 VDD.n619 VDD.t466 4.428
R1782 VDD.n620 VDD.t469 4.428
R1783 VDD.n620 VDD.t454 4.428
R1784 VDD.n621 VDD.t451 4.428
R1785 VDD.n621 VDD.t457 4.428
R1786 VDD.n622 VDD.t481 4.428
R1787 VDD.n622 VDD.t448 4.428
R1788 VDD.n623 VDD.t460 4.428
R1789 VDD.n623 VDD.t478 4.428
R1790 VDD.n571 VDD.t60 4.428
R1791 VDD.n571 VDD.t417 4.428
R1792 VDD.n561 VDD.t347 4.428
R1793 VDD.n561 VDD.t423 4.428
R1794 VDD.n562 VDD.t387 4.428
R1795 VDD.n562 VDD.t413 4.428
R1796 VDD.n563 VDD.t35 4.428
R1797 VDD.n563 VDD.t97 4.428
R1798 VDD.n564 VDD.t435 4.428
R1799 VDD.n564 VDD.t80 4.428
R1800 VDD.n565 VDD.t135 4.428
R1801 VDD.n565 VDD.t431 4.428
R1802 VDD.n345 VDD.t121 4.428
R1803 VDD.n345 VDD.t204 4.428
R1804 VDD.n332 VDD.t381 4.428
R1805 VDD.n332 VDD.t314 4.428
R1806 VDD.n331 VDD.t7 4.428
R1807 VDD.n331 VDD.t379 4.428
R1808 VDD.n330 VDD.t427 4.428
R1809 VDD.n330 VDD.t49 4.428
R1810 VDD.n329 VDD.t403 4.428
R1811 VDD.n329 VDD.t405 4.428
R1812 VDD.n328 VDD.t333 4.428
R1813 VDD.n328 VDD.t71 4.428
R1814 VDD.n327 VDD.t399 4.428
R1815 VDD.n327 VDD.t401 4.428
R1816 VDD.n326 VDD.t43 4.428
R1817 VDD.n326 VDD.t365 4.428
R1818 VDD.n325 VDD.t419 4.428
R1819 VDD.n325 VDD.t351 4.428
R1820 VDD.n324 VDD.t104 4.428
R1821 VDD.n324 VDD.t397 4.428
R1822 VDD.n323 VDD.t377 4.428
R1823 VDD.n323 VDD.t102 4.428
R1824 VDD.n322 VDD.t439 4.428
R1825 VDD.n322 VDD.t90 4.428
R1826 VDD.n321 VDD.t164 4.428
R1827 VDD.n321 VDD.t226 4.428
R1828 VDD.n287 VDD.t47 4.428
R1829 VDD.n287 VDD.t115 4.428
R1830 VDD.n288 VDD.t241 4.428
R1831 VDD.n288 VDD.t201 4.428
R1832 VDD.n289 VDD.t395 4.428
R1833 VDD.n289 VDD.t189 4.428
R1834 VDD.n290 VDD.t65 4.428
R1835 VDD.n290 VDD.t69 4.428
R1836 VDD.n291 VDD.t39 4.428
R1837 VDD.n291 VDD.t55 4.428
R1838 VDD.n292 VDD.t175 4.428
R1839 VDD.n292 VDD.t179 4.428
R1840 VDD.n293 VDD.t82 4.428
R1841 VDD.n293 VDD.t95 4.428
R1842 VDD.n294 VDD.t208 4.428
R1843 VDD.n294 VDD.t76 4.428
R1844 VDD.n295 VDD.t133 4.428
R1845 VDD.n295 VDD.t216 4.428
R1846 VDD.n296 VDD.t111 4.428
R1847 VDD.n296 VDD.t191 4.428
R1848 VDD.n297 VDD.t249 4.428
R1849 VDD.n297 VDD.t297 4.428
R1850 VDD.n298 VDD.t45 4.428
R1851 VDD.n298 VDD.t361 4.428
R1852 VDD.n299 VDD.t318 4.428
R1853 VDD.n299 VDD.t233 4.428
R1854 VDD.n300 VDD.t239 4.428
R1855 VDD.n300 VDD.t283 4.428
R1856 VDD.n301 VDD.t228 4.428
R1857 VDD.n301 VDD.t31 4.428
R1858 VDD.n302 VDD.t169 4.428
R1859 VDD.n302 VDD.t173 4.428
R1860 VDD.n303 VDD.t123 4.428
R1861 VDD.n303 VDD.t275 4.428
R1862 VDD.n279 VDD.t445 4.428
R1863 VDD.n279 VDD.t493 4.428
R1864 VDD.n282 VDD.t5 4.428
R1865 VDD.n282 VDD.t1 4.428
R1866 VDD.n280 VDD.t487 4.428
R1867 VDD.n280 VDD.t3 4.428
R1868 VDD.n71 VDD.t212 4.428
R1869 VDD.n71 VDD.t222 4.428
R1870 VDD.n13 VDD.t119 4.428
R1871 VDD.n13 VDD.t206 4.428
R1872 VDD.n14 VDD.t255 4.428
R1873 VDD.n14 VDD.t306 4.428
R1874 VDD.n15 VDD.t243 4.428
R1875 VDD.n15 VDD.t29 4.428
R1876 VDD.n16 VDD.t329 4.428
R1877 VDD.n16 VDD.t148 4.428
R1878 VDD.n17 VDD.t320 4.428
R1879 VDD.n17 VDD.t285 4.428
R1880 VDD.n18 VDD.t53 4.428
R1881 VDD.n18 VDD.t277 4.428
R1882 VDD.n19 VDD.t177 4.428
R1883 VDD.n19 VDD.t181 4.428
R1884 VDD.n20 VDD.t139 4.428
R1885 VDD.n20 VDD.t160 4.428
R1886 VDD.n21 VDD.t210 4.428
R1887 VDD.n21 VDD.t271 4.428
R1888 VDD.n22 VDD.t150 4.428
R1889 VDD.n22 VDD.t218 4.428
R1890 VDD.n23 VDD.t299 4.428
R1891 VDD.n23 VDD.t197 4.428
R1892 VDD.n24 VDD.t363 4.428
R1893 VDD.n24 VDD.t295 4.428
R1894 VDD.n25 VDD.t27 4.428
R1895 VDD.n25 VDD.t287 4.428
R1896 VDD.n26 VDD.t322 4.428
R1897 VDD.n26 VDD.t355 4.428
R1898 VDD.n27 VDD.t311 4.428
R1899 VDD.n27 VDD.t389 4.428
R1900 VDD.n28 VDD.t373 4.428
R1901 VDD.n28 VDD.t375 4.428
R1902 VDD.n29 VDD.t316 4.428
R1903 VDD.n29 VDD.t339 4.428
R1904 VDD.n30 VDD.t308 4.428
R1905 VDD.n30 VDD.t129 4.428
R1906 VDD.n31 VDD.t257 4.428
R1907 VDD.n31 VDD.t261 4.428
R1908 VDD.n32 VDD.t245 4.428
R1909 VDD.n32 VDD.t337 4.428
R1910 VDD.n33 VDD.t291 4.428
R1911 VDD.n33 VDD.t331 4.428
R1912 VDD.n34 VDD.t359 4.428
R1913 VDD.n34 VDD.t393 4.428
R1914 VDD.n35 VDD.t353 4.428
R1915 VDD.n35 VDD.t281 4.428
R1916 VDD.n36 VDD.t415 4.428
R1917 VDD.n36 VDD.t345 4.428
R1918 VDD.n37 VDD.t409 4.428
R1919 VDD.n37 VDD.t411 4.428
R1920 VDD.n38 VDD.t371 4.428
R1921 VDD.n38 VDD.t407 4.428
R1922 VDD.n39 VDD.t429 4.428
R1923 VDD.n39 VDD.t433 4.428
R1924 VDD.n40 VDD.t301 4.428
R1925 VDD.n40 VDD.t425 4.428
R1926 VDD.n41 VDD.t367 4.428
R1927 VDD.n41 VDD.t251 4.428
R1928 VDD.n987 VDD.t127 4.428
R1929 VDD.n987 VDD.t214 4.428
R1930 VDD.n975 VDD.t183 4.428
R1931 VDD.n975 VDD.t41 4.428
R1932 VDD.n974 VDD.t162 4.428
R1933 VDD.n974 VDD.t437 4.428
R1934 VDD.n973 VDD.t78 4.428
R1935 VDD.n973 VDD.t84 4.428
R1936 VDD.n972 VDD.t51 4.428
R1937 VDD.n972 VDD.t146 4.428
R1938 VDD.n971 VDD.t154 4.428
R1939 VDD.n971 VDD.t199 4.428
R1940 VDD.n970 VDD.t74 4.428
R1941 VDD.n970 VDD.t113 4.428
R1942 VDD.n969 VDD.t67 4.428
R1943 VDD.n969 VDD.t357 4.428
R1944 VDD.n968 VDD.t109 4.428
R1945 VDD.n968 VDD.t421 4.428
R1946 VDD.n967 VDD.t385 4.428
R1947 VDD.n967 VDD.t106 4.428
R1948 VDD.n966 VDD.t33 4.428
R1949 VDD.n966 VDD.t93 4.428
R1950 VDD.n965 VDD.t171 4.428
R1951 VDD.n965 VDD.t231 4.428
R1952 VDD.n929 VDD.t263 4.428
R1953 VDD.n929 VDD.t131 4.428
R1954 VDD.n930 VDD.t247 4.428
R1955 VDD.n930 VDD.t259 4.428
R1956 VDD.n931 VDD.t193 4.428
R1957 VDD.n931 VDD.t195 4.428
R1958 VDD.n932 VDD.t289 4.428
R1959 VDD.n932 VDD.t293 4.428
R1960 VDD.n933 VDD.t62 4.428
R1961 VDD.n933 VDD.t25 4.428
R1962 VDD.n934 VDD.t185 4.428
R1963 VDD.n934 VDD.t187 4.428
R1964 VDD.n935 VDD.t166 4.428
R1965 VDD.n935 VDD.t100 4.428
R1966 VDD.n936 VDD.t224 4.428
R1967 VDD.n936 VDD.t86 4.428
R1968 VDD.n937 VDD.t158 4.428
R1969 VDD.n937 VDD.t220 4.428
R1970 VDD.n938 VDD.t117 4.428
R1971 VDD.n938 VDD.t156 4.428
R1972 VDD.n939 VDD.t253 4.428
R1973 VDD.n939 VDD.t303 4.428
R1974 VDD.n940 VDD.t237 4.428
R1975 VDD.n940 VDD.t369 4.428
R1976 VDD.n941 VDD.t327 4.428
R1977 VDD.n941 VDD.t235 4.428
R1978 VDD.n942 VDD.t391 4.428
R1979 VDD.n942 VDD.t324 4.428
R1980 VDD.n943 VDD.t383 4.428
R1981 VDD.n943 VDD.t273 4.428
R1982 VDD.n944 VDD.t152 4.428
R1983 VDD.n944 VDD.t342 4.428
R1984 VDD.n945 VDD.t137 4.428
R1985 VDD.n945 VDD.t279 4.428
R1986 VDD.n946 VDD.t267 4.428
R1987 VDD.n946 VDD.t269 4.428
R1988 VDD.n75 VDD.n74 4.139
R1989 VDD.n688 sky130_asc_res_xhigh_po_2p85_1_8/VPWR 4.129
R1990 VDD.n590 sky130_asc_res_xhigh_po_2p85_1_0/VPWR 4.129
R1991 sky130_asc_res_xhigh_po_2p85_1_19/VPWR VDD.n863 4.128
R1992 VDD.n878 sky130_asc_cap_mim_m3_1_0/VPWR 4.08
R1993 sky130_asc_res_xhigh_po_2p85_1_11/VPWR sky130_asc_res_xhigh_po_2p85_1_13/VPWR 3.978
R1994 VDD.n252 VDD.n251 3.891
R1995 VDD.n524 sky130_asc_res_xhigh_po_2p85_1_18/VPWR 3.72
R1996 VDD.n377 VDD.n376 3.657
R1997 VDD.n411 VDD.n410 3.657
R1998 VDD.n446 VDD.n445 3.657
R1999 VDD.n480 VDD.n479 3.657
R2000 VDD.n115 VDD.n114 3.657
R2001 VDD.n149 VDD.n148 3.657
R2002 VDD.n183 VDD.n182 3.657
R2003 VDD.n217 VDD.n216 3.657
R2004 VDD.n1024 VDD.n1023 3.657
R2005 VDD.n1058 VDD.n1057 3.657
R2006 VDD.n1093 VDD.n1092 3.657
R2007 VDD.n1127 VDD.n1126 3.657
R2008 sky130_asc_cap_mim_m3_1_3/VPWR VDD.n878 3.648
R2009 VDD.n884 VDD.n883 3.471
R2010 VDD.n877 VDD.n876 3.471
R2011 VDD.n869 VDD.n868 3.471
R2012 sky130_asc_res_xhigh_po_2p85_1_29/VPWR sky130_asc_res_xhigh_po_2p85_2_0/VPWR 3.465
R2013 sky130_asc_res_xhigh_po_2p85_1_27/VPWR sky130_asc_res_xhigh_po_2p85_2_1/VPWR 3.465
R2014 VDD.n882 VDD.n879 3.427
R2015 VDD.n875 VDD.n871 3.427
R2016 VDD.n867 VDD.n864 3.427
R2017 VDD.n881 VDD.n880 3.41
R2018 VDD.n874 VDD.n872 3.41
R2019 VDD.n866 VDD.n865 3.41
R2020 VDD.n1176 sky130_asc_res_xhigh_po_2p85_1_3/VPWR 3.21
R2021 VDD.n1175 sky130_asc_res_xhigh_po_2p85_1_4/VPWR 3.21
R2022 sky130_asc_res_xhigh_po_2p85_1_1/VPWR VDD.n1177 3.2
R2023 VDD.n1173 VDD.n3 3.193
R2024 VDD.n574 sky130_asc_res_xhigh_po_2p85_1_7/VPWR 3.145
R2025 VDD.n76 sky130_asc_cap_mim_m3_1_2/VPWR 3.091
R2026 VDD.n665 VDD.n630 3.04
R2027 VDD.n1160 VDD.n1159 2.974
R2028 VDD.n993 VDD.n990 2.874
R2029 sky130_asc_res_xhigh_po_2p85_1_12/VPWR sky130_asc_res_xhigh_po_2p85_1_14/VPWR 2.855
R2030 sky130_asc_res_xhigh_po_2p85_1_14/VPWR sky130_asc_res_xhigh_po_2p85_1_10/VPWR 2.855
R2031 sky130_asc_res_xhigh_po_2p85_1_10/VPWR sky130_asc_res_xhigh_po_2p85_1_30/VPWR 2.855
R2032 sky130_asc_res_xhigh_po_2p85_1_30/VPWR sky130_asc_res_xhigh_po_2p85_1_29/VPWR 2.855
R2033 sky130_asc_res_xhigh_po_2p85_1_21/VPWR sky130_asc_res_xhigh_po_2p85_1_24/VPWR 2.855
R2034 sky130_asc_res_xhigh_po_2p85_1_24/VPWR sky130_asc_res_xhigh_po_2p85_1_3/VPWR 2.855
R2035 sky130_asc_res_xhigh_po_2p85_1_9/VPWR sky130_asc_res_xhigh_po_2p85_1_2/VPWR 2.855
R2036 sky130_asc_res_xhigh_po_2p85_1_2/VPWR sky130_asc_res_xhigh_po_2p85_1_4/VPWR 2.855
R2037 sky130_asc_res_xhigh_po_2p85_1_6/VPWR sky130_asc_res_xhigh_po_2p85_1_5/VPWR 2.855
R2038 sky130_asc_res_xhigh_po_2p85_1_18/VPWR sky130_asc_res_xhigh_po_2p85_1_20/VPWR 2.855
R2039 sky130_asc_res_xhigh_po_2p85_1_15/VPWR sky130_asc_res_xhigh_po_2p85_1_11/VPWR 2.855
R2040 sky130_asc_res_xhigh_po_2p85_1_13/VPWR sky130_asc_res_xhigh_po_2p85_1_28/VPWR 2.855
R2041 sky130_asc_res_xhigh_po_2p85_1_28/VPWR sky130_asc_res_xhigh_po_2p85_1_26/VPWR 2.855
R2042 sky130_asc_res_xhigh_po_2p85_1_26/VPWR sky130_asc_res_xhigh_po_2p85_1_23/VPWR 2.855
R2043 sky130_asc_res_xhigh_po_2p85_1_23/VPWR sky130_asc_res_xhigh_po_2p85_1_25/VPWR 2.855
R2044 sky130_asc_res_xhigh_po_2p85_1_25/VPWR sky130_asc_res_xhigh_po_2p85_1_27/VPWR 2.855
R2045 sky130_asc_cap_mim_m3_1_8/VPWR sky130_asc_res_xhigh_po_2p85_1_21/VPWR 2.836
R2046 sky130_asc_cap_mim_m3_1_6/VPWR sky130_asc_res_xhigh_po_2p85_1_9/VPWR 2.836
R2047 sky130_asc_cap_mim_m3_1_7/VPWR sky130_asc_res_xhigh_po_2p85_1_6/VPWR 2.836
R2048 VDD.n515 VDD.n512 2.5
R2049 VDD.n78 VDD.n75 2.242
R2050 sky130_asc_cap_mim_m3_1_5/VPWR VDD.n687 2.141
R2051 sky130_asc_cap_mim_m3_1_9/VPWR VDD.n589 2.141
R2052 sky130_asc_nfet_01v8_lvt_9_2/VPWR sky130_asc_pnp_05v5_W3p40L3p40_1_0/VPWR 2.04
R2053 sky130_asc_res_xhigh_po_2p85_1_20/VPWR VDD.n523 2.007
R2054 VDD.n1172 sky130_asc_res_xhigh_po_2p85_1_7/VPWR 1.985
R2055 VDD.n1170 sky130_asc_cap_mim_m3_1_2/VPWR 1.864
R2056 VDD.n573 VDD.n572 1.835
R2057 sky130_asc_pnp_05v5_W3p40L3p40_8_0/VPWR VDD.n737 1.783
R2058 sky130_asc_nfet_01v8_lvt_1_1/VPWR sky130_asc_pnp_05v5_W3p40L3p40_7_0/VPWR 1.766
R2059 VDD.n522 VDD.n284 1.766
R2060 VDD.n1171 VDD.n6 1.458
R2061 VDD.n421 VDD.n346 1.403
R2062 VDD.n84 VDD.n72 1.403
R2063 VDD.n1060 VDD.n988 1.403
R2064 VDD.n878 VDD.n877 1.369
R2065 VDD.n885 VDD.n884 1.368
R2066 VDD.n870 VDD.n869 1.368
R2067 VDD.n1174 sky130_asc_nfet_01v8_lvt_9_0/VPWR 1.25
R2068 VDD.n1168 sky130_asc_nfet_01v8_lvt_1_0/VPWR 1.218
R2069 VDD.n1169 sky130_asc_cap_mim_m3_1_1/VPWR 1.15
R2070 VDD.n284 VDD.n279 1.024
R2071 VDD.n346 VDD.n345 1.023
R2072 VDD.n72 VDD.n71 1.023
R2073 VDD.n988 VDD.n987 1.023
R2074 VDD.t325 sky130_asc_cap_mim_m3_1_2/Cin 0.982
R2075 VDD.t37 sky130_asc_cap_mim_m3_1_1/Cin 0.982
R2076 VDD.t20 sky130_asc_cap_mim_m3_1_3/Cin 0.982
R2077 VDD.t348 sky130_asc_cap_mim_m3_1_0/Cin 0.982
R2078 VDD.t19 sky130_asc_cap_mim_m3_1_4/Cin 0.982
R2079 VDD.n572 VDD.n571 0.958
R2080 VDD.n884 VDD.n879 0.852
R2081 VDD.n877 VDD.n871 0.852
R2082 VDD.n869 VDD.n864 0.852
R2083 VDD.n883 VDD.n882 0.851
R2084 VDD.n876 VDD.n875 0.851
R2085 VDD.n868 VDD.n867 0.851
R2086 sky130_asc_cap_mim_m3_1_4/VPWR sky130_asc_nfet_01v8_lvt_1_0/VPWR 0.849
R2087 VDD.n816 VDD.n0 0.816
R2088 VDD.n1168 VDD.n1167 0.808
R2089 VDD.n1167 VDD.n1166 0.485
R2090 VDD.n1167 VDD.n923 0.485
R2091 VDD.n1167 VDD.n919 0.485
R2092 VDD.n1167 VDD.n904 0.481
R2093 VDD.n1167 VDD.n909 0.481
R2094 VDD.n1167 VDD.n911 0.481
R2095 VDD.n881 VDD.t340 0.447
R2096 VDD.n866 VDD.t36 0.447
R2097 VDD.n512 VDD.n511 0.439
R2098 VDD.n1159 VDD.n1158 0.439
R2099 VDD.n251 VDD.n248 0.439
R2100 VDD.n895 VDD.n892 0.438
R2101 VDD.n687 VDD.n686 0.438
R2102 VDD.n589 VDD.n588 0.438
R2103 VDD.n874 VDD.n873 0.435
R2104 VDD.n870 sky130_asc_nfet_01v8_lvt_1_1/VPWR 0.422
R2105 VDD.n735 VDD.n734 0.416
R2106 VDD.n734 VDD.n722 0.416
R2107 VDD.n729 VDD.n722 0.416
R2108 VDD.n729 VDD.n728 0.416
R2109 VDD.n728 VDD.n727 0.416
R2110 VDD.n686 VDD.n684 0.416
R2111 VDD.n684 VDD.n682 0.416
R2112 VDD.n682 VDD.n680 0.416
R2113 VDD.n680 VDD.n676 0.416
R2114 VDD.n676 VDD.n674 0.416
R2115 VDD.n674 VDD.n672 0.416
R2116 VDD.n667 VDD.n3 0.416
R2117 VDD.n588 VDD.n552 0.416
R2118 VDD.n584 VDD.n552 0.416
R2119 VDD.n584 VDD.n583 0.416
R2120 VDD.n583 VDD.n554 0.416
R2121 VDD.n579 VDD.n554 0.416
R2122 VDD.n579 VDD.n578 0.416
R2123 VDD.n578 VDD.n556 0.416
R2124 VDD.n521 VDD.n517 0.416
R2125 VDD.n517 VDD.n515 0.416
R2126 VDD.n511 VDD.n509 0.416
R2127 VDD.n509 VDD.n507 0.416
R2128 VDD.n507 VDD.n503 0.416
R2129 VDD.n503 VDD.n501 0.416
R2130 VDD.n501 VDD.n499 0.416
R2131 VDD.n499 VDD.n497 0.416
R2132 VDD.n497 VDD.n493 0.416
R2133 VDD.n493 VDD.n491 0.416
R2134 VDD.n491 VDD.n489 0.416
R2135 VDD.n489 VDD.n485 0.416
R2136 VDD.n485 VDD.n483 0.416
R2137 VDD.n483 VDD.n481 0.416
R2138 VDD.n481 VDD.n477 0.416
R2139 VDD.n477 VDD.n475 0.416
R2140 VDD.n475 VDD.n473 0.416
R2141 VDD.n473 VDD.n469 0.416
R2142 VDD.n469 VDD.n467 0.416
R2143 VDD.n467 VDD.n465 0.416
R2144 VDD.n465 VDD.n463 0.416
R2145 VDD.n463 VDD.n459 0.416
R2146 VDD.n459 VDD.n457 0.416
R2147 VDD.n457 VDD.n455 0.416
R2148 VDD.n455 VDD.n451 0.416
R2149 VDD.n451 VDD.n449 0.416
R2150 VDD.n449 VDD.n447 0.416
R2151 VDD.n447 VDD.n443 0.416
R2152 VDD.n443 VDD.n441 0.416
R2153 VDD.n441 VDD.n439 0.416
R2154 VDD.n439 VDD.n435 0.416
R2155 VDD.n435 VDD.n433 0.416
R2156 VDD.n433 VDD.n431 0.416
R2157 VDD.n431 VDD.n429 0.416
R2158 VDD.n429 VDD.n425 0.416
R2159 VDD.n425 VDD.n423 0.416
R2160 VDD.n420 VDD.n416 0.416
R2161 VDD.n416 VDD.n414 0.416
R2162 VDD.n414 VDD.n412 0.416
R2163 VDD.n412 VDD.n408 0.416
R2164 VDD.n408 VDD.n406 0.416
R2165 VDD.n406 VDD.n404 0.416
R2166 VDD.n404 VDD.n400 0.416
R2167 VDD.n400 VDD.n398 0.416
R2168 VDD.n398 VDD.n396 0.416
R2169 VDD.n396 VDD.n394 0.416
R2170 VDD.n394 VDD.n390 0.416
R2171 VDD.n390 VDD.n388 0.416
R2172 VDD.n388 VDD.n386 0.416
R2173 VDD.n386 VDD.n382 0.416
R2174 VDD.n382 VDD.n380 0.416
R2175 VDD.n380 VDD.n378 0.416
R2176 VDD.n378 VDD.n374 0.416
R2177 VDD.n374 VDD.n372 0.416
R2178 VDD.n372 VDD.n370 0.416
R2179 VDD.n370 VDD.n366 0.416
R2180 VDD.n366 VDD.n364 0.416
R2181 VDD.n364 VDD.n362 0.416
R2182 VDD.n362 VDD.n360 0.416
R2183 VDD.n360 VDD.n356 0.416
R2184 VDD.n356 VDD.n354 0.416
R2185 VDD.n354 VDD.n352 0.416
R2186 VDD.n352 VDD.n348 0.416
R2187 VDD.n348 VDD.n6 0.416
R2188 VDD.n248 VDD.n246 0.416
R2189 VDD.n246 VDD.n244 0.416
R2190 VDD.n244 VDD.n240 0.416
R2191 VDD.n240 VDD.n238 0.416
R2192 VDD.n238 VDD.n236 0.416
R2193 VDD.n236 VDD.n234 0.416
R2194 VDD.n234 VDD.n230 0.416
R2195 VDD.n230 VDD.n228 0.416
R2196 VDD.n228 VDD.n226 0.416
R2197 VDD.n226 VDD.n222 0.416
R2198 VDD.n222 VDD.n220 0.416
R2199 VDD.n220 VDD.n218 0.416
R2200 VDD.n218 VDD.n214 0.416
R2201 VDD.n214 VDD.n212 0.416
R2202 VDD.n212 VDD.n210 0.416
R2203 VDD.n210 VDD.n206 0.416
R2204 VDD.n206 VDD.n204 0.416
R2205 VDD.n204 VDD.n202 0.416
R2206 VDD.n202 VDD.n200 0.416
R2207 VDD.n200 VDD.n196 0.416
R2208 VDD.n196 VDD.n194 0.416
R2209 VDD.n194 VDD.n192 0.416
R2210 VDD.n192 VDD.n188 0.416
R2211 VDD.n188 VDD.n186 0.416
R2212 VDD.n186 VDD.n184 0.416
R2213 VDD.n184 VDD.n180 0.416
R2214 VDD.n180 VDD.n178 0.416
R2215 VDD.n178 VDD.n176 0.416
R2216 VDD.n176 VDD.n172 0.416
R2217 VDD.n172 VDD.n170 0.416
R2218 VDD.n170 VDD.n168 0.416
R2219 VDD.n168 VDD.n166 0.416
R2220 VDD.n166 VDD.n162 0.416
R2221 VDD.n162 VDD.n160 0.416
R2222 VDD.n160 VDD.n158 0.416
R2223 VDD.n158 VDD.n154 0.416
R2224 VDD.n154 VDD.n152 0.416
R2225 VDD.n152 VDD.n150 0.416
R2226 VDD.n150 VDD.n146 0.416
R2227 VDD.n146 VDD.n144 0.416
R2228 VDD.n144 VDD.n142 0.416
R2229 VDD.n142 VDD.n138 0.416
R2230 VDD.n138 VDD.n136 0.416
R2231 VDD.n136 VDD.n134 0.416
R2232 VDD.n134 VDD.n132 0.416
R2233 VDD.n132 VDD.n128 0.416
R2234 VDD.n128 VDD.n126 0.416
R2235 VDD.n126 VDD.n124 0.416
R2236 VDD.n124 VDD.n120 0.416
R2237 VDD.n120 VDD.n118 0.416
R2238 VDD.n118 VDD.n116 0.416
R2239 VDD.n116 VDD.n112 0.416
R2240 VDD.n112 VDD.n110 0.416
R2241 VDD.n110 VDD.n108 0.416
R2242 VDD.n108 VDD.n104 0.416
R2243 VDD.n104 VDD.n102 0.416
R2244 VDD.n102 VDD.n100 0.416
R2245 VDD.n100 VDD.n98 0.416
R2246 VDD.n98 VDD.n94 0.416
R2247 VDD.n94 VDD.n92 0.416
R2248 VDD.n92 VDD.n90 0.416
R2249 VDD.n90 VDD.n86 0.416
R2250 VDD.n1158 VDD.n1156 0.416
R2251 VDD.n1156 VDD.n1154 0.416
R2252 VDD.n1154 VDD.n1150 0.416
R2253 VDD.n1150 VDD.n1148 0.416
R2254 VDD.n1148 VDD.n1146 0.416
R2255 VDD.n1146 VDD.n1144 0.416
R2256 VDD.n1144 VDD.n1140 0.416
R2257 VDD.n1140 VDD.n1138 0.416
R2258 VDD.n1138 VDD.n1136 0.416
R2259 VDD.n1136 VDD.n1132 0.416
R2260 VDD.n1132 VDD.n1130 0.416
R2261 VDD.n1130 VDD.n1128 0.416
R2262 VDD.n1128 VDD.n1124 0.416
R2263 VDD.n1124 VDD.n1122 0.416
R2264 VDD.n1122 VDD.n1120 0.416
R2265 VDD.n1120 VDD.n1116 0.416
R2266 VDD.n1116 VDD.n1114 0.416
R2267 VDD.n1114 VDD.n1112 0.416
R2268 VDD.n1112 VDD.n1110 0.416
R2269 VDD.n1110 VDD.n1106 0.416
R2270 VDD.n1106 VDD.n1104 0.416
R2271 VDD.n1104 VDD.n1102 0.416
R2272 VDD.n1102 VDD.n1098 0.416
R2273 VDD.n1098 VDD.n1096 0.416
R2274 VDD.n1096 VDD.n1094 0.416
R2275 VDD.n1094 VDD.n1090 0.416
R2276 VDD.n1090 VDD.n1088 0.416
R2277 VDD.n1088 VDD.n1086 0.416
R2278 VDD.n1086 VDD.n1082 0.416
R2279 VDD.n1082 VDD.n1080 0.416
R2280 VDD.n1080 VDD.n1078 0.416
R2281 VDD.n1078 VDD.n1076 0.416
R2282 VDD.n1076 VDD.n1072 0.416
R2283 VDD.n1072 VDD.n1070 0.416
R2284 VDD.n1070 VDD.n1068 0.416
R2285 VDD.n1068 VDD.n1064 0.416
R2286 VDD.n1064 VDD.n1062 0.416
R2287 VDD.n1059 VDD.n1055 0.416
R2288 VDD.n1055 VDD.n1053 0.416
R2289 VDD.n1053 VDD.n1051 0.416
R2290 VDD.n1051 VDD.n1047 0.416
R2291 VDD.n1047 VDD.n1045 0.416
R2292 VDD.n1045 VDD.n1043 0.416
R2293 VDD.n1043 VDD.n1041 0.416
R2294 VDD.n1041 VDD.n1037 0.416
R2295 VDD.n1037 VDD.n1035 0.416
R2296 VDD.n1035 VDD.n1033 0.416
R2297 VDD.n1033 VDD.n1029 0.416
R2298 VDD.n1029 VDD.n1027 0.416
R2299 VDD.n1027 VDD.n1025 0.416
R2300 VDD.n1025 VDD.n1021 0.416
R2301 VDD.n1021 VDD.n1019 0.416
R2302 VDD.n1019 VDD.n1017 0.416
R2303 VDD.n1017 VDD.n1013 0.416
R2304 VDD.n1013 VDD.n1011 0.416
R2305 VDD.n1011 VDD.n1009 0.416
R2306 VDD.n1009 VDD.n1007 0.416
R2307 VDD.n1007 VDD.n1003 0.416
R2308 VDD.n1003 VDD.n1001 0.416
R2309 VDD.n1001 VDD.n999 0.416
R2310 VDD.n999 VDD.n995 0.416
R2311 VDD.n995 VDD.n993 0.416
R2312 VDD.n1060 VDD.n1059 0.408
R2313 VDD.n77 VDD.n76 0.404
R2314 VDD.n737 VDD.n736 0.389
R2315 VDD.n672 VDD.n668 0.368
R2316 VDD.n668 VDD.n665 0.365
R2317 VDD.n885 sky130_asc_cap_mim_m3_1_3/VPWR 0.362
R2318 VDD.n522 VDD.n521 0.345
R2319 VDD.n84 VDD.n83 0.339
R2320 VDD.n423 VDD.n421 0.3
R2321 VDD.n574 VDD.n573 0.25
R2322 VDD.n573 VDD.n556 0.166
R2323 VDD.n421 VDD.n420 0.116
R2324 VDD.n818 VDD.n815 0.115
R2325 VDD.n821 VDD.n788 0.115
R2326 VDD.n824 VDD.n761 0.115
R2327 VDD.n827 VDD.n711 0.115
R2328 VDD.n830 VDD.n613 0.115
R2329 VDD.n833 VDD.n547 0.115
R2330 VDD.n836 VDD.n275 0.115
R2331 VDD.n840 VDD.n839 0.115
R2332 VDD.n894 VDD.n893 0.106
R2333 VDD.n838 VDD.n837 0.106
R2334 VDD.n835 VDD.n834 0.106
R2335 VDD.n832 VDD.n831 0.106
R2336 VDD.n829 VDD.n828 0.106
R2337 VDD.n826 VDD.n825 0.106
R2338 VDD.n823 VDD.n822 0.106
R2339 VDD.n820 VDD.n819 0.106
R2340 VDD.n817 VDD.n816 0.106
R2341 VDD.n1169 VDD.n1168 0.106
R2342 VDD.n1170 VDD.n1169 0.106
R2343 VDD.n1171 VDD.n1170 0.106
R2344 VDD.n1172 VDD.n1171 0.106
R2345 VDD.n1173 VDD.n1172 0.106
R2346 VDD.n1174 VDD.n1173 0.106
R2347 VDD.n1175 VDD.n1174 0.106
R2348 VDD.n1176 VDD.n1175 0.106
R2349 VDD.n1177 VDD.n1176 0.106
R2350 VDD.n1177 VDD.n0 0.1
R2351 VDD.n523 VDD.n522 0.092
R2352 VDD.n86 VDD.n84 0.077
R2353 VDD.n0 VDD 0.073
R2354 VDD.n668 VDD.n667 0.047
R2355 VDD.n75 VDD.n73 0.041
R2356 VDD.n736 VDD.n735 0.027
R2357 VDD.n1163 VDD.n1162 0.026
R2358 VDD.n843 VDD.n842 0.025
R2359 VDD.n273 VDD.n272 0.025
R2360 VDD.n545 VDD.n544 0.025
R2361 VDD.n611 VDD.n610 0.025
R2362 VDD.n709 VDD.n708 0.025
R2363 VDD.n759 VDD.n758 0.025
R2364 VDD.n786 VDD.n785 0.025
R2365 VDD.n813 VDD.n812 0.025
R2366 VDD.n811 VDD.n810 0.025
R2367 VDD.n784 VDD.n783 0.025
R2368 VDD.n757 VDD.n756 0.025
R2369 VDD.n707 VDD.n706 0.025
R2370 VDD.n609 VDD.n608 0.025
R2371 VDD.n543 VDD.n542 0.025
R2372 VDD.n271 VDD.n270 0.025
R2373 VDD.n845 VDD.n844 0.025
R2374 VDD.n1165 VDD.n1164 0.025
R2375 VDD.n899 VDD.n898 0.025
R2376 VDD.n901 VDD.n900 0.025
R2377 VDD.n914 VDD.n913 0.025
R2378 VDD.t15 VDD.t58 0.025
R2379 VDD.t10 VDD.t15 0.025
R2380 VDD.t334 VDD.t10 0.025
R2381 VDD.t98 VDD.t334 0.025
R2382 VDD.t63 VDD.t56 0.025
R2383 VDD.t56 VDD.t142 0.025
R2384 VDD.t142 VDD.t22 0.025
R2385 VDD.t22 VDD.t325 0.025
R2386 VDD.t340 VDD.t143 0.025
R2387 VDD.t143 VDD.t23 0.025
R2388 VDD.t23 VDD.t88 0.025
R2389 VDD.t88 VDD.t72 0.025
R2390 VDD.t72 VDD.t202 0.025
R2391 VDD.t202 VDD.t124 0.025
R2392 VDD.t124 VDD.t309 0.025
R2393 VDD.t309 VDD.t91 0.025
R2394 VDD.t91 VDD.t37 0.025
R2395 VDD.t144 VDD.t17 0.025
R2396 VDD.t304 VDD.t144 0.025
R2397 VDD.t87 VDD.t304 0.025
R2398 VDD.t265 VDD.t87 0.025
R2399 VDD.t9 VDD.t12 0.025
R2400 VDD.t12 VDD.t264 0.025
R2401 VDD.t264 VDD.t141 0.025
R2402 VDD.t141 VDD.t20 0.025
R2403 VDD.t36 VDD.t229 0.025
R2404 VDD.t229 VDD.t343 0.025
R2405 VDD.t343 VDD.t312 0.025
R2406 VDD.t312 VDD.t107 0.025
R2407 VDD.t107 VDD.t14 0.025
R2408 VDD.t14 VDD.t349 0.025
R2409 VDD.t349 VDD.t57 0.025
R2410 VDD.t57 VDD.t13 0.025
R2411 VDD.t13 VDD.t348 0.025
R2412 VDD.t8 VDD.t18 0.025
R2413 VDD.t11 VDD.t167 0.025
R2414 VDD.t167 VDD.t125 0.025
R2415 VDD.t125 VDD.t16 0.025
R2416 VDD.t16 VDD.t21 0.025
R2417 VDD.t21 VDD.t335 0.025
R2418 VDD.t335 VDD.t140 0.025
R2419 VDD.t140 VDD.t19 0.025
R2420 VDD.n861 VDD.n860 0.023
R2421 VDD.n255 VDD.n254 0.023
R2422 VDD.n527 VDD.n526 0.023
R2423 VDD.n593 VDD.n592 0.023
R2424 VDD.n691 VDD.n690 0.023
R2425 VDD.n741 VDD.n740 0.023
R2426 VDD.n768 VDD.n767 0.023
R2427 VDD.n795 VDD.n794 0.023
R2428 VDD.n797 VDD.n791 0.021
R2429 VDD.n770 VDD.n764 0.021
R2430 VDD.n743 VDD.n714 0.021
R2431 VDD.n693 VDD.n616 0.021
R2432 VDD.n595 VDD.n550 0.021
R2433 VDD.n529 VDD.n278 0.021
R2434 VDD.n257 VDD.n12 0.021
R2435 VDD.n858 VDD.n7 0.021
R2436 VDD.n906 VDD.n905 0.021
R2437 VDD.n901 VDD.n896 0.021
R2438 VDD.n1165 VDD.n926 0.021
R2439 VDD.n892 VDD.n891 0.021
R2440 VDD.n887 VDD.n886 0.021
R2441 VDD.n882 VDD.n881 0.021
R2442 VDD.n875 VDD.n874 0.021
R2443 VDD.n867 VDD.n866 0.021
R2444 VDD.n797 VDD.n796 0.02
R2445 VDD.n770 VDD.n769 0.02
R2446 VDD.n743 VDD.n742 0.02
R2447 VDD.n693 VDD.n692 0.02
R2448 VDD.n595 VDD.n594 0.02
R2449 VDD.n529 VDD.n528 0.02
R2450 VDD.n257 VDD.n256 0.02
R2451 VDD.n859 VDD.n858 0.02
R2452 VDD.n841 VDD.n840 0.019
R2453 VDD.n275 VDD.n274 0.019
R2454 VDD.n547 VDD.n546 0.019
R2455 VDD.n613 VDD.n612 0.019
R2456 VDD.n711 VDD.n710 0.019
R2457 VDD.n761 VDD.n760 0.019
R2458 VDD.n788 VDD.n787 0.019
R2459 VDD.n815 VDD.n814 0.019
R2460 VDD.n904 VDD.n903 0.019
R2461 VDD.n909 VDD.n908 0.019
R2462 VDD.n892 VDD.n890 0.019
R2463 VDD.n79 VDD.n78 0.015
R2464 VDD.n814 VDD.n813 0.014
R2465 VDD.n787 VDD.n786 0.014
R2466 VDD.n760 VDD.n759 0.014
R2467 VDD.n710 VDD.n709 0.014
R2468 VDD.n612 VDD.n611 0.014
R2469 VDD.n546 VDD.n545 0.014
R2470 VDD.n274 VDD.n273 0.014
R2471 VDD.n842 VDD.n841 0.014
R2472 VDD.n890 VDD.n889 0.014
R2473 VDD.n911 VDD.n910 0.014
R2474 VDD.n909 VDD.n906 0.014
R2475 VDD.n904 VDD.n901 0.014
R2476 VDD.n794 VDD.n793 0.013
R2477 VDD.n767 VDD.n766 0.013
R2478 VDD.n740 VDD.n739 0.013
R2479 VDD.n690 VDD.n689 0.013
R2480 VDD.n592 VDD.n591 0.013
R2481 VDD.n526 VDD.n525 0.013
R2482 VDD.n254 VDD.n253 0.013
R2483 VDD.n862 VDD.n861 0.013
R2484 VDD.n74 VDD.t98 0.013
R2485 VDD.n873 VDD.t265 0.013
R2486 VDD.n989 VDD.t8 0.013
R2487 VDD.n809 VDD.n808 0.012
R2488 VDD.n805 VDD.n804 0.012
R2489 VDD.n801 VDD.n800 0.012
R2490 VDD.n782 VDD.n781 0.012
R2491 VDD.n778 VDD.n777 0.012
R2492 VDD.n774 VDD.n773 0.012
R2493 VDD.n755 VDD.n754 0.012
R2494 VDD.n751 VDD.n750 0.012
R2495 VDD.n747 VDD.n746 0.012
R2496 VDD.n705 VDD.n704 0.012
R2497 VDD.n701 VDD.n700 0.012
R2498 VDD.n697 VDD.n696 0.012
R2499 VDD.n607 VDD.n606 0.012
R2500 VDD.n603 VDD.n602 0.012
R2501 VDD.n599 VDD.n598 0.012
R2502 VDD.n541 VDD.n540 0.012
R2503 VDD.n537 VDD.n536 0.012
R2504 VDD.n533 VDD.n532 0.012
R2505 VDD.n269 VDD.n268 0.012
R2506 VDD.n265 VDD.n264 0.012
R2507 VDD.n261 VDD.n260 0.012
R2508 VDD.n847 VDD.n846 0.012
R2509 VDD.n851 VDD.n850 0.012
R2510 VDD.n855 VDD.n854 0.012
R2511 VDD.n889 VDD.n888 0.012
R2512 VDD.n916 VDD.n915 0.012
R2513 VDD.n74 VDD.t63 0.012
R2514 VDD.n873 VDD.t9 0.012
R2515 VDD.n989 VDD.t11 0.012
R2516 VDD.n80 VDD.n79 0.012
R2517 VDD.n857 VDD.n856 0.011
R2518 VDD.n853 VDD.n852 0.011
R2519 VDD.n849 VDD.n848 0.011
R2520 VDD.n259 VDD.n258 0.011
R2521 VDD.n263 VDD.n262 0.011
R2522 VDD.n267 VDD.n266 0.011
R2523 VDD.n531 VDD.n530 0.011
R2524 VDD.n535 VDD.n534 0.011
R2525 VDD.n539 VDD.n538 0.011
R2526 VDD.n597 VDD.n596 0.011
R2527 VDD.n601 VDD.n600 0.011
R2528 VDD.n605 VDD.n604 0.011
R2529 VDD.n695 VDD.n694 0.011
R2530 VDD.n699 VDD.n698 0.011
R2531 VDD.n703 VDD.n702 0.011
R2532 VDD.n745 VDD.n744 0.011
R2533 VDD.n749 VDD.n748 0.011
R2534 VDD.n753 VDD.n752 0.011
R2535 VDD.n772 VDD.n771 0.011
R2536 VDD.n776 VDD.n775 0.011
R2537 VDD.n780 VDD.n779 0.011
R2538 VDD.n799 VDD.n798 0.011
R2539 VDD.n803 VDD.n802 0.011
R2540 VDD.n807 VDD.n806 0.011
R2541 VDD.n1166 VDD.n925 0.011
R2542 VDD.n923 VDD.n921 0.011
R2543 VDD.n919 VDD.n917 0.011
R2544 VDD.n78 VDD.n77 0.011
R2545 VDD.n796 VDD.n795 0.01
R2546 VDD.n769 VDD.n768 0.01
R2547 VDD.n742 VDD.n741 0.01
R2548 VDD.n692 VDD.n691 0.01
R2549 VDD.n594 VDD.n593 0.01
R2550 VDD.n528 VDD.n527 0.01
R2551 VDD.n256 VDD.n255 0.01
R2552 VDD.n860 VDD.n859 0.01
R2553 VDD.n839 VDD.n838 0.009
R2554 VDD.n836 VDD.n835 0.009
R2555 VDD.n833 VDD.n832 0.009
R2556 VDD.n830 VDD.n829 0.009
R2557 VDD.n827 VDD.n826 0.009
R2558 VDD.n824 VDD.n823 0.009
R2559 VDD.n821 VDD.n820 0.009
R2560 VDD.n818 VDD.n817 0.009
R2561 VDD.n806 VDD.n805 0.009
R2562 VDD.n802 VDD.n801 0.009
R2563 VDD.n798 VDD.n797 0.009
R2564 VDD.n779 VDD.n778 0.009
R2565 VDD.n775 VDD.n774 0.009
R2566 VDD.n771 VDD.n770 0.009
R2567 VDD.n752 VDD.n751 0.009
R2568 VDD.n748 VDD.n747 0.009
R2569 VDD.n744 VDD.n743 0.009
R2570 VDD.n702 VDD.n701 0.009
R2571 VDD.n698 VDD.n697 0.009
R2572 VDD.n694 VDD.n693 0.009
R2573 VDD.n604 VDD.n603 0.009
R2574 VDD.n600 VDD.n599 0.009
R2575 VDD.n596 VDD.n595 0.009
R2576 VDD.n538 VDD.n537 0.009
R2577 VDD.n534 VDD.n533 0.009
R2578 VDD.n530 VDD.n529 0.009
R2579 VDD.n266 VDD.n265 0.009
R2580 VDD.n262 VDD.n261 0.009
R2581 VDD.n258 VDD.n257 0.009
R2582 VDD.n850 VDD.n849 0.009
R2583 VDD.n854 VDD.n853 0.009
R2584 VDD.n858 VDD.n857 0.009
R2585 VDD.n919 VDD.n918 0.009
R2586 VDD.n923 VDD.n922 0.009
R2587 VDD.n1166 VDD.n1165 0.009
R2588 VDD.n1062 VDD.n1060 0.008
R2589 VDD.n812 VDD.n811 0.007
R2590 VDD.n810 VDD.n809 0.007
R2591 VDD.n785 VDD.n784 0.007
R2592 VDD.n783 VDD.n782 0.007
R2593 VDD.n758 VDD.n757 0.007
R2594 VDD.n756 VDD.n755 0.007
R2595 VDD.n708 VDD.n707 0.007
R2596 VDD.n706 VDD.n705 0.007
R2597 VDD.n610 VDD.n609 0.007
R2598 VDD.n608 VDD.n607 0.007
R2599 VDD.n544 VDD.n543 0.007
R2600 VDD.n542 VDD.n541 0.007
R2601 VDD.n272 VDD.n271 0.007
R2602 VDD.n270 VDD.n269 0.007
R2603 VDD.n844 VDD.n843 0.007
R2604 VDD.n846 VDD.n845 0.007
R2605 VDD.n900 VDD.n899 0.007
R2606 VDD.n915 VDD.n914 0.007
R2607 VDD.n1164 VDD.n1163 0.007
R2608 VDD.n808 VDD.n807 0.007
R2609 VDD.n804 VDD.n803 0.007
R2610 VDD.n800 VDD.n799 0.007
R2611 VDD.n781 VDD.n780 0.007
R2612 VDD.n777 VDD.n776 0.007
R2613 VDD.n773 VDD.n772 0.007
R2614 VDD.n754 VDD.n753 0.007
R2615 VDD.n750 VDD.n749 0.007
R2616 VDD.n746 VDD.n745 0.007
R2617 VDD.n704 VDD.n703 0.007
R2618 VDD.n700 VDD.n699 0.007
R2619 VDD.n696 VDD.n695 0.007
R2620 VDD.n606 VDD.n605 0.007
R2621 VDD.n602 VDD.n601 0.007
R2622 VDD.n598 VDD.n597 0.007
R2623 VDD.n540 VDD.n539 0.007
R2624 VDD.n536 VDD.n535 0.007
R2625 VDD.n532 VDD.n531 0.007
R2626 VDD.n268 VDD.n267 0.007
R2627 VDD.n264 VDD.n263 0.007
R2628 VDD.n260 VDD.n259 0.007
R2629 VDD.n848 VDD.n847 0.007
R2630 VDD.n852 VDD.n851 0.007
R2631 VDD.n856 VDD.n855 0.007
R2632 VDD.n888 VDD.n887 0.007
R2633 VDD.n908 VDD.n907 0.007
R2634 VDD.n903 VDD.n902 0.007
R2635 VDD.n917 VDD.n916 0.007
R2636 VDD.n921 VDD.n920 0.007
R2637 VDD.n925 VDD.n924 0.007
R2638 VDD.n883 VDD.n880 0.006
R2639 VDD.n876 VDD.n872 0.006
R2640 VDD.n868 VDD.n865 0.006
R2641 VDD.n1162 VDD.n1161 0.006
R2642 VDD.n837 VDD.n836 0.005
R2643 VDD.n834 VDD.n833 0.005
R2644 VDD.n831 VDD.n830 0.005
R2645 VDD.n828 VDD.n827 0.005
R2646 VDD.n825 VDD.n824 0.005
R2647 VDD.n822 VDD.n821 0.005
R2648 VDD.n819 VDD.n818 0.005
R2649 VDD.n880 VDD.n879 0.005
R2650 VDD.n872 VDD.n871 0.005
R2651 VDD.n865 VDD.n864 0.005
R2652 VDD.n895 VDD.n894 0.001
R2653 VDD.n1167 VDD.n895 0.001
R2654 VDD.n811 VDD.n790 0.001
R2655 VDD.n793 VDD.n792 0.001
R2656 VDD.n813 VDD.n789 0.001
R2657 VDD.n784 VDD.n763 0.001
R2658 VDD.n766 VDD.n765 0.001
R2659 VDD.n786 VDD.n762 0.001
R2660 VDD.n757 VDD.n713 0.001
R2661 VDD.n739 VDD.n738 0.001
R2662 VDD.n759 VDD.n712 0.001
R2663 VDD.n707 VDD.n615 0.001
R2664 VDD.n689 VDD.n688 0.001
R2665 VDD.n709 VDD.n614 0.001
R2666 VDD.n609 VDD.n549 0.001
R2667 VDD.n591 VDD.n590 0.001
R2668 VDD.n611 VDD.n548 0.001
R2669 VDD.n543 VDD.n277 0.001
R2670 VDD.n525 VDD.n524 0.001
R2671 VDD.n545 VDD.n276 0.001
R2672 VDD.n271 VDD.n11 0.001
R2673 VDD.n253 VDD.n252 0.001
R2674 VDD.n273 VDD.n10 0.001
R2675 VDD.n844 VDD.n8 0.001
R2676 VDD.n863 VDD.n862 0.001
R2677 VDD.n842 VDD.n9 0.001
R2678 VDD.n913 VDD.n912 0.001
R2679 VDD.n1161 VDD.n1160 0.001
R2680 VDD.n899 VDD.n897 0.001
R2681 VSS.n14750 VSS.n14749 3048.36
R2682 VSS.n12768 VSS.n12736 3048.36
R2683 VSS.n7863 VSS.n7657 3048.36
R2684 VSS.n6853 VSS.n6852 3048.36
R2685 VSS.n4221 VSS.n4189 3048.36
R2686 VSS.n1991 VSS.n1990 3048.36
R2687 VSS.n15971 VSS.n14025 2962.09
R2688 VSS.n12186 VSS.n12074 2962.09
R2689 VSS.n7200 VSS.n6991 2962.09
R2690 VSS.n6877 VSS.n6876 2962.09
R2691 VSS.n5634 VSS.n5633 2962.09
R2692 VSS.n3018 VSS.n3017 2962.09
R2693 VSS.n6828 VSS.n6827 2875.82
R2694 VSS.n6804 VSS.n6803 2760.78
R2695 VSS.n14725 VSS.n14724 2674.51
R2696 VSS.n12795 VSS.n12722 2674.51
R2697 VSS.n7839 VSS.n7838 2674.51
R2698 VSS.n4248 VSS.n4175 2674.51
R2699 VSS.n1966 VSS.n1965 2674.51
R2700 VSS.n15953 VSS.n14037 2588.24
R2701 VSS.n15954 VSS.n15953 2588.24
R2702 VSS.n15955 VSS.n15954 2588.24
R2703 VSS.n15955 VSS.n14033 2588.24
R2704 VSS.n15961 VSS.n14033 2588.24
R2705 VSS.n15962 VSS.n15961 2588.24
R2706 VSS.n15963 VSS.n15962 2588.24
R2707 VSS.n15963 VSS.n14029 2588.24
R2708 VSS.n15969 VSS.n14029 2588.24
R2709 VSS.n15970 VSS.n15969 2588.24
R2710 VSS.n15971 VSS.n15970 2588.24
R2711 VSS.n15995 VSS.n15994 2588.24
R2712 VSS.n15994 VSS.n15993 2588.24
R2713 VSS.n15993 VSS.n14017 2588.24
R2714 VSS.n15987 VSS.n14017 2588.24
R2715 VSS.n15987 VSS.n15986 2588.24
R2716 VSS.n15986 VSS.n15985 2588.24
R2717 VSS.n15985 VSS.n14021 2588.24
R2718 VSS.n15979 VSS.n14021 2588.24
R2719 VSS.n15979 VSS.n15978 2588.24
R2720 VSS.n15978 VSS.n15977 2588.24
R2721 VSS.n15977 VSS.n14025 2588.24
R2722 VSS.n15920 VSS.n14052 2588.24
R2723 VSS.n15926 VSS.n14052 2588.24
R2724 VSS.n15927 VSS.n15926 2588.24
R2725 VSS.n15928 VSS.n15927 2588.24
R2726 VSS.n15928 VSS.n14048 2588.24
R2727 VSS.n15934 VSS.n14048 2588.24
R2728 VSS.n15935 VSS.n15934 2588.24
R2729 VSS.n15937 VSS.n15935 2588.24
R2730 VSS.n15937 VSS.n15936 2588.24
R2731 VSS.n15936 VSS.n14044 2588.24
R2732 VSS.n15944 VSS.n14044 2588.24
R2733 VSS.n14193 VSS.n14159 2588.24
R2734 VSS.n14187 VSS.n14159 2588.24
R2735 VSS.n14187 VSS.n14186 2588.24
R2736 VSS.n14186 VSS.n14185 2588.24
R2737 VSS.n14185 VSS.n14163 2588.24
R2738 VSS.n14179 VSS.n14163 2588.24
R2739 VSS.n14179 VSS.n14178 2588.24
R2740 VSS.n14178 VSS.n14177 2588.24
R2741 VSS.n14177 VSS.n14167 2588.24
R2742 VSS.n14171 VSS.n14167 2588.24
R2743 VSS.n14171 VSS.n14056 2588.24
R2744 VSS.n15391 VSS.n15390 2588.24
R2745 VSS.n15391 VSS.n14202 2588.24
R2746 VSS.n15397 VSS.n14202 2588.24
R2747 VSS.n15398 VSS.n15397 2588.24
R2748 VSS.n15399 VSS.n15398 2588.24
R2749 VSS.n15399 VSS.n14198 2588.24
R2750 VSS.n15405 VSS.n14198 2588.24
R2751 VSS.n15406 VSS.n15405 2588.24
R2752 VSS.n15407 VSS.n15406 2588.24
R2753 VSS.n15407 VSS.n14194 2588.24
R2754 VSS.n15413 VSS.n14194 2588.24
R2755 VSS.n15363 VSS.n15362 2588.24
R2756 VSS.n15364 VSS.n15363 2588.24
R2757 VSS.n15364 VSS.n14217 2588.24
R2758 VSS.n15370 VSS.n14217 2588.24
R2759 VSS.n15371 VSS.n15370 2588.24
R2760 VSS.n15372 VSS.n15371 2588.24
R2761 VSS.n15372 VSS.n14213 2588.24
R2762 VSS.n15379 VSS.n14213 2588.24
R2763 VSS.n15380 VSS.n15379 2588.24
R2764 VSS.n15381 VSS.n15380 2588.24
R2765 VSS.n15381 VSS.n14206 2588.24
R2766 VSS.n14834 VSS.n14801 2588.24
R2767 VSS.n14805 VSS.n14801 2588.24
R2768 VSS.n14827 VSS.n14805 2588.24
R2769 VSS.n14827 VSS.n14826 2588.24
R2770 VSS.n14826 VSS.n14825 2588.24
R2771 VSS.n14825 VSS.n14806 2588.24
R2772 VSS.n14819 VSS.n14806 2588.24
R2773 VSS.n14819 VSS.n14818 2588.24
R2774 VSS.n14818 VSS.n14817 2588.24
R2775 VSS.n14817 VSS.n14810 2588.24
R2776 VSS.n14811 VSS.n14810 2588.24
R2777 VSS.n14783 VSS.n14333 2588.24
R2778 VSS.n14784 VSS.n14783 2588.24
R2779 VSS.n14785 VSS.n14784 2588.24
R2780 VSS.n14785 VSS.n14329 2588.24
R2781 VSS.n14791 VSS.n14329 2588.24
R2782 VSS.n14792 VSS.n14791 2588.24
R2783 VSS.n14793 VSS.n14792 2588.24
R2784 VSS.n14793 VSS.n14325 2588.24
R2785 VSS.n14799 VSS.n14325 2588.24
R2786 VSS.n14800 VSS.n14799 2588.24
R2787 VSS.n14836 VSS.n14800 2588.24
R2788 VSS.n14750 VSS.n14348 2588.24
R2789 VSS.n14756 VSS.n14348 2588.24
R2790 VSS.n14757 VSS.n14756 2588.24
R2791 VSS.n14758 VSS.n14757 2588.24
R2792 VSS.n14758 VSS.n14344 2588.24
R2793 VSS.n14764 VSS.n14344 2588.24
R2794 VSS.n14765 VSS.n14764 2588.24
R2795 VSS.n14767 VSS.n14765 2588.24
R2796 VSS.n14767 VSS.n14766 2588.24
R2797 VSS.n14766 VSS.n14340 2588.24
R2798 VSS.n14774 VSS.n14340 2588.24
R2799 VSS.n14726 VSS.n14360 2588.24
R2800 VSS.n14732 VSS.n14360 2588.24
R2801 VSS.n14733 VSS.n14732 2588.24
R2802 VSS.n14734 VSS.n14733 2588.24
R2803 VSS.n14734 VSS.n14356 2588.24
R2804 VSS.n14740 VSS.n14356 2588.24
R2805 VSS.n14741 VSS.n14740 2588.24
R2806 VSS.n14742 VSS.n14741 2588.24
R2807 VSS.n14742 VSS.n14352 2588.24
R2808 VSS.n14748 VSS.n14352 2588.24
R2809 VSS.n14749 VSS.n14748 2588.24
R2810 VSS.n12168 VSS.n12086 2588.24
R2811 VSS.n12169 VSS.n12168 2588.24
R2812 VSS.n12170 VSS.n12169 2588.24
R2813 VSS.n12170 VSS.n12082 2588.24
R2814 VSS.n12176 VSS.n12082 2588.24
R2815 VSS.n12177 VSS.n12176 2588.24
R2816 VSS.n12178 VSS.n12177 2588.24
R2817 VSS.n12178 VSS.n12078 2588.24
R2818 VSS.n12184 VSS.n12078 2588.24
R2819 VSS.n12185 VSS.n12184 2588.24
R2820 VSS.n12186 VSS.n12185 2588.24
R2821 VSS.n12210 VSS.n12209 2588.24
R2822 VSS.n12209 VSS.n12208 2588.24
R2823 VSS.n12208 VSS.n12066 2588.24
R2824 VSS.n12202 VSS.n12066 2588.24
R2825 VSS.n12202 VSS.n12201 2588.24
R2826 VSS.n12201 VSS.n12200 2588.24
R2827 VSS.n12200 VSS.n12070 2588.24
R2828 VSS.n12194 VSS.n12070 2588.24
R2829 VSS.n12194 VSS.n12193 2588.24
R2830 VSS.n12193 VSS.n12192 2588.24
R2831 VSS.n12192 VSS.n12074 2588.24
R2832 VSS.n12135 VSS.n12134 2588.24
R2833 VSS.n12141 VSS.n12134 2588.24
R2834 VSS.n12142 VSS.n12141 2588.24
R2835 VSS.n12143 VSS.n12142 2588.24
R2836 VSS.n12143 VSS.n12130 2588.24
R2837 VSS.n12149 VSS.n12130 2588.24
R2838 VSS.n12150 VSS.n12149 2588.24
R2839 VSS.n12152 VSS.n12150 2588.24
R2840 VSS.n12152 VSS.n12151 2588.24
R2841 VSS.n12151 VSS.n12126 2588.24
R2842 VSS.n12159 VSS.n12126 2588.24
R2843 VSS.n12455 VSS.n11510 2588.24
R2844 VSS.n12455 VSS.n12454 2588.24
R2845 VSS.n12454 VSS.n12453 2588.24
R2846 VSS.n12453 VSS.n11517 2588.24
R2847 VSS.n12447 VSS.n11517 2588.24
R2848 VSS.n12447 VSS.n12446 2588.24
R2849 VSS.n12446 VSS.n12445 2588.24
R2850 VSS.n12445 VSS.n11522 2588.24
R2851 VSS.n12439 VSS.n11522 2588.24
R2852 VSS.n12439 VSS.n12438 2588.24
R2853 VSS.n12438 VSS.n12437 2588.24
R2854 VSS.n12487 VSS.n11498 2588.24
R2855 VSS.n12481 VSS.n11498 2588.24
R2856 VSS.n12481 VSS.n12480 2588.24
R2857 VSS.n12480 VSS.n12479 2588.24
R2858 VSS.n12479 VSS.n11502 2588.24
R2859 VSS.n12473 VSS.n11502 2588.24
R2860 VSS.n12473 VSS.n12472 2588.24
R2861 VSS.n12472 VSS.n12471 2588.24
R2862 VSS.n12471 VSS.n11506 2588.24
R2863 VSS.n12465 VSS.n11506 2588.24
R2864 VSS.n12465 VSS.n12464 2588.24
R2865 VSS.n13347 VSS.n13346 2588.24
R2866 VSS.n13347 VSS.n12496 2588.24
R2867 VSS.n13353 VSS.n12496 2588.24
R2868 VSS.n13354 VSS.n13353 2588.24
R2869 VSS.n13355 VSS.n13354 2588.24
R2870 VSS.n13355 VSS.n12492 2588.24
R2871 VSS.n13361 VSS.n12492 2588.24
R2872 VSS.n13362 VSS.n13361 2588.24
R2873 VSS.n13363 VSS.n13362 2588.24
R2874 VSS.n13363 VSS.n12488 2588.24
R2875 VSS.n13369 VSS.n12488 2588.24
R2876 VSS.n12628 VSS.n12599 2588.24
R2877 VSS.n12622 VSS.n12599 2588.24
R2878 VSS.n12622 VSS.n12621 2588.24
R2879 VSS.n12621 VSS.n12620 2588.24
R2880 VSS.n12620 VSS.n12603 2588.24
R2881 VSS.n12614 VSS.n12603 2588.24
R2882 VSS.n12614 VSS.n12613 2588.24
R2883 VSS.n12613 VSS.n12612 2588.24
R2884 VSS.n12612 VSS.n12607 2588.24
R2885 VSS.n12607 VSS.n12501 2588.24
R2886 VSS.n13344 VSS.n12501 2588.24
R2887 VSS.n13098 VSS.n13097 2588.24
R2888 VSS.n13098 VSS.n12637 2588.24
R2889 VSS.n13104 VSS.n12637 2588.24
R2890 VSS.n13105 VSS.n13104 2588.24
R2891 VSS.n13106 VSS.n13105 2588.24
R2892 VSS.n13106 VSS.n12633 2588.24
R2893 VSS.n13112 VSS.n12633 2588.24
R2894 VSS.n13113 VSS.n13112 2588.24
R2895 VSS.n13114 VSS.n13113 2588.24
R2896 VSS.n13114 VSS.n12629 2588.24
R2897 VSS.n13120 VSS.n12629 2588.24
R2898 VSS.n12762 VSS.n12736 2588.24
R2899 VSS.n12762 VSS.n12761 2588.24
R2900 VSS.n12761 VSS.n12760 2588.24
R2901 VSS.n12760 VSS.n12740 2588.24
R2902 VSS.n12754 VSS.n12740 2588.24
R2903 VSS.n12754 VSS.n12753 2588.24
R2904 VSS.n12753 VSS.n12752 2588.24
R2905 VSS.n12752 VSS.n12744 2588.24
R2906 VSS.n12746 VSS.n12744 2588.24
R2907 VSS.n12746 VSS.n12642 2588.24
R2908 VSS.n13095 VSS.n12642 2588.24
R2909 VSS.n12786 VSS.n12725 2588.24
R2910 VSS.n12786 VSS.n12785 2588.24
R2911 VSS.n12785 VSS.n12784 2588.24
R2912 VSS.n12784 VSS.n12727 2588.24
R2913 VSS.n12778 VSS.n12727 2588.24
R2914 VSS.n12778 VSS.n12777 2588.24
R2915 VSS.n12777 VSS.n12776 2588.24
R2916 VSS.n12776 VSS.n12732 2588.24
R2917 VSS.n12770 VSS.n12732 2588.24
R2918 VSS.n12770 VSS.n12769 2588.24
R2919 VSS.n12769 VSS.n12768 2588.24
R2920 VSS.n7224 VSS.n7223 2588.24
R2921 VSS.n7223 VSS.n7222 2588.24
R2922 VSS.n7222 VSS.n6983 2588.24
R2923 VSS.n7216 VSS.n6983 2588.24
R2924 VSS.n7216 VSS.n7215 2588.24
R2925 VSS.n7215 VSS.n7214 2588.24
R2926 VSS.n7214 VSS.n6987 2588.24
R2927 VSS.n7208 VSS.n6987 2588.24
R2928 VSS.n7208 VSS.n7207 2588.24
R2929 VSS.n7207 VSS.n7206 2588.24
R2930 VSS.n7206 VSS.n6991 2588.24
R2931 VSS.n7182 VSS.n7003 2588.24
R2932 VSS.n7183 VSS.n7182 2588.24
R2933 VSS.n7184 VSS.n7183 2588.24
R2934 VSS.n7184 VSS.n6999 2588.24
R2935 VSS.n7190 VSS.n6999 2588.24
R2936 VSS.n7191 VSS.n7190 2588.24
R2937 VSS.n7192 VSS.n7191 2588.24
R2938 VSS.n7192 VSS.n6995 2588.24
R2939 VSS.n7198 VSS.n6995 2588.24
R2940 VSS.n7199 VSS.n7198 2588.24
R2941 VSS.n7200 VSS.n7199 2588.24
R2942 VSS.n8807 VSS.n7237 2588.24
R2943 VSS.n8808 VSS.n8807 2588.24
R2944 VSS.n8809 VSS.n8808 2588.24
R2945 VSS.n8809 VSS.n7233 2588.24
R2946 VSS.n8815 VSS.n7233 2588.24
R2947 VSS.n8816 VSS.n8815 2588.24
R2948 VSS.n8817 VSS.n8816 2588.24
R2949 VSS.n8817 VSS.n7229 2588.24
R2950 VSS.n8823 VSS.n7229 2588.24
R2951 VSS.n8824 VSS.n8823 2588.24
R2952 VSS.n8825 VSS.n8824 2588.24
R2953 VSS.n7364 VSS.n7363 2588.24
R2954 VSS.n7363 VSS.n7362 2588.24
R2955 VSS.n7362 VSS.n7339 2588.24
R2956 VSS.n7356 VSS.n7339 2588.24
R2957 VSS.n7356 VSS.n7355 2588.24
R2958 VSS.n7355 VSS.n7354 2588.24
R2959 VSS.n7354 VSS.n7343 2588.24
R2960 VSS.n7348 VSS.n7343 2588.24
R2961 VSS.n7348 VSS.n7347 2588.24
R2962 VSS.n7347 VSS.n7243 2588.24
R2963 VSS.n8800 VSS.n7243 2588.24
R2964 VSS.n8585 VSS.n7377 2588.24
R2965 VSS.n8586 VSS.n8585 2588.24
R2966 VSS.n8587 VSS.n8586 2588.24
R2967 VSS.n8587 VSS.n7373 2588.24
R2968 VSS.n8593 VSS.n7373 2588.24
R2969 VSS.n8594 VSS.n8593 2588.24
R2970 VSS.n8595 VSS.n8594 2588.24
R2971 VSS.n8595 VSS.n7369 2588.24
R2972 VSS.n8601 VSS.n7369 2588.24
R2973 VSS.n8602 VSS.n8601 2588.24
R2974 VSS.n8603 VSS.n8602 2588.24
R2975 VSS.n7504 VSS.n7503 2588.24
R2976 VSS.n7503 VSS.n7502 2588.24
R2977 VSS.n7502 VSS.n7479 2588.24
R2978 VSS.n7496 VSS.n7479 2588.24
R2979 VSS.n7496 VSS.n7495 2588.24
R2980 VSS.n7495 VSS.n7494 2588.24
R2981 VSS.n7494 VSS.n7483 2588.24
R2982 VSS.n7488 VSS.n7483 2588.24
R2983 VSS.n7488 VSS.n7487 2588.24
R2984 VSS.n7487 VSS.n7383 2588.24
R2985 VSS.n8578 VSS.n7383 2588.24
R2986 VSS.n8227 VSS.n7517 2588.24
R2987 VSS.n8228 VSS.n8227 2588.24
R2988 VSS.n8229 VSS.n8228 2588.24
R2989 VSS.n8229 VSS.n7513 2588.24
R2990 VSS.n8235 VSS.n7513 2588.24
R2991 VSS.n8236 VSS.n8235 2588.24
R2992 VSS.n8237 VSS.n8236 2588.24
R2993 VSS.n8237 VSS.n7509 2588.24
R2994 VSS.n8243 VSS.n7509 2588.24
R2995 VSS.n8244 VSS.n8243 2588.24
R2996 VSS.n8245 VSS.n8244 2588.24
R2997 VSS.n7644 VSS.n7643 2588.24
R2998 VSS.n7643 VSS.n7642 2588.24
R2999 VSS.n7642 VSS.n7619 2588.24
R3000 VSS.n7636 VSS.n7619 2588.24
R3001 VSS.n7636 VSS.n7635 2588.24
R3002 VSS.n7635 VSS.n7634 2588.24
R3003 VSS.n7634 VSS.n7623 2588.24
R3004 VSS.n7628 VSS.n7623 2588.24
R3005 VSS.n7628 VSS.n7627 2588.24
R3006 VSS.n7627 VSS.n7523 2588.24
R3007 VSS.n8220 VSS.n7523 2588.24
R3008 VSS.n7869 VSS.n7657 2588.24
R3009 VSS.n7870 VSS.n7869 2588.24
R3010 VSS.n7871 VSS.n7870 2588.24
R3011 VSS.n7871 VSS.n7653 2588.24
R3012 VSS.n7877 VSS.n7653 2588.24
R3013 VSS.n7878 VSS.n7877 2588.24
R3014 VSS.n7879 VSS.n7878 2588.24
R3015 VSS.n7879 VSS.n7649 2588.24
R3016 VSS.n7885 VSS.n7649 2588.24
R3017 VSS.n7886 VSS.n7885 2588.24
R3018 VSS.n7887 VSS.n7886 2588.24
R3019 VSS.n7845 VSS.n7669 2588.24
R3020 VSS.n7846 VSS.n7845 2588.24
R3021 VSS.n7847 VSS.n7846 2588.24
R3022 VSS.n7847 VSS.n7665 2588.24
R3023 VSS.n7853 VSS.n7665 2588.24
R3024 VSS.n7854 VSS.n7853 2588.24
R3025 VSS.n7855 VSS.n7854 2588.24
R3026 VSS.n7855 VSS.n7661 2588.24
R3027 VSS.n7861 VSS.n7661 2588.24
R3028 VSS.n7862 VSS.n7861 2588.24
R3029 VSS.n7863 VSS.n7862 2588.24
R3030 VSS.n6827 VSS.n6759 2588.24
R3031 VSS.n6821 VSS.n6759 2588.24
R3032 VSS.n6821 VSS.n6820 2588.24
R3033 VSS.n6820 VSS.n6819 2588.24
R3034 VSS.n6819 VSS.n6763 2588.24
R3035 VSS.n6813 VSS.n6763 2588.24
R3036 VSS.n6813 VSS.n6812 2588.24
R3037 VSS.n6812 VSS.n6811 2588.24
R3038 VSS.n6811 VSS.n6766 2588.24
R3039 VSS.n6805 VSS.n6766 2588.24
R3040 VSS.n6805 VSS.n6804 2588.24
R3041 VSS.n6797 VSS.n6771 2588.24
R3042 VSS.n6797 VSS.n6796 2588.24
R3043 VSS.n6796 VSS.n6795 2588.24
R3044 VSS.n6795 VSS.n6775 2588.24
R3045 VSS.n6789 VSS.n6775 2588.24
R3046 VSS.n6789 VSS.n6788 2588.24
R3047 VSS.n6788 VSS.n6787 2588.24
R3048 VSS.n6787 VSS.n6779 2588.24
R3049 VSS.n6781 VSS.n6779 2588.24
R3050 VSS.n6781 VSS.n6733 2588.24
R3051 VSS.n6877 VSS.n6733 2588.24
R3052 VSS.n6853 VSS.n6742 2588.24
R3053 VSS.n6859 VSS.n6742 2588.24
R3054 VSS.n6860 VSS.n6859 2588.24
R3055 VSS.n6861 VSS.n6860 2588.24
R3056 VSS.n6861 VSS.n6738 2588.24
R3057 VSS.n6867 VSS.n6738 2588.24
R3058 VSS.n6868 VSS.n6867 2588.24
R3059 VSS.n6869 VSS.n6868 2588.24
R3060 VSS.n6869 VSS.n6734 2588.24
R3061 VSS.n6875 VSS.n6734 2588.24
R3062 VSS.n6876 VSS.n6875 2588.24
R3063 VSS.n6829 VSS.n6754 2588.24
R3064 VSS.n6835 VSS.n6754 2588.24
R3065 VSS.n6836 VSS.n6835 2588.24
R3066 VSS.n6837 VSS.n6836 2588.24
R3067 VSS.n6837 VSS.n6750 2588.24
R3068 VSS.n6843 VSS.n6750 2588.24
R3069 VSS.n6844 VSS.n6843 2588.24
R3070 VSS.n6845 VSS.n6844 2588.24
R3071 VSS.n6845 VSS.n6746 2588.24
R3072 VSS.n6851 VSS.n6746 2588.24
R3073 VSS.n6852 VSS.n6851 2588.24
R3074 VSS.n5611 VSS.n5610 2588.24
R3075 VSS.n5611 VSS.n3667 2588.24
R3076 VSS.n5617 VSS.n3667 2588.24
R3077 VSS.n5618 VSS.n5617 2588.24
R3078 VSS.n5619 VSS.n5618 2588.24
R3079 VSS.n5619 VSS.n3663 2588.24
R3080 VSS.n5625 VSS.n3663 2588.24
R3081 VSS.n5626 VSS.n5625 2588.24
R3082 VSS.n5627 VSS.n5626 2588.24
R3083 VSS.n5627 VSS.n3659 2588.24
R3084 VSS.n5633 VSS.n3659 2588.24
R3085 VSS.n5657 VSS.n3642 2588.24
R3086 VSS.n5651 VSS.n3642 2588.24
R3087 VSS.n5651 VSS.n5650 2588.24
R3088 VSS.n5650 VSS.n5649 2588.24
R3089 VSS.n5649 VSS.n3651 2588.24
R3090 VSS.n5643 VSS.n3651 2588.24
R3091 VSS.n5643 VSS.n5642 2588.24
R3092 VSS.n5642 VSS.n5641 2588.24
R3093 VSS.n5641 VSS.n3655 2588.24
R3094 VSS.n5635 VSS.n3655 2588.24
R3095 VSS.n5635 VSS.n5634 2588.24
R3096 VSS.n3799 VSS.n3770 2588.24
R3097 VSS.n3793 VSS.n3770 2588.24
R3098 VSS.n3793 VSS.n3792 2588.24
R3099 VSS.n3792 VSS.n3791 2588.24
R3100 VSS.n3791 VSS.n3774 2588.24
R3101 VSS.n3785 VSS.n3774 2588.24
R3102 VSS.n3785 VSS.n3784 2588.24
R3103 VSS.n3784 VSS.n3783 2588.24
R3104 VSS.n3783 VSS.n3778 2588.24
R3105 VSS.n3778 VSS.n3672 2588.24
R3106 VSS.n5608 VSS.n3672 2588.24
R3107 VSS.n5265 VSS.n5264 2588.24
R3108 VSS.n5265 VSS.n3808 2588.24
R3109 VSS.n5271 VSS.n3808 2588.24
R3110 VSS.n5272 VSS.n5271 2588.24
R3111 VSS.n5273 VSS.n5272 2588.24
R3112 VSS.n5273 VSS.n3804 2588.24
R3113 VSS.n5279 VSS.n3804 2588.24
R3114 VSS.n5280 VSS.n5279 2588.24
R3115 VSS.n5281 VSS.n5280 2588.24
R3116 VSS.n5281 VSS.n3800 2588.24
R3117 VSS.n5287 VSS.n3800 2588.24
R3118 VSS.n3940 VSS.n3911 2588.24
R3119 VSS.n3934 VSS.n3911 2588.24
R3120 VSS.n3934 VSS.n3933 2588.24
R3121 VSS.n3933 VSS.n3932 2588.24
R3122 VSS.n3932 VSS.n3915 2588.24
R3123 VSS.n3926 VSS.n3915 2588.24
R3124 VSS.n3926 VSS.n3925 2588.24
R3125 VSS.n3925 VSS.n3924 2588.24
R3126 VSS.n3924 VSS.n3919 2588.24
R3127 VSS.n3919 VSS.n3813 2588.24
R3128 VSS.n5262 VSS.n3813 2588.24
R3129 VSS.n4908 VSS.n4907 2588.24
R3130 VSS.n4908 VSS.n3949 2588.24
R3131 VSS.n4914 VSS.n3949 2588.24
R3132 VSS.n4915 VSS.n4914 2588.24
R3133 VSS.n4916 VSS.n4915 2588.24
R3134 VSS.n4916 VSS.n3945 2588.24
R3135 VSS.n4922 VSS.n3945 2588.24
R3136 VSS.n4923 VSS.n4922 2588.24
R3137 VSS.n4924 VSS.n4923 2588.24
R3138 VSS.n4924 VSS.n3941 2588.24
R3139 VSS.n4930 VSS.n3941 2588.24
R3140 VSS.n4081 VSS.n4052 2588.24
R3141 VSS.n4075 VSS.n4052 2588.24
R3142 VSS.n4075 VSS.n4074 2588.24
R3143 VSS.n4074 VSS.n4073 2588.24
R3144 VSS.n4073 VSS.n4056 2588.24
R3145 VSS.n4067 VSS.n4056 2588.24
R3146 VSS.n4067 VSS.n4066 2588.24
R3147 VSS.n4066 VSS.n4065 2588.24
R3148 VSS.n4065 VSS.n4060 2588.24
R3149 VSS.n4060 VSS.n3954 2588.24
R3150 VSS.n4905 VSS.n3954 2588.24
R3151 VSS.n4551 VSS.n4550 2588.24
R3152 VSS.n4551 VSS.n4090 2588.24
R3153 VSS.n4557 VSS.n4090 2588.24
R3154 VSS.n4558 VSS.n4557 2588.24
R3155 VSS.n4559 VSS.n4558 2588.24
R3156 VSS.n4559 VSS.n4086 2588.24
R3157 VSS.n4565 VSS.n4086 2588.24
R3158 VSS.n4566 VSS.n4565 2588.24
R3159 VSS.n4567 VSS.n4566 2588.24
R3160 VSS.n4567 VSS.n4082 2588.24
R3161 VSS.n4573 VSS.n4082 2588.24
R3162 VSS.n4215 VSS.n4189 2588.24
R3163 VSS.n4215 VSS.n4214 2588.24
R3164 VSS.n4214 VSS.n4213 2588.24
R3165 VSS.n4213 VSS.n4193 2588.24
R3166 VSS.n4207 VSS.n4193 2588.24
R3167 VSS.n4207 VSS.n4206 2588.24
R3168 VSS.n4206 VSS.n4205 2588.24
R3169 VSS.n4205 VSS.n4197 2588.24
R3170 VSS.n4199 VSS.n4197 2588.24
R3171 VSS.n4199 VSS.n4095 2588.24
R3172 VSS.n4548 VSS.n4095 2588.24
R3173 VSS.n4239 VSS.n4178 2588.24
R3174 VSS.n4239 VSS.n4238 2588.24
R3175 VSS.n4238 VSS.n4237 2588.24
R3176 VSS.n4237 VSS.n4180 2588.24
R3177 VSS.n4231 VSS.n4180 2588.24
R3178 VSS.n4231 VSS.n4230 2588.24
R3179 VSS.n4230 VSS.n4229 2588.24
R3180 VSS.n4229 VSS.n4185 2588.24
R3181 VSS.n4223 VSS.n4185 2588.24
R3182 VSS.n4223 VSS.n4222 2588.24
R3183 VSS.n4222 VSS.n4221 2588.24
R3184 VSS.n3041 VSS.n3040 2588.24
R3185 VSS.n3040 VSS.n1273 2588.24
R3186 VSS.n3034 VSS.n1273 2588.24
R3187 VSS.n3034 VSS.n3033 2588.24
R3188 VSS.n3033 VSS.n3032 2588.24
R3189 VSS.n3032 VSS.n1277 2588.24
R3190 VSS.n3026 VSS.n1277 2588.24
R3191 VSS.n3026 VSS.n3025 2588.24
R3192 VSS.n3025 VSS.n3024 2588.24
R3193 VSS.n3024 VSS.n1281 2588.24
R3194 VSS.n3018 VSS.n1281 2588.24
R3195 VSS.n2994 VSS.n1293 2588.24
R3196 VSS.n3000 VSS.n1293 2588.24
R3197 VSS.n3001 VSS.n3000 2588.24
R3198 VSS.n3002 VSS.n3001 2588.24
R3199 VSS.n3002 VSS.n1289 2588.24
R3200 VSS.n3008 VSS.n1289 2588.24
R3201 VSS.n3009 VSS.n3008 2588.24
R3202 VSS.n3010 VSS.n3009 2588.24
R3203 VSS.n3010 VSS.n1285 2588.24
R3204 VSS.n3016 VSS.n1285 2588.24
R3205 VSS.n3017 VSS.n3016 2588.24
R3206 VSS.n1434 VSS.n1400 2588.24
R3207 VSS.n1428 VSS.n1400 2588.24
R3208 VSS.n1428 VSS.n1427 2588.24
R3209 VSS.n1427 VSS.n1426 2588.24
R3210 VSS.n1426 VSS.n1404 2588.24
R3211 VSS.n1420 VSS.n1404 2588.24
R3212 VSS.n1420 VSS.n1419 2588.24
R3213 VSS.n1419 VSS.n1418 2588.24
R3214 VSS.n1418 VSS.n1408 2588.24
R3215 VSS.n1412 VSS.n1408 2588.24
R3216 VSS.n1412 VSS.n1297 2588.24
R3217 VSS.n2632 VSS.n2631 2588.24
R3218 VSS.n2632 VSS.n1443 2588.24
R3219 VSS.n2638 VSS.n1443 2588.24
R3220 VSS.n2639 VSS.n2638 2588.24
R3221 VSS.n2640 VSS.n2639 2588.24
R3222 VSS.n2640 VSS.n1439 2588.24
R3223 VSS.n2646 VSS.n1439 2588.24
R3224 VSS.n2647 VSS.n2646 2588.24
R3225 VSS.n2648 VSS.n2647 2588.24
R3226 VSS.n2648 VSS.n1435 2588.24
R3227 VSS.n2654 VSS.n1435 2588.24
R3228 VSS.n2604 VSS.n2603 2588.24
R3229 VSS.n2605 VSS.n2604 2588.24
R3230 VSS.n2605 VSS.n1458 2588.24
R3231 VSS.n2611 VSS.n1458 2588.24
R3232 VSS.n2612 VSS.n2611 2588.24
R3233 VSS.n2613 VSS.n2612 2588.24
R3234 VSS.n2613 VSS.n1454 2588.24
R3235 VSS.n2620 VSS.n1454 2588.24
R3236 VSS.n2621 VSS.n2620 2588.24
R3237 VSS.n2622 VSS.n2621 2588.24
R3238 VSS.n2622 VSS.n1447 2588.24
R3239 VSS.n2075 VSS.n2042 2588.24
R3240 VSS.n2046 VSS.n2042 2588.24
R3241 VSS.n2068 VSS.n2046 2588.24
R3242 VSS.n2068 VSS.n2067 2588.24
R3243 VSS.n2067 VSS.n2066 2588.24
R3244 VSS.n2066 VSS.n2047 2588.24
R3245 VSS.n2060 VSS.n2047 2588.24
R3246 VSS.n2060 VSS.n2059 2588.24
R3247 VSS.n2059 VSS.n2058 2588.24
R3248 VSS.n2058 VSS.n2051 2588.24
R3249 VSS.n2052 VSS.n2051 2588.24
R3250 VSS.n2024 VSS.n1574 2588.24
R3251 VSS.n2025 VSS.n2024 2588.24
R3252 VSS.n2026 VSS.n2025 2588.24
R3253 VSS.n2026 VSS.n1570 2588.24
R3254 VSS.n2032 VSS.n1570 2588.24
R3255 VSS.n2033 VSS.n2032 2588.24
R3256 VSS.n2034 VSS.n2033 2588.24
R3257 VSS.n2034 VSS.n1566 2588.24
R3258 VSS.n2040 VSS.n1566 2588.24
R3259 VSS.n2041 VSS.n2040 2588.24
R3260 VSS.n2077 VSS.n2041 2588.24
R3261 VSS.n1991 VSS.n1589 2588.24
R3262 VSS.n1997 VSS.n1589 2588.24
R3263 VSS.n1998 VSS.n1997 2588.24
R3264 VSS.n1999 VSS.n1998 2588.24
R3265 VSS.n1999 VSS.n1585 2588.24
R3266 VSS.n2005 VSS.n1585 2588.24
R3267 VSS.n2006 VSS.n2005 2588.24
R3268 VSS.n2008 VSS.n2006 2588.24
R3269 VSS.n2008 VSS.n2007 2588.24
R3270 VSS.n2007 VSS.n1581 2588.24
R3271 VSS.n2015 VSS.n1581 2588.24
R3272 VSS.n1967 VSS.n1601 2588.24
R3273 VSS.n1973 VSS.n1601 2588.24
R3274 VSS.n1974 VSS.n1973 2588.24
R3275 VSS.n1975 VSS.n1974 2588.24
R3276 VSS.n1975 VSS.n1597 2588.24
R3277 VSS.n1981 VSS.n1597 2588.24
R3278 VSS.n1982 VSS.n1981 2588.24
R3279 VSS.n1983 VSS.n1982 2588.24
R3280 VSS.n1983 VSS.n1593 2588.24
R3281 VSS.n1989 VSS.n1593 2588.24
R3282 VSS.n1990 VSS.n1989 2588.24
R3283 VSS.n16005 VSS.n14011 2473.2
R3284 VSS.n12220 VSS.n12060 2473.2
R3285 VSS.n7171 VSS.n7170 2473.2
R3286 VSS.n5659 VSS.n5658 2473.2
R3287 VSS.n3042 VSS.n1272 2473.2
R3288 VSS.n15794 VSS.n15793 2099.35
R3289 VSS.n15782 VSS.n15680 2099.35
R3290 VSS.n15780 VSS.n15689 2099.35
R3291 VSS.n15771 VSS.n15770 2099.35
R3292 VSS.n15759 VSS.n15699 2099.35
R3293 VSS.n15757 VSS.n15708 2099.35
R3294 VSS.n15749 VSS.n15748 2099.35
R3295 VSS.n15737 VSS.n15718 2099.35
R3296 VSS.n15735 VSS.n15727 2099.35
R3297 VSS.n16019 VSS.n16018 2099.35
R3298 VSS.n16007 VSS.n14002 2099.35
R3299 VSS.n15886 VSS.n15885 2099.35
R3300 VSS.n15874 VSS.n15568 2099.35
R3301 VSS.n15872 VSS.n15577 2099.35
R3302 VSS.n15863 VSS.n15862 2099.35
R3303 VSS.n15851 VSS.n15587 2099.35
R3304 VSS.n15849 VSS.n15596 2099.35
R3305 VSS.n15841 VSS.n15840 2099.35
R3306 VSS.n15829 VSS.n15606 2099.35
R3307 VSS.n15827 VSS.n15615 2099.35
R3308 VSS.n15818 VSS.n15817 2099.35
R3309 VSS.n15806 VSS.n15625 2099.35
R3310 VSS.n15462 VSS.n15461 2099.35
R3311 VSS.n15472 VSS.n15471 2099.35
R3312 VSS.n15483 VSS.n14118 2099.35
R3313 VSS.n15485 VSS.n14111 2099.35
R3314 VSS.n15497 VSS.n15496 2099.35
R3315 VSS.n15507 VSS.n15506 2099.35
R3316 VSS.n15517 VSS.n14097 2099.35
R3317 VSS.n15519 VSS.n14090 2099.35
R3318 VSS.n15531 VSS.n15530 2099.35
R3319 VSS.n15541 VSS.n15540 2099.35
R3320 VSS.n15552 VSS.n14076 2099.35
R3321 VSS.n15227 VSS.n15226 2099.35
R3322 VSS.n15215 VSS.n15093 2099.35
R3323 VSS.n15213 VSS.n15102 2099.35
R3324 VSS.n15204 VSS.n15203 2099.35
R3325 VSS.n15192 VSS.n15112 2099.35
R3326 VSS.n15190 VSS.n15121 2099.35
R3327 VSS.n15182 VSS.n15181 2099.35
R3328 VSS.n15170 VSS.n15131 2099.35
R3329 VSS.n15168 VSS.n15140 2099.35
R3330 VSS.n15159 VSS.n15158 2099.35
R3331 VSS.n15445 VSS.n14143 2099.35
R3332 VSS.n15319 VSS.n15318 2099.35
R3333 VSS.n15307 VSS.n14981 2099.35
R3334 VSS.n15305 VSS.n14990 2099.35
R3335 VSS.n15296 VSS.n15295 2099.35
R3336 VSS.n15284 VSS.n15000 2099.35
R3337 VSS.n15282 VSS.n15009 2099.35
R3338 VSS.n15274 VSS.n15273 2099.35
R3339 VSS.n15262 VSS.n15019 2099.35
R3340 VSS.n15260 VSS.n15028 2099.35
R3341 VSS.n15251 VSS.n15250 2099.35
R3342 VSS.n15239 VSS.n15038 2099.35
R3343 VSS.n14885 VSS.n14295 2099.35
R3344 VSS.n14887 VSS.n14288 2099.35
R3345 VSS.n14899 VSS.n14898 2099.35
R3346 VSS.n14909 VSS.n14908 2099.35
R3347 VSS.n14920 VSS.n14274 2099.35
R3348 VSS.n14922 VSS.n14267 2099.35
R3349 VSS.n14933 VSS.n14932 2099.35
R3350 VSS.n14943 VSS.n14942 2099.35
R3351 VSS.n14954 VSS.n14253 2099.35
R3352 VSS.n14956 VSS.n14246 2099.35
R3353 VSS.n14968 VSS.n14967 2099.35
R3354 VSS.n14626 VSS.n14625 2099.35
R3355 VSS.n14614 VSS.n14484 2099.35
R3356 VSS.n14612 VSS.n14493 2099.35
R3357 VSS.n14603 VSS.n14602 2099.35
R3358 VSS.n14591 VSS.n14503 2099.35
R3359 VSS.n14589 VSS.n14512 2099.35
R3360 VSS.n14581 VSS.n14580 2099.35
R3361 VSS.n14569 VSS.n14522 2099.35
R3362 VSS.n14567 VSS.n14531 2099.35
R3363 VSS.n14558 VSS.n14557 2099.35
R3364 VSS.n14544 VSS.n14541 2099.35
R3365 VSS.n14718 VSS.n14717 2099.35
R3366 VSS.n14706 VSS.n14371 2099.35
R3367 VSS.n14704 VSS.n14381 2099.35
R3368 VSS.n14695 VSS.n14694 2099.35
R3369 VSS.n14683 VSS.n14391 2099.35
R3370 VSS.n14681 VSS.n14400 2099.35
R3371 VSS.n14673 VSS.n14672 2099.35
R3372 VSS.n14661 VSS.n14410 2099.35
R3373 VSS.n14659 VSS.n14419 2099.35
R3374 VSS.n14650 VSS.n14649 2099.35
R3375 VSS.n14638 VSS.n14429 2099.35
R3376 VSS.n12302 VSS.n12301 2099.35
R3377 VSS.n12290 VSS.n11994 2099.35
R3378 VSS.n12288 VSS.n12003 2099.35
R3379 VSS.n12279 VSS.n12278 2099.35
R3380 VSS.n12267 VSS.n12013 2099.35
R3381 VSS.n12265 VSS.n12022 2099.35
R3382 VSS.n12257 VSS.n12256 2099.35
R3383 VSS.n12245 VSS.n12032 2099.35
R3384 VSS.n12243 VSS.n12041 2099.35
R3385 VSS.n12234 VSS.n12233 2099.35
R3386 VSS.n12222 VSS.n12051 2099.35
R3387 VSS.n12394 VSS.n12393 2099.35
R3388 VSS.n12382 VSS.n11915 2099.35
R3389 VSS.n12380 VSS.n11924 2099.35
R3390 VSS.n12371 VSS.n12370 2099.35
R3391 VSS.n12359 VSS.n11934 2099.35
R3392 VSS.n12357 VSS.n11943 2099.35
R3393 VSS.n12349 VSS.n12348 2099.35
R3394 VSS.n12337 VSS.n11953 2099.35
R3395 VSS.n12335 VSS.n11962 2099.35
R3396 VSS.n12326 VSS.n12325 2099.35
R3397 VSS.n12314 VSS.n11972 2099.35
R3398 VSS.n11819 VSS.n11600 2099.35
R3399 VSS.n11821 VSS.n11593 2099.35
R3400 VSS.n11833 VSS.n11832 2099.35
R3401 VSS.n11843 VSS.n11842 2099.35
R3402 VSS.n11854 VSS.n11579 2099.35
R3403 VSS.n11856 VSS.n11572 2099.35
R3404 VSS.n11867 VSS.n11866 2099.35
R3405 VSS.n11877 VSS.n11876 2099.35
R3406 VSS.n11888 VSS.n11558 2099.35
R3407 VSS.n11890 VSS.n11551 2099.35
R3408 VSS.n11902 VSS.n11901 2099.35
R3409 VSS.n11675 VSS.n11665 2099.35
R3410 VSS.n11687 VSS.n11686 2099.35
R3411 VSS.n11697 VSS.n11696 2099.35
R3412 VSS.n11708 VSS.n11651 2099.35
R3413 VSS.n11710 VSS.n11644 2099.35
R3414 VSS.n11722 VSS.n11721 2099.35
R3415 VSS.n11731 VSS.n11730 2099.35
R3416 VSS.n11742 VSS.n11630 2099.35
R3417 VSS.n11744 VSS.n11623 2099.35
R3418 VSS.n11756 VSS.n11755 2099.35
R3419 VSS.n11766 VSS.n11765 2099.35
R3420 VSS.n13294 VSS.n13255 2099.35
R3421 VSS.n13292 VSS.n13256 2099.35
R3422 VSS.n13283 VSS.n13282 2099.35
R3423 VSS.n13269 VSS.n13266 2099.35
R3424 VSS.n13453 VSS.n13452 2099.35
R3425 VSS.n13441 VSS.n11436 2099.35
R3426 VSS.n13439 VSS.n11445 2099.35
R3427 VSS.n13431 VSS.n13430 2099.35
R3428 VSS.n13419 VSS.n11455 2099.35
R3429 VSS.n13417 VSS.n11464 2099.35
R3430 VSS.n13408 VSS.n13407 2099.35
R3431 VSS.n13154 VSS.n12574 2099.35
R3432 VSS.n13166 VSS.n13165 2099.35
R3433 VSS.n13176 VSS.n13175 2099.35
R3434 VSS.n13187 VSS.n12560 2099.35
R3435 VSS.n13189 VSS.n12553 2099.35
R3436 VSS.n13201 VSS.n13200 2099.35
R3437 VSS.n13210 VSS.n13209 2099.35
R3438 VSS.n13221 VSS.n12539 2099.35
R3439 VSS.n13223 VSS.n12532 2099.35
R3440 VSS.n13236 VSS.n13234 2099.35
R3441 VSS.n13247 VSS.n12524 2099.35
R3442 VSS.n13045 VSS.n12898 2099.35
R3443 VSS.n13043 VSS.n12899 2099.35
R3444 VSS.n13034 VSS.n13033 2099.35
R3445 VSS.n13022 VSS.n12909 2099.35
R3446 VSS.n13020 VSS.n12918 2099.35
R3447 VSS.n13011 VSS.n13010 2099.35
R3448 VSS.n13000 VSS.n12928 2099.35
R3449 VSS.n12998 VSS.n12937 2099.35
R3450 VSS.n12989 VSS.n12988 2099.35
R3451 VSS.n12977 VSS.n12947 2099.35
R3452 VSS.n12975 VSS.n12956 2099.35
R3453 VSS.n12797 VSS.n12715 2099.35
R3454 VSS.n12809 VSS.n12808 2099.35
R3455 VSS.n12819 VSS.n12818 2099.35
R3456 VSS.n12830 VSS.n12701 2099.35
R3457 VSS.n12832 VSS.n12694 2099.35
R3458 VSS.n12844 VSS.n12843 2099.35
R3459 VSS.n12853 VSS.n12852 2099.35
R3460 VSS.n12864 VSS.n12680 2099.35
R3461 VSS.n12866 VSS.n12673 2099.35
R3462 VSS.n12879 VSS.n12877 2099.35
R3463 VSS.n12890 VSS.n12665 2099.35
R3464 VSS.n7078 VSS.n7077 2099.35
R3465 VSS.n7088 VSS.n7087 2099.35
R3466 VSS.n7099 VSS.n7053 2099.35
R3467 VSS.n7101 VSS.n7046 2099.35
R3468 VSS.n7113 VSS.n7112 2099.35
R3469 VSS.n7123 VSS.n7122 2099.35
R3470 VSS.n7133 VSS.n7032 2099.35
R3471 VSS.n7135 VSS.n7025 2099.35
R3472 VSS.n7147 VSS.n7146 2099.35
R3473 VSS.n7157 VSS.n7156 2099.35
R3474 VSS.n7168 VSS.n7011 2099.35
R3475 VSS.n8759 VSS.n8758 2099.35
R3476 VSS.n8752 VSS.n8751 2099.35
R3477 VSS.n8925 VSS.n8924 2099.35
R3478 VSS.n8913 VSS.n6908 2099.35
R3479 VSS.n8911 VSS.n6917 2099.35
R3480 VSS.n8902 VSS.n8901 2099.35
R3481 VSS.n8891 VSS.n6927 2099.35
R3482 VSS.n8889 VSS.n6936 2099.35
R3483 VSS.n8880 VSS.n8879 2099.35
R3484 VSS.n8868 VSS.n6946 2099.35
R3485 VSS.n8866 VSS.n6955 2099.35
R3486 VSS.n8646 VSS.n7314 2099.35
R3487 VSS.n8648 VSS.n7307 2099.35
R3488 VSS.n8660 VSS.n8659 2099.35
R3489 VSS.n8670 VSS.n8669 2099.35
R3490 VSS.n8681 VSS.n7293 2099.35
R3491 VSS.n8683 VSS.n7286 2099.35
R3492 VSS.n8694 VSS.n8693 2099.35
R3493 VSS.n8704 VSS.n8703 2099.35
R3494 VSS.n8715 VSS.n7272 2099.35
R3495 VSS.n8717 VSS.n7265 2099.35
R3496 VSS.n8729 VSS.n8728 2099.35
R3497 VSS.n8537 VSS.n8536 2099.35
R3498 VSS.n8530 VSS.n8529 2099.35
R3499 VSS.n8518 VSS.n8390 2099.35
R3500 VSS.n8516 VSS.n8400 2099.35
R3501 VSS.n8507 VSS.n8506 2099.35
R3502 VSS.n8495 VSS.n8410 2099.35
R3503 VSS.n8493 VSS.n8419 2099.35
R3504 VSS.n8485 VSS.n8484 2099.35
R3505 VSS.n8473 VSS.n8429 2099.35
R3506 VSS.n8471 VSS.n8438 2099.35
R3507 VSS.n8462 VSS.n8461 2099.35
R3508 VSS.n8288 VSS.n7454 2099.35
R3509 VSS.n8290 VSS.n7447 2099.35
R3510 VSS.n8302 VSS.n8301 2099.35
R3511 VSS.n8312 VSS.n8311 2099.35
R3512 VSS.n8323 VSS.n7433 2099.35
R3513 VSS.n8325 VSS.n7426 2099.35
R3514 VSS.n8336 VSS.n8335 2099.35
R3515 VSS.n8346 VSS.n8345 2099.35
R3516 VSS.n8357 VSS.n7412 2099.35
R3517 VSS.n8359 VSS.n7405 2099.35
R3518 VSS.n8371 VSS.n8370 2099.35
R3519 VSS.n8179 VSS.n8178 2099.35
R3520 VSS.n8172 VSS.n8171 2099.35
R3521 VSS.n8160 VSS.n8032 2099.35
R3522 VSS.n8158 VSS.n8042 2099.35
R3523 VSS.n8149 VSS.n8148 2099.35
R3524 VSS.n8137 VSS.n8052 2099.35
R3525 VSS.n8135 VSS.n8061 2099.35
R3526 VSS.n8127 VSS.n8126 2099.35
R3527 VSS.n8115 VSS.n8071 2099.35
R3528 VSS.n8113 VSS.n8080 2099.35
R3529 VSS.n8104 VSS.n8103 2099.35
R3530 VSS.n7930 VSS.n7594 2099.35
R3531 VSS.n7932 VSS.n7587 2099.35
R3532 VSS.n7944 VSS.n7943 2099.35
R3533 VSS.n7954 VSS.n7953 2099.35
R3534 VSS.n7965 VSS.n7573 2099.35
R3535 VSS.n7967 VSS.n7566 2099.35
R3536 VSS.n7978 VSS.n7977 2099.35
R3537 VSS.n7988 VSS.n7987 2099.35
R3538 VSS.n7999 VSS.n7552 2099.35
R3539 VSS.n8001 VSS.n7545 2099.35
R3540 VSS.n8013 VSS.n8012 2099.35
R3541 VSS.n7832 VSS.n7831 2099.35
R3542 VSS.n7820 VSS.n7678 2099.35
R3543 VSS.n7818 VSS.n7688 2099.35
R3544 VSS.n7809 VSS.n7808 2099.35
R3545 VSS.n7797 VSS.n7698 2099.35
R3546 VSS.n7795 VSS.n7707 2099.35
R3547 VSS.n7787 VSS.n7786 2099.35
R3548 VSS.n7775 VSS.n7717 2099.35
R3549 VSS.n7773 VSS.n7726 2099.35
R3550 VSS.n7764 VSS.n7763 2099.35
R3551 VSS.n7752 VSS.n7736 2099.35
R3552 VSS.n5558 VSS.n5422 2099.35
R3553 VSS.n5556 VSS.n5423 2099.35
R3554 VSS.n5547 VSS.n5546 2099.35
R3555 VSS.n5535 VSS.n5433 2099.35
R3556 VSS.n5533 VSS.n5442 2099.35
R3557 VSS.n5524 VSS.n5523 2099.35
R3558 VSS.n5513 VSS.n5452 2099.35
R3559 VSS.n5511 VSS.n5461 2099.35
R3560 VSS.n5502 VSS.n5501 2099.35
R3561 VSS.n5490 VSS.n5471 2099.35
R3562 VSS.n5488 VSS.n5480 2099.35
R3563 VSS.n5321 VSS.n3745 2099.35
R3564 VSS.n5333 VSS.n5332 2099.35
R3565 VSS.n5343 VSS.n5342 2099.35
R3566 VSS.n5354 VSS.n3731 2099.35
R3567 VSS.n5356 VSS.n3724 2099.35
R3568 VSS.n5368 VSS.n5367 2099.35
R3569 VSS.n5377 VSS.n5376 2099.35
R3570 VSS.n5388 VSS.n3710 2099.35
R3571 VSS.n5390 VSS.n3703 2099.35
R3572 VSS.n5403 VSS.n5401 2099.35
R3573 VSS.n5414 VSS.n3695 2099.35
R3574 VSS.n5212 VSS.n5065 2099.35
R3575 VSS.n5210 VSS.n5066 2099.35
R3576 VSS.n5201 VSS.n5200 2099.35
R3577 VSS.n5189 VSS.n5076 2099.35
R3578 VSS.n5187 VSS.n5085 2099.35
R3579 VSS.n5178 VSS.n5177 2099.35
R3580 VSS.n5167 VSS.n5095 2099.35
R3581 VSS.n5165 VSS.n5104 2099.35
R3582 VSS.n5156 VSS.n5155 2099.35
R3583 VSS.n5144 VSS.n5114 2099.35
R3584 VSS.n5142 VSS.n5123 2099.35
R3585 VSS.n4964 VSS.n3886 2099.35
R3586 VSS.n4976 VSS.n4975 2099.35
R3587 VSS.n4986 VSS.n4985 2099.35
R3588 VSS.n4997 VSS.n3872 2099.35
R3589 VSS.n4999 VSS.n3865 2099.35
R3590 VSS.n5011 VSS.n5010 2099.35
R3591 VSS.n5020 VSS.n5019 2099.35
R3592 VSS.n5031 VSS.n3851 2099.35
R3593 VSS.n5033 VSS.n3844 2099.35
R3594 VSS.n5046 VSS.n5044 2099.35
R3595 VSS.n5057 VSS.n3836 2099.35
R3596 VSS.n4855 VSS.n4708 2099.35
R3597 VSS.n4853 VSS.n4709 2099.35
R3598 VSS.n4844 VSS.n4843 2099.35
R3599 VSS.n4832 VSS.n4719 2099.35
R3600 VSS.n4830 VSS.n4728 2099.35
R3601 VSS.n4821 VSS.n4820 2099.35
R3602 VSS.n4810 VSS.n4738 2099.35
R3603 VSS.n4808 VSS.n4747 2099.35
R3604 VSS.n4799 VSS.n4798 2099.35
R3605 VSS.n4787 VSS.n4757 2099.35
R3606 VSS.n4785 VSS.n4766 2099.35
R3607 VSS.n4607 VSS.n4027 2099.35
R3608 VSS.n4619 VSS.n4618 2099.35
R3609 VSS.n4629 VSS.n4628 2099.35
R3610 VSS.n4640 VSS.n4013 2099.35
R3611 VSS.n4642 VSS.n4006 2099.35
R3612 VSS.n4654 VSS.n4653 2099.35
R3613 VSS.n4663 VSS.n4662 2099.35
R3614 VSS.n4674 VSS.n3992 2099.35
R3615 VSS.n4676 VSS.n3985 2099.35
R3616 VSS.n4689 VSS.n4687 2099.35
R3617 VSS.n4700 VSS.n3977 2099.35
R3618 VSS.n4498 VSS.n4351 2099.35
R3619 VSS.n4496 VSS.n4352 2099.35
R3620 VSS.n4487 VSS.n4486 2099.35
R3621 VSS.n4475 VSS.n4362 2099.35
R3622 VSS.n4473 VSS.n4371 2099.35
R3623 VSS.n4464 VSS.n4463 2099.35
R3624 VSS.n4453 VSS.n4381 2099.35
R3625 VSS.n4451 VSS.n4390 2099.35
R3626 VSS.n4442 VSS.n4441 2099.35
R3627 VSS.n4430 VSS.n4400 2099.35
R3628 VSS.n4428 VSS.n4409 2099.35
R3629 VSS.n4250 VSS.n4168 2099.35
R3630 VSS.n4262 VSS.n4261 2099.35
R3631 VSS.n4272 VSS.n4271 2099.35
R3632 VSS.n4283 VSS.n4154 2099.35
R3633 VSS.n4285 VSS.n4147 2099.35
R3634 VSS.n4297 VSS.n4296 2099.35
R3635 VSS.n4306 VSS.n4305 2099.35
R3636 VSS.n4317 VSS.n4133 2099.35
R3637 VSS.n4319 VSS.n4126 2099.35
R3638 VSS.n4332 VSS.n4330 2099.35
R3639 VSS.n4343 VSS.n4118 2099.35
R3640 VSS.n2960 VSS.n2959 2099.35
R3641 VSS.n2948 VSS.n2809 2099.35
R3642 VSS.n2946 VSS.n2818 2099.35
R3643 VSS.n2937 VSS.n2936 2099.35
R3644 VSS.n2925 VSS.n2828 2099.35
R3645 VSS.n2923 VSS.n2837 2099.35
R3646 VSS.n2915 VSS.n2914 2099.35
R3647 VSS.n2903 VSS.n2847 2099.35
R3648 VSS.n2901 VSS.n2856 2099.35
R3649 VSS.n2892 VSS.n2891 2099.35
R3650 VSS.n2880 VSS.n2866 2099.35
R3651 VSS.n2703 VSS.n2702 2099.35
R3652 VSS.n2713 VSS.n2712 2099.35
R3653 VSS.n2724 VSS.n1359 2099.35
R3654 VSS.n2726 VSS.n1352 2099.35
R3655 VSS.n2738 VSS.n2737 2099.35
R3656 VSS.n2748 VSS.n2747 2099.35
R3657 VSS.n2758 VSS.n1338 2099.35
R3658 VSS.n2760 VSS.n1331 2099.35
R3659 VSS.n2772 VSS.n2771 2099.35
R3660 VSS.n2782 VSS.n2781 2099.35
R3661 VSS.n2793 VSS.n1317 2099.35
R3662 VSS.n2468 VSS.n2467 2099.35
R3663 VSS.n2456 VSS.n2334 2099.35
R3664 VSS.n2454 VSS.n2343 2099.35
R3665 VSS.n2445 VSS.n2444 2099.35
R3666 VSS.n2433 VSS.n2353 2099.35
R3667 VSS.n2431 VSS.n2362 2099.35
R3668 VSS.n2423 VSS.n2422 2099.35
R3669 VSS.n2411 VSS.n2372 2099.35
R3670 VSS.n2409 VSS.n2381 2099.35
R3671 VSS.n2400 VSS.n2399 2099.35
R3672 VSS.n2686 VSS.n1384 2099.35
R3673 VSS.n2560 VSS.n2559 2099.35
R3674 VSS.n2548 VSS.n2222 2099.35
R3675 VSS.n2546 VSS.n2231 2099.35
R3676 VSS.n2537 VSS.n2536 2099.35
R3677 VSS.n2525 VSS.n2241 2099.35
R3678 VSS.n2523 VSS.n2250 2099.35
R3679 VSS.n2515 VSS.n2514 2099.35
R3680 VSS.n2503 VSS.n2260 2099.35
R3681 VSS.n2501 VSS.n2269 2099.35
R3682 VSS.n2492 VSS.n2491 2099.35
R3683 VSS.n2480 VSS.n2279 2099.35
R3684 VSS.n2126 VSS.n1536 2099.35
R3685 VSS.n2128 VSS.n1529 2099.35
R3686 VSS.n2140 VSS.n2139 2099.35
R3687 VSS.n2150 VSS.n2149 2099.35
R3688 VSS.n2161 VSS.n1515 2099.35
R3689 VSS.n2163 VSS.n1508 2099.35
R3690 VSS.n2174 VSS.n2173 2099.35
R3691 VSS.n2184 VSS.n2183 2099.35
R3692 VSS.n2195 VSS.n1494 2099.35
R3693 VSS.n2197 VSS.n1487 2099.35
R3694 VSS.n2209 VSS.n2208 2099.35
R3695 VSS.n1867 VSS.n1866 2099.35
R3696 VSS.n1855 VSS.n1725 2099.35
R3697 VSS.n1853 VSS.n1734 2099.35
R3698 VSS.n1844 VSS.n1843 2099.35
R3699 VSS.n1832 VSS.n1744 2099.35
R3700 VSS.n1830 VSS.n1753 2099.35
R3701 VSS.n1822 VSS.n1821 2099.35
R3702 VSS.n1810 VSS.n1763 2099.35
R3703 VSS.n1808 VSS.n1772 2099.35
R3704 VSS.n1799 VSS.n1798 2099.35
R3705 VSS.n1785 VSS.n1782 2099.35
R3706 VSS.n1959 VSS.n1958 2099.35
R3707 VSS.n1947 VSS.n1612 2099.35
R3708 VSS.n1945 VSS.n1622 2099.35
R3709 VSS.n1936 VSS.n1935 2099.35
R3710 VSS.n1924 VSS.n1632 2099.35
R3711 VSS.n1922 VSS.n1641 2099.35
R3712 VSS.n1914 VSS.n1913 2099.35
R3713 VSS.n1902 VSS.n1651 2099.35
R3714 VSS.n1900 VSS.n1660 2099.35
R3715 VSS.n1891 VSS.n1890 2099.35
R3716 VSS.n1879 VSS.n1670 2099.35
R3717 VSS.n15667 VSS.n15666 1294.12
R3718 VSS.n15666 VSS.n15665 1294.12
R3719 VSS.n15665 VSS.n15639 1294.12
R3720 VSS.n15659 VSS.n15639 1294.12
R3721 VSS.n15659 VSS.n15658 1294.12
R3722 VSS.n15658 VSS.n15657 1294.12
R3723 VSS.n15657 VSS.n15643 1294.12
R3724 VSS.n15651 VSS.n15643 1294.12
R3725 VSS.n15651 VSS.n15650 1294.12
R3726 VSS.n15650 VSS.n15649 1294.12
R3727 VSS.n15649 VSS.n14043 1294.12
R3728 VSS.n15946 VSS.n14043 1294.12
R3729 VSS.n15895 VSS.n15894 1294.12
R3730 VSS.n15896 VSS.n15895 1294.12
R3731 VSS.n15896 VSS.n14065 1294.12
R3732 VSS.n15902 VSS.n14065 1294.12
R3733 VSS.n15903 VSS.n15902 1294.12
R3734 VSS.n15904 VSS.n15903 1294.12
R3735 VSS.n15904 VSS.n14061 1294.12
R3736 VSS.n15910 VSS.n14061 1294.12
R3737 VSS.n15911 VSS.n15910 1294.12
R3738 VSS.n15912 VSS.n15911 1294.12
R3739 VSS.n15912 VSS.n14057 1294.12
R3740 VSS.n15918 VSS.n14057 1294.12
R3741 VSS.n15439 VSS.n15438 1294.12
R3742 VSS.n15438 VSS.n15437 1294.12
R3743 VSS.n15437 VSS.n14146 1294.12
R3744 VSS.n15431 VSS.n14146 1294.12
R3745 VSS.n15431 VSS.n15430 1294.12
R3746 VSS.n15430 VSS.n15429 1294.12
R3747 VSS.n15429 VSS.n14151 1294.12
R3748 VSS.n15423 VSS.n14151 1294.12
R3749 VSS.n15423 VSS.n15422 1294.12
R3750 VSS.n15422 VSS.n15421 1294.12
R3751 VSS.n15421 VSS.n14155 1294.12
R3752 VSS.n15415 VSS.n14155 1294.12
R3753 VSS.n15080 VSS.n15079 1294.12
R3754 VSS.n15079 VSS.n15078 1294.12
R3755 VSS.n15078 VSS.n15052 1294.12
R3756 VSS.n15072 VSS.n15052 1294.12
R3757 VSS.n15072 VSS.n15071 1294.12
R3758 VSS.n15071 VSS.n15070 1294.12
R3759 VSS.n15070 VSS.n15056 1294.12
R3760 VSS.n15064 VSS.n15056 1294.12
R3761 VSS.n15064 VSS.n15063 1294.12
R3762 VSS.n15063 VSS.n15062 1294.12
R3763 VSS.n15062 VSS.n14207 1294.12
R3764 VSS.n15388 VSS.n14207 1294.12
R3765 VSS.n15332 VSS.n14234 1294.12
R3766 VSS.n15338 VSS.n14234 1294.12
R3767 VSS.n15339 VSS.n15338 1294.12
R3768 VSS.n15340 VSS.n15339 1294.12
R3769 VSS.n15340 VSS.n14230 1294.12
R3770 VSS.n15346 VSS.n14230 1294.12
R3771 VSS.n15347 VSS.n15346 1294.12
R3772 VSS.n15348 VSS.n15347 1294.12
R3773 VSS.n15348 VSS.n14226 1294.12
R3774 VSS.n15354 VSS.n14226 1294.12
R3775 VSS.n15355 VSS.n15354 1294.12
R3776 VSS.n15356 VSS.n15355 1294.12
R3777 VSS.n14861 VSS.n14301 1294.12
R3778 VSS.n14861 VSS.n14860 1294.12
R3779 VSS.n14860 VSS.n14859 1294.12
R3780 VSS.n14859 VSS.n14310 1294.12
R3781 VSS.n14853 VSS.n14310 1294.12
R3782 VSS.n14853 VSS.n14852 1294.12
R3783 VSS.n14852 VSS.n14851 1294.12
R3784 VSS.n14851 VSS.n14315 1294.12
R3785 VSS.n14845 VSS.n14315 1294.12
R3786 VSS.n14845 VSS.n14844 1294.12
R3787 VSS.n14844 VSS.n14843 1294.12
R3788 VSS.n14843 VSS.n14319 1294.12
R3789 VSS.n14471 VSS.n14470 1294.12
R3790 VSS.n14470 VSS.n14469 1294.12
R3791 VSS.n14469 VSS.n14443 1294.12
R3792 VSS.n14463 VSS.n14443 1294.12
R3793 VSS.n14463 VSS.n14462 1294.12
R3794 VSS.n14462 VSS.n14461 1294.12
R3795 VSS.n14461 VSS.n14447 1294.12
R3796 VSS.n14455 VSS.n14447 1294.12
R3797 VSS.n14455 VSS.n14454 1294.12
R3798 VSS.n14454 VSS.n14453 1294.12
R3799 VSS.n14453 VSS.n14339 1294.12
R3800 VSS.n14776 VSS.n14339 1294.12
R3801 VSS.n12102 VSS.n12100 1294.12
R3802 VSS.n12108 VSS.n12100 1294.12
R3803 VSS.n12109 VSS.n12108 1294.12
R3804 VSS.n12110 VSS.n12109 1294.12
R3805 VSS.n12110 VSS.n12096 1294.12
R3806 VSS.n12116 VSS.n12096 1294.12
R3807 VSS.n12117 VSS.n12116 1294.12
R3808 VSS.n12118 VSS.n12117 1294.12
R3809 VSS.n12118 VSS.n12092 1294.12
R3810 VSS.n12124 VSS.n12092 1294.12
R3811 VSS.n12125 VSS.n12124 1294.12
R3812 VSS.n12161 VSS.n12125 1294.12
R3813 VSS.n12407 VSS.n11539 1294.12
R3814 VSS.n12413 VSS.n11539 1294.12
R3815 VSS.n12414 VSS.n12413 1294.12
R3816 VSS.n12415 VSS.n12414 1294.12
R3817 VSS.n12415 VSS.n11535 1294.12
R3818 VSS.n12421 VSS.n11535 1294.12
R3819 VSS.n12422 VSS.n12421 1294.12
R3820 VSS.n12423 VSS.n12422 1294.12
R3821 VSS.n12423 VSS.n11531 1294.12
R3822 VSS.n12429 VSS.n11531 1294.12
R3823 VSS.n12430 VSS.n12429 1294.12
R3824 VSS.n12431 VSS.n12430 1294.12
R3825 VSS.n11806 VSS.n11607 1294.12
R3826 VSS.n11800 VSS.n11607 1294.12
R3827 VSS.n11800 VSS.n11799 1294.12
R3828 VSS.n11799 VSS.n11798 1294.12
R3829 VSS.n11798 VSS.n11778 1294.12
R3830 VSS.n11792 VSS.n11778 1294.12
R3831 VSS.n11792 VSS.n11791 1294.12
R3832 VSS.n11791 VSS.n11790 1294.12
R3833 VSS.n11790 VSS.n11782 1294.12
R3834 VSS.n11784 VSS.n11782 1294.12
R3835 VSS.n11784 VSS.n11511 1294.12
R3836 VSS.n12462 VSS.n11511 1294.12
R3837 VSS.n13395 VSS.n13394 1294.12
R3838 VSS.n13394 VSS.n13393 1294.12
R3839 VSS.n13393 VSS.n11486 1294.12
R3840 VSS.n13387 VSS.n11486 1294.12
R3841 VSS.n13387 VSS.n13386 1294.12
R3842 VSS.n13386 VSS.n13385 1294.12
R3843 VSS.n13385 VSS.n11490 1294.12
R3844 VSS.n13379 VSS.n11490 1294.12
R3845 VSS.n13379 VSS.n13378 1294.12
R3846 VSS.n13378 VSS.n13377 1294.12
R3847 VSS.n13377 VSS.n11494 1294.12
R3848 VSS.n13371 VSS.n11494 1294.12
R3849 VSS.n13318 VSS.n12515 1294.12
R3850 VSS.n13319 VSS.n13318 1294.12
R3851 VSS.n13320 VSS.n13319 1294.12
R3852 VSS.n13320 VSS.n12511 1294.12
R3853 VSS.n13326 VSS.n12511 1294.12
R3854 VSS.n13327 VSS.n13326 1294.12
R3855 VSS.n13328 VSS.n13327 1294.12
R3856 VSS.n13328 VSS.n12507 1294.12
R3857 VSS.n13335 VSS.n12507 1294.12
R3858 VSS.n13336 VSS.n13335 1294.12
R3859 VSS.n13337 VSS.n13336 1294.12
R3860 VSS.n13337 VSS.n12500 1294.12
R3861 VSS.n13146 VSS.n13145 1294.12
R3862 VSS.n13145 VSS.n13144 1294.12
R3863 VSS.n13144 VSS.n12587 1294.12
R3864 VSS.n13138 VSS.n12587 1294.12
R3865 VSS.n13138 VSS.n13137 1294.12
R3866 VSS.n13137 VSS.n13136 1294.12
R3867 VSS.n13136 VSS.n12591 1294.12
R3868 VSS.n13130 VSS.n12591 1294.12
R3869 VSS.n13130 VSS.n13129 1294.12
R3870 VSS.n13129 VSS.n13128 1294.12
R3871 VSS.n13128 VSS.n12595 1294.12
R3872 VSS.n13122 VSS.n12595 1294.12
R3873 VSS.n13069 VSS.n12656 1294.12
R3874 VSS.n13070 VSS.n13069 1294.12
R3875 VSS.n13071 VSS.n13070 1294.12
R3876 VSS.n13071 VSS.n12652 1294.12
R3877 VSS.n13077 VSS.n12652 1294.12
R3878 VSS.n13078 VSS.n13077 1294.12
R3879 VSS.n13079 VSS.n13078 1294.12
R3880 VSS.n13079 VSS.n12648 1294.12
R3881 VSS.n13086 VSS.n12648 1294.12
R3882 VSS.n13087 VSS.n13086 1294.12
R3883 VSS.n13088 VSS.n13087 1294.12
R3884 VSS.n13088 VSS.n12641 1294.12
R3885 VSS.n8855 VSS.n6966 1294.12
R3886 VSS.n8849 VSS.n6966 1294.12
R3887 VSS.n8849 VSS.n8848 1294.12
R3888 VSS.n8848 VSS.n8847 1294.12
R3889 VSS.n8847 VSS.n6971 1294.12
R3890 VSS.n8841 VSS.n6971 1294.12
R3891 VSS.n8841 VSS.n8840 1294.12
R3892 VSS.n8840 VSS.n8839 1294.12
R3893 VSS.n8839 VSS.n6975 1294.12
R3894 VSS.n8833 VSS.n6975 1294.12
R3895 VSS.n8833 VSS.n8832 1294.12
R3896 VSS.n8832 VSS.n8831 1294.12
R3897 VSS.n8774 VSS.n8773 1294.12
R3898 VSS.n8774 VSS.n7252 1294.12
R3899 VSS.n8780 VSS.n7252 1294.12
R3900 VSS.n8781 VSS.n8780 1294.12
R3901 VSS.n8782 VSS.n8781 1294.12
R3902 VSS.n8782 VSS.n7248 1294.12
R3903 VSS.n8788 VSS.n7248 1294.12
R3904 VSS.n8789 VSS.n8788 1294.12
R3905 VSS.n8791 VSS.n8789 1294.12
R3906 VSS.n8791 VSS.n8790 1294.12
R3907 VSS.n8790 VSS.n7244 1294.12
R3908 VSS.n8798 VSS.n7244 1294.12
R3909 VSS.n8633 VSS.n7321 1294.12
R3910 VSS.n8627 VSS.n7321 1294.12
R3911 VSS.n8627 VSS.n8626 1294.12
R3912 VSS.n8626 VSS.n8625 1294.12
R3913 VSS.n8625 VSS.n7327 1294.12
R3914 VSS.n8619 VSS.n7327 1294.12
R3915 VSS.n8619 VSS.n8618 1294.12
R3916 VSS.n8618 VSS.n8617 1294.12
R3917 VSS.n8617 VSS.n7331 1294.12
R3918 VSS.n8611 VSS.n7331 1294.12
R3919 VSS.n8611 VSS.n8610 1294.12
R3920 VSS.n8610 VSS.n8609 1294.12
R3921 VSS.n8552 VSS.n8551 1294.12
R3922 VSS.n8552 VSS.n7392 1294.12
R3923 VSS.n8558 VSS.n7392 1294.12
R3924 VSS.n8559 VSS.n8558 1294.12
R3925 VSS.n8560 VSS.n8559 1294.12
R3926 VSS.n8560 VSS.n7388 1294.12
R3927 VSS.n8566 VSS.n7388 1294.12
R3928 VSS.n8567 VSS.n8566 1294.12
R3929 VSS.n8569 VSS.n8567 1294.12
R3930 VSS.n8569 VSS.n8568 1294.12
R3931 VSS.n8568 VSS.n7384 1294.12
R3932 VSS.n8576 VSS.n7384 1294.12
R3933 VSS.n8275 VSS.n7461 1294.12
R3934 VSS.n8269 VSS.n7461 1294.12
R3935 VSS.n8269 VSS.n8268 1294.12
R3936 VSS.n8268 VSS.n8267 1294.12
R3937 VSS.n8267 VSS.n7467 1294.12
R3938 VSS.n8261 VSS.n7467 1294.12
R3939 VSS.n8261 VSS.n8260 1294.12
R3940 VSS.n8260 VSS.n8259 1294.12
R3941 VSS.n8259 VSS.n7471 1294.12
R3942 VSS.n8253 VSS.n7471 1294.12
R3943 VSS.n8253 VSS.n8252 1294.12
R3944 VSS.n8252 VSS.n8251 1294.12
R3945 VSS.n8194 VSS.n8193 1294.12
R3946 VSS.n8194 VSS.n7532 1294.12
R3947 VSS.n8200 VSS.n7532 1294.12
R3948 VSS.n8201 VSS.n8200 1294.12
R3949 VSS.n8202 VSS.n8201 1294.12
R3950 VSS.n8202 VSS.n7528 1294.12
R3951 VSS.n8208 VSS.n7528 1294.12
R3952 VSS.n8209 VSS.n8208 1294.12
R3953 VSS.n8211 VSS.n8209 1294.12
R3954 VSS.n8211 VSS.n8210 1294.12
R3955 VSS.n8210 VSS.n7524 1294.12
R3956 VSS.n8218 VSS.n7524 1294.12
R3957 VSS.n7917 VSS.n7601 1294.12
R3958 VSS.n7911 VSS.n7601 1294.12
R3959 VSS.n7911 VSS.n7910 1294.12
R3960 VSS.n7910 VSS.n7909 1294.12
R3961 VSS.n7909 VSS.n7607 1294.12
R3962 VSS.n7903 VSS.n7607 1294.12
R3963 VSS.n7903 VSS.n7902 1294.12
R3964 VSS.n7902 VSS.n7901 1294.12
R3965 VSS.n7901 VSS.n7611 1294.12
R3966 VSS.n7895 VSS.n7611 1294.12
R3967 VSS.n7895 VSS.n7894 1294.12
R3968 VSS.n7894 VSS.n7893 1294.12
R3969 VSS.n5582 VSS.n3686 1294.12
R3970 VSS.n5583 VSS.n5582 1294.12
R3971 VSS.n5584 VSS.n5583 1294.12
R3972 VSS.n5584 VSS.n3682 1294.12
R3973 VSS.n5590 VSS.n3682 1294.12
R3974 VSS.n5591 VSS.n5590 1294.12
R3975 VSS.n5592 VSS.n5591 1294.12
R3976 VSS.n5592 VSS.n3678 1294.12
R3977 VSS.n5599 VSS.n3678 1294.12
R3978 VSS.n5600 VSS.n5599 1294.12
R3979 VSS.n5601 VSS.n5600 1294.12
R3980 VSS.n5601 VSS.n3671 1294.12
R3981 VSS.n5313 VSS.n5312 1294.12
R3982 VSS.n5312 VSS.n5311 1294.12
R3983 VSS.n5311 VSS.n3758 1294.12
R3984 VSS.n5305 VSS.n3758 1294.12
R3985 VSS.n5305 VSS.n5304 1294.12
R3986 VSS.n5304 VSS.n5303 1294.12
R3987 VSS.n5303 VSS.n3762 1294.12
R3988 VSS.n5297 VSS.n3762 1294.12
R3989 VSS.n5297 VSS.n5296 1294.12
R3990 VSS.n5296 VSS.n5295 1294.12
R3991 VSS.n5295 VSS.n3766 1294.12
R3992 VSS.n5289 VSS.n3766 1294.12
R3993 VSS.n5236 VSS.n3827 1294.12
R3994 VSS.n5237 VSS.n5236 1294.12
R3995 VSS.n5238 VSS.n5237 1294.12
R3996 VSS.n5238 VSS.n3823 1294.12
R3997 VSS.n5244 VSS.n3823 1294.12
R3998 VSS.n5245 VSS.n5244 1294.12
R3999 VSS.n5246 VSS.n5245 1294.12
R4000 VSS.n5246 VSS.n3819 1294.12
R4001 VSS.n5253 VSS.n3819 1294.12
R4002 VSS.n5254 VSS.n5253 1294.12
R4003 VSS.n5255 VSS.n5254 1294.12
R4004 VSS.n5255 VSS.n3812 1294.12
R4005 VSS.n4956 VSS.n4955 1294.12
R4006 VSS.n4955 VSS.n4954 1294.12
R4007 VSS.n4954 VSS.n3899 1294.12
R4008 VSS.n4948 VSS.n3899 1294.12
R4009 VSS.n4948 VSS.n4947 1294.12
R4010 VSS.n4947 VSS.n4946 1294.12
R4011 VSS.n4946 VSS.n3903 1294.12
R4012 VSS.n4940 VSS.n3903 1294.12
R4013 VSS.n4940 VSS.n4939 1294.12
R4014 VSS.n4939 VSS.n4938 1294.12
R4015 VSS.n4938 VSS.n3907 1294.12
R4016 VSS.n4932 VSS.n3907 1294.12
R4017 VSS.n4879 VSS.n3968 1294.12
R4018 VSS.n4880 VSS.n4879 1294.12
R4019 VSS.n4881 VSS.n4880 1294.12
R4020 VSS.n4881 VSS.n3964 1294.12
R4021 VSS.n4887 VSS.n3964 1294.12
R4022 VSS.n4888 VSS.n4887 1294.12
R4023 VSS.n4889 VSS.n4888 1294.12
R4024 VSS.n4889 VSS.n3960 1294.12
R4025 VSS.n4896 VSS.n3960 1294.12
R4026 VSS.n4897 VSS.n4896 1294.12
R4027 VSS.n4898 VSS.n4897 1294.12
R4028 VSS.n4898 VSS.n3953 1294.12
R4029 VSS.n4599 VSS.n4598 1294.12
R4030 VSS.n4598 VSS.n4597 1294.12
R4031 VSS.n4597 VSS.n4040 1294.12
R4032 VSS.n4591 VSS.n4040 1294.12
R4033 VSS.n4591 VSS.n4590 1294.12
R4034 VSS.n4590 VSS.n4589 1294.12
R4035 VSS.n4589 VSS.n4044 1294.12
R4036 VSS.n4583 VSS.n4044 1294.12
R4037 VSS.n4583 VSS.n4582 1294.12
R4038 VSS.n4582 VSS.n4581 1294.12
R4039 VSS.n4581 VSS.n4048 1294.12
R4040 VSS.n4575 VSS.n4048 1294.12
R4041 VSS.n4522 VSS.n4109 1294.12
R4042 VSS.n4523 VSS.n4522 1294.12
R4043 VSS.n4524 VSS.n4523 1294.12
R4044 VSS.n4524 VSS.n4105 1294.12
R4045 VSS.n4530 VSS.n4105 1294.12
R4046 VSS.n4531 VSS.n4530 1294.12
R4047 VSS.n4532 VSS.n4531 1294.12
R4048 VSS.n4532 VSS.n4101 1294.12
R4049 VSS.n4539 VSS.n4101 1294.12
R4050 VSS.n4540 VSS.n4539 1294.12
R4051 VSS.n4541 VSS.n4540 1294.12
R4052 VSS.n4541 VSS.n4094 1294.12
R4053 VSS.n2969 VSS.n2968 1294.12
R4054 VSS.n2970 VSS.n2969 1294.12
R4055 VSS.n2970 VSS.n1306 1294.12
R4056 VSS.n2976 VSS.n1306 1294.12
R4057 VSS.n2977 VSS.n2976 1294.12
R4058 VSS.n2978 VSS.n2977 1294.12
R4059 VSS.n2978 VSS.n1302 1294.12
R4060 VSS.n2984 VSS.n1302 1294.12
R4061 VSS.n2985 VSS.n2984 1294.12
R4062 VSS.n2986 VSS.n2985 1294.12
R4063 VSS.n2986 VSS.n1298 1294.12
R4064 VSS.n2992 VSS.n1298 1294.12
R4065 VSS.n2680 VSS.n2679 1294.12
R4066 VSS.n2679 VSS.n2678 1294.12
R4067 VSS.n2678 VSS.n1387 1294.12
R4068 VSS.n2672 VSS.n1387 1294.12
R4069 VSS.n2672 VSS.n2671 1294.12
R4070 VSS.n2671 VSS.n2670 1294.12
R4071 VSS.n2670 VSS.n1392 1294.12
R4072 VSS.n2664 VSS.n1392 1294.12
R4073 VSS.n2664 VSS.n2663 1294.12
R4074 VSS.n2663 VSS.n2662 1294.12
R4075 VSS.n2662 VSS.n1396 1294.12
R4076 VSS.n2656 VSS.n1396 1294.12
R4077 VSS.n2321 VSS.n2320 1294.12
R4078 VSS.n2320 VSS.n2319 1294.12
R4079 VSS.n2319 VSS.n2293 1294.12
R4080 VSS.n2313 VSS.n2293 1294.12
R4081 VSS.n2313 VSS.n2312 1294.12
R4082 VSS.n2312 VSS.n2311 1294.12
R4083 VSS.n2311 VSS.n2297 1294.12
R4084 VSS.n2305 VSS.n2297 1294.12
R4085 VSS.n2305 VSS.n2304 1294.12
R4086 VSS.n2304 VSS.n2303 1294.12
R4087 VSS.n2303 VSS.n1448 1294.12
R4088 VSS.n2629 VSS.n1448 1294.12
R4089 VSS.n2573 VSS.n1475 1294.12
R4090 VSS.n2579 VSS.n1475 1294.12
R4091 VSS.n2580 VSS.n2579 1294.12
R4092 VSS.n2581 VSS.n2580 1294.12
R4093 VSS.n2581 VSS.n1471 1294.12
R4094 VSS.n2587 VSS.n1471 1294.12
R4095 VSS.n2588 VSS.n2587 1294.12
R4096 VSS.n2589 VSS.n2588 1294.12
R4097 VSS.n2589 VSS.n1467 1294.12
R4098 VSS.n2595 VSS.n1467 1294.12
R4099 VSS.n2596 VSS.n2595 1294.12
R4100 VSS.n2597 VSS.n2596 1294.12
R4101 VSS.n2102 VSS.n1542 1294.12
R4102 VSS.n2102 VSS.n2101 1294.12
R4103 VSS.n2101 VSS.n2100 1294.12
R4104 VSS.n2100 VSS.n1551 1294.12
R4105 VSS.n2094 VSS.n1551 1294.12
R4106 VSS.n2094 VSS.n2093 1294.12
R4107 VSS.n2093 VSS.n2092 1294.12
R4108 VSS.n2092 VSS.n1556 1294.12
R4109 VSS.n2086 VSS.n1556 1294.12
R4110 VSS.n2086 VSS.n2085 1294.12
R4111 VSS.n2085 VSS.n2084 1294.12
R4112 VSS.n2084 VSS.n1560 1294.12
R4113 VSS.n1712 VSS.n1711 1294.12
R4114 VSS.n1711 VSS.n1710 1294.12
R4115 VSS.n1710 VSS.n1684 1294.12
R4116 VSS.n1704 VSS.n1684 1294.12
R4117 VSS.n1704 VSS.n1703 1294.12
R4118 VSS.n1703 VSS.n1702 1294.12
R4119 VSS.n1702 VSS.n1688 1294.12
R4120 VSS.n1696 VSS.n1688 1294.12
R4121 VSS.n1696 VSS.n1695 1294.12
R4122 VSS.n1695 VSS.n1694 1294.12
R4123 VSS.n1694 VSS.n1580 1294.12
R4124 VSS.n2017 VSS.n1580 1294.12
R4125 VSS.n15946 VSS.n15945 1193.46
R4126 VSS.n15919 VSS.n15918 1193.46
R4127 VSS.n15415 VSS.n15414 1193.46
R4128 VSS.n15389 VSS.n15388 1193.46
R4129 VSS.n15356 VSS.n14221 1193.46
R4130 VSS.n14835 VSS.n14319 1193.46
R4131 VSS.n14776 VSS.n14775 1193.46
R4132 VSS.n12161 VSS.n12160 1193.46
R4133 VSS.n12431 VSS.n11526 1193.46
R4134 VSS.n12463 VSS.n12462 1193.46
R4135 VSS.n13371 VSS.n13370 1193.46
R4136 VSS.n13345 VSS.n12500 1193.46
R4137 VSS.n13122 VSS.n13121 1193.46
R4138 VSS.n13096 VSS.n12641 1193.46
R4139 VSS.n8831 VSS.n6979 1193.46
R4140 VSS.n8799 VSS.n8798 1193.46
R4141 VSS.n8609 VSS.n7335 1193.46
R4142 VSS.n8577 VSS.n8576 1193.46
R4143 VSS.n8251 VSS.n7475 1193.46
R4144 VSS.n8219 VSS.n8218 1193.46
R4145 VSS.n7893 VSS.n7615 1193.46
R4146 VSS.n5609 VSS.n3671 1193.46
R4147 VSS.n5289 VSS.n5288 1193.46
R4148 VSS.n5263 VSS.n3812 1193.46
R4149 VSS.n4932 VSS.n4931 1193.46
R4150 VSS.n4906 VSS.n3953 1193.46
R4151 VSS.n4575 VSS.n4574 1193.46
R4152 VSS.n4549 VSS.n4094 1193.46
R4153 VSS.n2993 VSS.n2992 1193.46
R4154 VSS.n2656 VSS.n2655 1193.46
R4155 VSS.n2630 VSS.n2629 1193.46
R4156 VSS.n2597 VSS.n1462 1193.46
R4157 VSS.n2076 VSS.n1560 1193.46
R4158 VSS.n2017 VSS.n2016 1193.46
R4159 VSS.n15995 VSS.n14011 1121.57
R4160 VSS.n12210 VSS.n12060 1121.57
R4161 VSS.n7170 VSS.n7003 1121.57
R4162 VSS.n6803 VSS.n6771 1121.57
R4163 VSS.n5658 VSS.n5657 1121.57
R4164 VSS.n3042 VSS.n3041 1121.57
R4165 VSS.n14726 VSS.n14725 1092.81
R4166 VSS.n12725 VSS.n12722 1092.81
R4167 VSS.n7839 VSS.n7669 1092.81
R4168 VSS.n6829 VSS.n6828 1092.81
R4169 VSS.n4178 VSS.n4175 1092.81
R4170 VSS.n1967 VSS.n1966 1092.81
R4171 VSS.n15945 VSS.n14037 690.196
R4172 VSS.n15920 VSS.n15919 690.196
R4173 VSS.n15414 VSS.n14193 690.196
R4174 VSS.n15390 VSS.n15389 690.196
R4175 VSS.n15362 VSS.n14221 690.196
R4176 VSS.n14835 VSS.n14834 690.196
R4177 VSS.n14775 VSS.n14333 690.196
R4178 VSS.n12160 VSS.n12086 690.196
R4179 VSS.n12135 VSS.n11526 690.196
R4180 VSS.n12463 VSS.n11510 690.196
R4181 VSS.n13370 VSS.n12487 690.196
R4182 VSS.n13346 VSS.n13345 690.196
R4183 VSS.n13121 VSS.n12628 690.196
R4184 VSS.n13097 VSS.n13096 690.196
R4185 VSS.n7224 VSS.n6979 690.196
R4186 VSS.n8799 VSS.n7237 690.196
R4187 VSS.n7364 VSS.n7335 690.196
R4188 VSS.n8577 VSS.n7377 690.196
R4189 VSS.n7504 VSS.n7475 690.196
R4190 VSS.n8219 VSS.n7517 690.196
R4191 VSS.n7644 VSS.n7615 690.196
R4192 VSS.n5610 VSS.n5609 690.196
R4193 VSS.n5288 VSS.n3799 690.196
R4194 VSS.n5264 VSS.n5263 690.196
R4195 VSS.n4931 VSS.n3940 690.196
R4196 VSS.n4907 VSS.n4906 690.196
R4197 VSS.n4574 VSS.n4081 690.196
R4198 VSS.n4550 VSS.n4549 690.196
R4199 VSS.n2994 VSS.n2993 690.196
R4200 VSS.n2655 VSS.n1434 690.196
R4201 VSS.n2631 VSS.n2630 690.196
R4202 VSS.n2603 VSS.n1462 690.196
R4203 VSS.n2076 VSS.n2075 690.196
R4204 VSS.n2016 VSS.n1574 690.196
R4205 VSS.n16009 VSS.n16008 585
R4206 VSS.n16008 VSS.n16007 585
R4207 VSS.n14004 VSS.n14000 585
R4208 VSS.n16018 VSS.n14000 585
R4209 VSS.n15729 VSS.n15728 585
R4210 VSS.n15728 VSS.n15727 585
R4211 VSS.n15739 VSS.n15738 585
R4212 VSS.n15738 VSS.n15737 585
R4213 VSS.n15720 VSS.n15716 585
R4214 VSS.n15748 VSS.n15716 585
R4215 VSS.n15712 VSS.n15709 585
R4216 VSS.n15709 VSS.n15708 585
R4217 VSS.n15761 VSS.n15760 585
R4218 VSS.n15760 VSS.n15759 585
R4219 VSS.n15701 VSS.n15697 585
R4220 VSS.n15770 VSS.n15697 585
R4221 VSS.n15693 VSS.n15690 585
R4222 VSS.n15690 VSS.n15689 585
R4223 VSS.n15784 VSS.n15783 585
R4224 VSS.n15783 VSS.n15782 585
R4225 VSS.n15682 VSS.n15675 585
R4226 VSS.n15793 VSS.n15675 585
R4227 VSS.n15677 VSS.n15676 585
R4228 VSS.n15678 VSS.n15677 585
R4229 VSS.n15808 VSS.n15807 585
R4230 VSS.n15807 VSS.n15806 585
R4231 VSS.n15627 VSS.n15623 585
R4232 VSS.n15817 VSS.n15623 585
R4233 VSS.n15619 VSS.n15616 585
R4234 VSS.n15616 VSS.n15615 585
R4235 VSS.n15831 VSS.n15830 585
R4236 VSS.n15830 VSS.n15829 585
R4237 VSS.n15608 VSS.n15604 585
R4238 VSS.n15840 VSS.n15604 585
R4239 VSS.n15600 VSS.n15597 585
R4240 VSS.n15597 VSS.n15596 585
R4241 VSS.n15853 VSS.n15852 585
R4242 VSS.n15852 VSS.n15851 585
R4243 VSS.n15589 VSS.n15585 585
R4244 VSS.n15862 VSS.n15585 585
R4245 VSS.n15581 VSS.n15578 585
R4246 VSS.n15578 VSS.n15577 585
R4247 VSS.n15876 VSS.n15875 585
R4248 VSS.n15875 VSS.n15874 585
R4249 VSS.n15570 VSS.n15564 585
R4250 VSS.n15885 VSS.n15564 585
R4251 VSS.n15565 VSS.n14071 585
R4252 VSS.n15566 VSS.n15565 585
R4253 VSS.n15551 VSS.n15550 585
R4254 VSS.n15552 VSS.n15551 585
R4255 VSS.n14081 VSS.n14080 585
R4256 VSS.n15541 VSS.n14081 585
R4257 VSS.n15533 VSS.n15532 585
R4258 VSS.n15532 VSS.n15531 585
R4259 VSS.n14092 VSS.n14091 585
R4260 VSS.n14091 VSS.n14090 585
R4261 VSS.n15516 VSS.n15515 585
R4262 VSS.n15517 VSS.n15516 585
R4263 VSS.n14102 VSS.n14101 585
R4264 VSS.n15507 VSS.n14102 585
R4265 VSS.n15499 VSS.n15498 585
R4266 VSS.n15498 VSS.n15497 585
R4267 VSS.n14113 VSS.n14112 585
R4268 VSS.n14112 VSS.n14111 585
R4269 VSS.n15482 VSS.n15481 585
R4270 VSS.n15483 VSS.n15482 585
R4271 VSS.n14123 VSS.n14122 585
R4272 VSS.n15472 VSS.n14123 585
R4273 VSS.n15464 VSS.n15463 585
R4274 VSS.n15463 VSS.n15462 585
R4275 VSS.n14134 VSS.n14133 585
R4276 VSS.n14133 VSS.n14132 585
R4277 VSS.n15447 VSS.n15446 585
R4278 VSS.n15446 VSS.n15445 585
R4279 VSS.n15150 VSS.n15148 585
R4280 VSS.n15158 VSS.n15148 585
R4281 VSS.n15144 VSS.n15141 585
R4282 VSS.n15141 VSS.n15140 585
R4283 VSS.n15172 VSS.n15171 585
R4284 VSS.n15171 VSS.n15170 585
R4285 VSS.n15133 VSS.n15129 585
R4286 VSS.n15181 VSS.n15129 585
R4287 VSS.n15125 VSS.n15122 585
R4288 VSS.n15122 VSS.n15121 585
R4289 VSS.n15194 VSS.n15193 585
R4290 VSS.n15193 VSS.n15192 585
R4291 VSS.n15114 VSS.n15110 585
R4292 VSS.n15203 VSS.n15110 585
R4293 VSS.n15106 VSS.n15103 585
R4294 VSS.n15103 VSS.n15102 585
R4295 VSS.n15217 VSS.n15216 585
R4296 VSS.n15216 VSS.n15215 585
R4297 VSS.n15095 VSS.n15088 585
R4298 VSS.n15226 VSS.n15088 585
R4299 VSS.n15090 VSS.n15089 585
R4300 VSS.n15091 VSS.n15090 585
R4301 VSS.n15241 VSS.n15240 585
R4302 VSS.n15240 VSS.n15239 585
R4303 VSS.n15040 VSS.n15036 585
R4304 VSS.n15250 VSS.n15036 585
R4305 VSS.n15032 VSS.n15029 585
R4306 VSS.n15029 VSS.n15028 585
R4307 VSS.n15264 VSS.n15263 585
R4308 VSS.n15263 VSS.n15262 585
R4309 VSS.n15021 VSS.n15017 585
R4310 VSS.n15273 VSS.n15017 585
R4311 VSS.n15013 VSS.n15010 585
R4312 VSS.n15010 VSS.n15009 585
R4313 VSS.n15286 VSS.n15285 585
R4314 VSS.n15285 VSS.n15284 585
R4315 VSS.n15002 VSS.n14998 585
R4316 VSS.n15295 VSS.n14998 585
R4317 VSS.n14994 VSS.n14991 585
R4318 VSS.n14991 VSS.n14990 585
R4319 VSS.n15309 VSS.n15308 585
R4320 VSS.n15308 VSS.n15307 585
R4321 VSS.n14983 VSS.n14979 585
R4322 VSS.n15318 VSS.n14979 585
R4323 VSS.n14977 VSS.n14976 585
R4324 VSS.n14977 VSS.n14238 585
R4325 VSS.n14970 VSS.n14969 585
R4326 VSS.n14969 VSS.n14968 585
R4327 VSS.n14248 VSS.n14247 585
R4328 VSS.n14247 VSS.n14246 585
R4329 VSS.n14953 VSS.n14952 585
R4330 VSS.n14954 VSS.n14953 585
R4331 VSS.n14258 VSS.n14257 585
R4332 VSS.n14943 VSS.n14258 585
R4333 VSS.n14935 VSS.n14934 585
R4334 VSS.n14934 VSS.n14933 585
R4335 VSS.n14269 VSS.n14268 585
R4336 VSS.n14268 VSS.n14267 585
R4337 VSS.n14919 VSS.n14918 585
R4338 VSS.n14920 VSS.n14919 585
R4339 VSS.n14279 VSS.n14278 585
R4340 VSS.n14909 VSS.n14279 585
R4341 VSS.n14901 VSS.n14900 585
R4342 VSS.n14900 VSS.n14899 585
R4343 VSS.n14290 VSS.n14289 585
R4344 VSS.n14289 VSS.n14288 585
R4345 VSS.n14884 VSS.n14883 585
R4346 VSS.n14885 VSS.n14884 585
R4347 VSS.n14300 VSS.n14299 585
R4348 VSS.n14874 VSS.n14300 585
R4349 VSS.n14546 VSS.n14545 585
R4350 VSS.n14545 VSS.n14544 585
R4351 VSS.n14543 VSS.n14539 585
R4352 VSS.n14557 VSS.n14539 585
R4353 VSS.n14535 VSS.n14532 585
R4354 VSS.n14532 VSS.n14531 585
R4355 VSS.n14571 VSS.n14570 585
R4356 VSS.n14570 VSS.n14569 585
R4357 VSS.n14524 VSS.n14520 585
R4358 VSS.n14580 VSS.n14520 585
R4359 VSS.n14516 VSS.n14513 585
R4360 VSS.n14513 VSS.n14512 585
R4361 VSS.n14593 VSS.n14592 585
R4362 VSS.n14592 VSS.n14591 585
R4363 VSS.n14505 VSS.n14501 585
R4364 VSS.n14602 VSS.n14501 585
R4365 VSS.n14497 VSS.n14494 585
R4366 VSS.n14494 VSS.n14493 585
R4367 VSS.n14616 VSS.n14615 585
R4368 VSS.n14615 VSS.n14614 585
R4369 VSS.n14486 VSS.n14479 585
R4370 VSS.n14625 VSS.n14479 585
R4371 VSS.n14481 VSS.n14480 585
R4372 VSS.n14482 VSS.n14481 585
R4373 VSS.n14640 VSS.n14639 585
R4374 VSS.n14639 VSS.n14638 585
R4375 VSS.n14431 VSS.n14427 585
R4376 VSS.n14649 VSS.n14427 585
R4377 VSS.n14423 VSS.n14420 585
R4378 VSS.n14420 VSS.n14419 585
R4379 VSS.n14663 VSS.n14662 585
R4380 VSS.n14662 VSS.n14661 585
R4381 VSS.n14412 VSS.n14408 585
R4382 VSS.n14672 VSS.n14408 585
R4383 VSS.n14404 VSS.n14401 585
R4384 VSS.n14401 VSS.n14400 585
R4385 VSS.n14685 VSS.n14684 585
R4386 VSS.n14684 VSS.n14683 585
R4387 VSS.n14393 VSS.n14389 585
R4388 VSS.n14694 VSS.n14389 585
R4389 VSS.n14385 VSS.n14382 585
R4390 VSS.n14382 VSS.n14381 585
R4391 VSS.n14708 VSS.n14707 585
R4392 VSS.n14707 VSS.n14706 585
R4393 VSS.n14373 VSS.n14370 585
R4394 VSS.n14717 VSS.n14370 585
R4395 VSS.n14723 VSS.n14722 585
R4396 VSS.n14724 VSS.n14723 585
R4397 VSS.n12224 VSS.n12223 585
R4398 VSS.n12223 VSS.n12222 585
R4399 VSS.n12053 VSS.n12049 585
R4400 VSS.n12233 VSS.n12049 585
R4401 VSS.n12045 VSS.n12042 585
R4402 VSS.n12042 VSS.n12041 585
R4403 VSS.n12247 VSS.n12246 585
R4404 VSS.n12246 VSS.n12245 585
R4405 VSS.n12034 VSS.n12030 585
R4406 VSS.n12256 VSS.n12030 585
R4407 VSS.n12026 VSS.n12023 585
R4408 VSS.n12023 VSS.n12022 585
R4409 VSS.n12269 VSS.n12268 585
R4410 VSS.n12268 VSS.n12267 585
R4411 VSS.n12015 VSS.n12011 585
R4412 VSS.n12278 VSS.n12011 585
R4413 VSS.n12007 VSS.n12004 585
R4414 VSS.n12004 VSS.n12003 585
R4415 VSS.n12292 VSS.n12291 585
R4416 VSS.n12291 VSS.n12290 585
R4417 VSS.n11996 VSS.n11989 585
R4418 VSS.n12301 VSS.n11989 585
R4419 VSS.n11991 VSS.n11990 585
R4420 VSS.n11992 VSS.n11991 585
R4421 VSS.n12316 VSS.n12315 585
R4422 VSS.n12315 VSS.n12314 585
R4423 VSS.n11974 VSS.n11970 585
R4424 VSS.n12325 VSS.n11970 585
R4425 VSS.n11966 VSS.n11963 585
R4426 VSS.n11963 VSS.n11962 585
R4427 VSS.n12339 VSS.n12338 585
R4428 VSS.n12338 VSS.n12337 585
R4429 VSS.n11955 VSS.n11951 585
R4430 VSS.n12348 VSS.n11951 585
R4431 VSS.n11947 VSS.n11944 585
R4432 VSS.n11944 VSS.n11943 585
R4433 VSS.n12361 VSS.n12360 585
R4434 VSS.n12360 VSS.n12359 585
R4435 VSS.n11936 VSS.n11932 585
R4436 VSS.n12370 VSS.n11932 585
R4437 VSS.n11928 VSS.n11925 585
R4438 VSS.n11925 VSS.n11924 585
R4439 VSS.n12384 VSS.n12383 585
R4440 VSS.n12383 VSS.n12382 585
R4441 VSS.n11917 VSS.n11913 585
R4442 VSS.n12393 VSS.n11913 585
R4443 VSS.n11911 VSS.n11910 585
R4444 VSS.n11911 VSS.n11543 585
R4445 VSS.n11904 VSS.n11903 585
R4446 VSS.n11903 VSS.n11902 585
R4447 VSS.n11553 VSS.n11552 585
R4448 VSS.n11552 VSS.n11551 585
R4449 VSS.n11887 VSS.n11886 585
R4450 VSS.n11888 VSS.n11887 585
R4451 VSS.n11563 VSS.n11562 585
R4452 VSS.n11877 VSS.n11563 585
R4453 VSS.n11869 VSS.n11868 585
R4454 VSS.n11868 VSS.n11867 585
R4455 VSS.n11574 VSS.n11573 585
R4456 VSS.n11573 VSS.n11572 585
R4457 VSS.n11853 VSS.n11852 585
R4458 VSS.n11854 VSS.n11853 585
R4459 VSS.n11584 VSS.n11583 585
R4460 VSS.n11843 VSS.n11584 585
R4461 VSS.n11835 VSS.n11834 585
R4462 VSS.n11834 VSS.n11833 585
R4463 VSS.n11595 VSS.n11594 585
R4464 VSS.n11594 VSS.n11593 585
R4465 VSS.n11818 VSS.n11817 585
R4466 VSS.n11819 VSS.n11818 585
R4467 VSS.n11605 VSS.n11604 585
R4468 VSS.n11808 VSS.n11605 585
R4469 VSS.n11617 VSS.n11613 585
R4470 VSS.n11766 VSS.n11613 585
R4471 VSS.n11758 VSS.n11757 585
R4472 VSS.n11757 VSS.n11756 585
R4473 VSS.n11625 VSS.n11624 585
R4474 VSS.n11624 VSS.n11623 585
R4475 VSS.n11741 VSS.n11740 585
R4476 VSS.n11742 VSS.n11741 585
R4477 VSS.n11635 VSS.n11634 585
R4478 VSS.n11731 VSS.n11635 585
R4479 VSS.n11724 VSS.n11723 585
R4480 VSS.n11723 VSS.n11722 585
R4481 VSS.n11646 VSS.n11645 585
R4482 VSS.n11645 VSS.n11644 585
R4483 VSS.n11707 VSS.n11706 585
R4484 VSS.n11708 VSS.n11707 585
R4485 VSS.n11656 VSS.n11655 585
R4486 VSS.n11697 VSS.n11656 585
R4487 VSS.n11689 VSS.n11688 585
R4488 VSS.n11688 VSS.n11687 585
R4489 VSS.n11667 VSS.n11666 585
R4490 VSS.n11666 VSS.n11665 585
R4491 VSS.n11672 VSS.n11481 585
R4492 VSS.n11673 VSS.n11672 585
R4493 VSS.n11476 VSS.n11472 585
R4494 VSS.n13407 VSS.n11472 585
R4495 VSS.n11468 VSS.n11465 585
R4496 VSS.n11465 VSS.n11464 585
R4497 VSS.n13421 VSS.n13420 585
R4498 VSS.n13420 VSS.n13419 585
R4499 VSS.n11457 VSS.n11453 585
R4500 VSS.n13430 VSS.n11453 585
R4501 VSS.n11449 VSS.n11446 585
R4502 VSS.n11446 VSS.n11445 585
R4503 VSS.n13443 VSS.n13442 585
R4504 VSS.n13442 VSS.n13441 585
R4505 VSS.n11438 VSS.n11434 585
R4506 VSS.n13452 VSS.n11434 585
R4507 VSS.n13271 VSS.n13270 585
R4508 VSS.n13270 VSS.n13269 585
R4509 VSS.n13268 VSS.n13264 585
R4510 VSS.n13282 VSS.n13264 585
R4511 VSS.n13260 VSS.n13257 585
R4512 VSS.n13257 VSS.n13256 585
R4513 VSS.n13296 VSS.n13295 585
R4514 VSS.n13295 VSS.n13294 585
R4515 VSS.n13304 VSS.n12517 585
R4516 VSS.n13305 VSS.n13304 585
R4517 VSS.n13246 VSS.n13245 585
R4518 VSS.n13247 VSS.n13246 585
R4519 VSS.n13238 VSS.n13237 585
R4520 VSS.n13237 VSS.n13236 585
R4521 VSS.n12534 VSS.n12533 585
R4522 VSS.n12533 VSS.n12532 585
R4523 VSS.n13220 VSS.n13219 585
R4524 VSS.n13221 VSS.n13220 585
R4525 VSS.n12544 VSS.n12543 585
R4526 VSS.n13210 VSS.n12544 585
R4527 VSS.n13203 VSS.n13202 585
R4528 VSS.n13202 VSS.n13201 585
R4529 VSS.n12555 VSS.n12554 585
R4530 VSS.n12554 VSS.n12553 585
R4531 VSS.n13186 VSS.n13185 585
R4532 VSS.n13187 VSS.n13186 585
R4533 VSS.n12565 VSS.n12564 585
R4534 VSS.n13176 VSS.n12565 585
R4535 VSS.n13168 VSS.n13167 585
R4536 VSS.n13167 VSS.n13166 585
R4537 VSS.n12576 VSS.n12575 585
R4538 VSS.n12575 VSS.n12574 585
R4539 VSS.n13151 VSS.n13150 585
R4540 VSS.n13152 VSS.n13151 585
R4541 VSS.n12961 VSS.n12957 585
R4542 VSS.n12957 VSS.n12956 585
R4543 VSS.n12979 VSS.n12978 585
R4544 VSS.n12978 VSS.n12977 585
R4545 VSS.n12949 VSS.n12945 585
R4546 VSS.n12988 VSS.n12945 585
R4547 VSS.n12941 VSS.n12938 585
R4548 VSS.n12938 VSS.n12937 585
R4549 VSS.n13002 VSS.n13001 585
R4550 VSS.n13001 VSS.n13000 585
R4551 VSS.n12930 VSS.n12926 585
R4552 VSS.n13010 VSS.n12926 585
R4553 VSS.n12922 VSS.n12919 585
R4554 VSS.n12919 VSS.n12918 585
R4555 VSS.n13024 VSS.n13023 585
R4556 VSS.n13023 VSS.n13022 585
R4557 VSS.n12911 VSS.n12907 585
R4558 VSS.n13033 VSS.n12907 585
R4559 VSS.n12903 VSS.n12900 585
R4560 VSS.n12900 VSS.n12899 585
R4561 VSS.n13047 VSS.n13046 585
R4562 VSS.n13046 VSS.n13045 585
R4563 VSS.n13055 VSS.n12658 585
R4564 VSS.n13056 VSS.n13055 585
R4565 VSS.n12889 VSS.n12888 585
R4566 VSS.n12890 VSS.n12889 585
R4567 VSS.n12881 VSS.n12880 585
R4568 VSS.n12880 VSS.n12879 585
R4569 VSS.n12675 VSS.n12674 585
R4570 VSS.n12674 VSS.n12673 585
R4571 VSS.n12863 VSS.n12862 585
R4572 VSS.n12864 VSS.n12863 585
R4573 VSS.n12685 VSS.n12684 585
R4574 VSS.n12853 VSS.n12685 585
R4575 VSS.n12846 VSS.n12845 585
R4576 VSS.n12845 VSS.n12844 585
R4577 VSS.n12696 VSS.n12695 585
R4578 VSS.n12695 VSS.n12694 585
R4579 VSS.n12829 VSS.n12828 585
R4580 VSS.n12830 VSS.n12829 585
R4581 VSS.n12706 VSS.n12705 585
R4582 VSS.n12819 VSS.n12706 585
R4583 VSS.n12811 VSS.n12810 585
R4584 VSS.n12810 VSS.n12809 585
R4585 VSS.n12717 VSS.n12716 585
R4586 VSS.n12716 VSS.n12715 585
R4587 VSS.n12794 VSS.n12793 585
R4588 VSS.n12795 VSS.n12794 585
R4589 VSS.n7167 VSS.n7166 585
R4590 VSS.n7168 VSS.n7167 585
R4591 VSS.n7016 VSS.n7015 585
R4592 VSS.n7157 VSS.n7016 585
R4593 VSS.n7149 VSS.n7148 585
R4594 VSS.n7148 VSS.n7147 585
R4595 VSS.n7027 VSS.n7026 585
R4596 VSS.n7026 VSS.n7025 585
R4597 VSS.n7132 VSS.n7131 585
R4598 VSS.n7133 VSS.n7132 585
R4599 VSS.n7037 VSS.n7036 585
R4600 VSS.n7123 VSS.n7037 585
R4601 VSS.n7115 VSS.n7114 585
R4602 VSS.n7114 VSS.n7113 585
R4603 VSS.n7048 VSS.n7047 585
R4604 VSS.n7047 VSS.n7046 585
R4605 VSS.n7098 VSS.n7097 585
R4606 VSS.n7099 VSS.n7098 585
R4607 VSS.n7058 VSS.n7057 585
R4608 VSS.n7088 VSS.n7058 585
R4609 VSS.n7080 VSS.n7079 585
R4610 VSS.n7079 VSS.n7078 585
R4611 VSS.n7068 VSS.n7067 585
R4612 VSS.n7067 VSS.n6965 585
R4613 VSS.n6959 VSS.n6956 585
R4614 VSS.n6956 VSS.n6955 585
R4615 VSS.n8870 VSS.n8869 585
R4616 VSS.n8869 VSS.n8868 585
R4617 VSS.n6948 VSS.n6944 585
R4618 VSS.n8879 VSS.n6944 585
R4619 VSS.n6940 VSS.n6937 585
R4620 VSS.n6937 VSS.n6936 585
R4621 VSS.n8893 VSS.n8892 585
R4622 VSS.n8892 VSS.n8891 585
R4623 VSS.n6929 VSS.n6925 585
R4624 VSS.n8901 VSS.n6925 585
R4625 VSS.n6921 VSS.n6918 585
R4626 VSS.n6918 VSS.n6917 585
R4627 VSS.n8915 VSS.n8914 585
R4628 VSS.n8914 VSS.n8913 585
R4629 VSS.n6910 VSS.n6906 585
R4630 VSS.n8924 VSS.n6906 585
R4631 VSS.n8750 VSS.n8749 585
R4632 VSS.n8751 VSS.n8750 585
R4633 VSS.n8757 VSS.n8756 585
R4634 VSS.n8758 VSS.n8757 585
R4635 VSS.n8763 VSS.n8762 585
R4636 VSS.n8762 VSS.n7256 585
R4637 VSS.n8731 VSS.n8730 585
R4638 VSS.n8730 VSS.n8729 585
R4639 VSS.n7267 VSS.n7266 585
R4640 VSS.n7266 VSS.n7265 585
R4641 VSS.n8714 VSS.n8713 585
R4642 VSS.n8715 VSS.n8714 585
R4643 VSS.n7277 VSS.n7276 585
R4644 VSS.n8704 VSS.n7277 585
R4645 VSS.n8696 VSS.n8695 585
R4646 VSS.n8695 VSS.n8694 585
R4647 VSS.n7288 VSS.n7287 585
R4648 VSS.n7287 VSS.n7286 585
R4649 VSS.n8680 VSS.n8679 585
R4650 VSS.n8681 VSS.n8680 585
R4651 VSS.n7298 VSS.n7297 585
R4652 VSS.n8670 VSS.n7298 585
R4653 VSS.n8662 VSS.n8661 585
R4654 VSS.n8661 VSS.n8660 585
R4655 VSS.n7309 VSS.n7308 585
R4656 VSS.n7308 VSS.n7307 585
R4657 VSS.n8645 VSS.n8644 585
R4658 VSS.n8646 VSS.n8645 585
R4659 VSS.n7319 VSS.n7318 585
R4660 VSS.n8635 VSS.n7319 585
R4661 VSS.n8449 VSS.n8446 585
R4662 VSS.n8461 VSS.n8446 585
R4663 VSS.n8442 VSS.n8439 585
R4664 VSS.n8439 VSS.n8438 585
R4665 VSS.n8475 VSS.n8474 585
R4666 VSS.n8474 VSS.n8473 585
R4667 VSS.n8431 VSS.n8427 585
R4668 VSS.n8484 VSS.n8427 585
R4669 VSS.n8423 VSS.n8420 585
R4670 VSS.n8420 VSS.n8419 585
R4671 VSS.n8497 VSS.n8496 585
R4672 VSS.n8496 VSS.n8495 585
R4673 VSS.n8412 VSS.n8408 585
R4674 VSS.n8506 VSS.n8408 585
R4675 VSS.n8404 VSS.n8401 585
R4676 VSS.n8401 VSS.n8400 585
R4677 VSS.n8520 VSS.n8519 585
R4678 VSS.n8519 VSS.n8518 585
R4679 VSS.n8392 VSS.n8389 585
R4680 VSS.n8529 VSS.n8389 585
R4681 VSS.n8535 VSS.n8534 585
R4682 VSS.n8536 VSS.n8535 585
R4683 VSS.n8541 VSS.n8540 585
R4684 VSS.n8540 VSS.n7396 585
R4685 VSS.n8373 VSS.n8372 585
R4686 VSS.n8372 VSS.n8371 585
R4687 VSS.n7407 VSS.n7406 585
R4688 VSS.n7406 VSS.n7405 585
R4689 VSS.n8356 VSS.n8355 585
R4690 VSS.n8357 VSS.n8356 585
R4691 VSS.n7417 VSS.n7416 585
R4692 VSS.n8346 VSS.n7417 585
R4693 VSS.n8338 VSS.n8337 585
R4694 VSS.n8337 VSS.n8336 585
R4695 VSS.n7428 VSS.n7427 585
R4696 VSS.n7427 VSS.n7426 585
R4697 VSS.n8322 VSS.n8321 585
R4698 VSS.n8323 VSS.n8322 585
R4699 VSS.n7438 VSS.n7437 585
R4700 VSS.n8312 VSS.n7438 585
R4701 VSS.n8304 VSS.n8303 585
R4702 VSS.n8303 VSS.n8302 585
R4703 VSS.n7449 VSS.n7448 585
R4704 VSS.n7448 VSS.n7447 585
R4705 VSS.n8287 VSS.n8286 585
R4706 VSS.n8288 VSS.n8287 585
R4707 VSS.n7459 VSS.n7458 585
R4708 VSS.n8277 VSS.n7459 585
R4709 VSS.n8091 VSS.n8088 585
R4710 VSS.n8103 VSS.n8088 585
R4711 VSS.n8084 VSS.n8081 585
R4712 VSS.n8081 VSS.n8080 585
R4713 VSS.n8117 VSS.n8116 585
R4714 VSS.n8116 VSS.n8115 585
R4715 VSS.n8073 VSS.n8069 585
R4716 VSS.n8126 VSS.n8069 585
R4717 VSS.n8065 VSS.n8062 585
R4718 VSS.n8062 VSS.n8061 585
R4719 VSS.n8139 VSS.n8138 585
R4720 VSS.n8138 VSS.n8137 585
R4721 VSS.n8054 VSS.n8050 585
R4722 VSS.n8148 VSS.n8050 585
R4723 VSS.n8046 VSS.n8043 585
R4724 VSS.n8043 VSS.n8042 585
R4725 VSS.n8162 VSS.n8161 585
R4726 VSS.n8161 VSS.n8160 585
R4727 VSS.n8034 VSS.n8031 585
R4728 VSS.n8171 VSS.n8031 585
R4729 VSS.n8177 VSS.n8176 585
R4730 VSS.n8178 VSS.n8177 585
R4731 VSS.n8183 VSS.n8182 585
R4732 VSS.n8182 VSS.n7536 585
R4733 VSS.n8015 VSS.n8014 585
R4734 VSS.n8014 VSS.n8013 585
R4735 VSS.n7547 VSS.n7546 585
R4736 VSS.n7546 VSS.n7545 585
R4737 VSS.n7998 VSS.n7997 585
R4738 VSS.n7999 VSS.n7998 585
R4739 VSS.n7557 VSS.n7556 585
R4740 VSS.n7988 VSS.n7557 585
R4741 VSS.n7980 VSS.n7979 585
R4742 VSS.n7979 VSS.n7978 585
R4743 VSS.n7568 VSS.n7567 585
R4744 VSS.n7567 VSS.n7566 585
R4745 VSS.n7964 VSS.n7963 585
R4746 VSS.n7965 VSS.n7964 585
R4747 VSS.n7578 VSS.n7577 585
R4748 VSS.n7954 VSS.n7578 585
R4749 VSS.n7946 VSS.n7945 585
R4750 VSS.n7945 VSS.n7944 585
R4751 VSS.n7589 VSS.n7588 585
R4752 VSS.n7588 VSS.n7587 585
R4753 VSS.n7929 VSS.n7928 585
R4754 VSS.n7930 VSS.n7929 585
R4755 VSS.n7599 VSS.n7598 585
R4756 VSS.n7919 VSS.n7599 585
R4757 VSS.n7754 VSS.n7753 585
R4758 VSS.n7753 VSS.n7752 585
R4759 VSS.n7738 VSS.n7734 585
R4760 VSS.n7763 VSS.n7734 585
R4761 VSS.n7730 VSS.n7727 585
R4762 VSS.n7727 VSS.n7726 585
R4763 VSS.n7777 VSS.n7776 585
R4764 VSS.n7776 VSS.n7775 585
R4765 VSS.n7719 VSS.n7715 585
R4766 VSS.n7786 VSS.n7715 585
R4767 VSS.n7711 VSS.n7708 585
R4768 VSS.n7708 VSS.n7707 585
R4769 VSS.n7799 VSS.n7798 585
R4770 VSS.n7798 VSS.n7797 585
R4771 VSS.n7700 VSS.n7696 585
R4772 VSS.n7808 VSS.n7696 585
R4773 VSS.n7692 VSS.n7689 585
R4774 VSS.n7689 VSS.n7688 585
R4775 VSS.n7822 VSS.n7821 585
R4776 VSS.n7821 VSS.n7820 585
R4777 VSS.n7680 VSS.n7677 585
R4778 VSS.n7831 VSS.n7677 585
R4779 VSS.n7837 VSS.n7836 585
R4780 VSS.n7838 VSS.n7837 585
R4781 VSS.n5482 VSS.n5481 585
R4782 VSS.n5481 VSS.n5480 585
R4783 VSS.n5492 VSS.n5491 585
R4784 VSS.n5491 VSS.n5490 585
R4785 VSS.n5473 VSS.n5469 585
R4786 VSS.n5501 VSS.n5469 585
R4787 VSS.n5465 VSS.n5462 585
R4788 VSS.n5462 VSS.n5461 585
R4789 VSS.n5515 VSS.n5514 585
R4790 VSS.n5514 VSS.n5513 585
R4791 VSS.n5454 VSS.n5450 585
R4792 VSS.n5523 VSS.n5450 585
R4793 VSS.n5446 VSS.n5443 585
R4794 VSS.n5443 VSS.n5442 585
R4795 VSS.n5537 VSS.n5536 585
R4796 VSS.n5536 VSS.n5535 585
R4797 VSS.n5435 VSS.n5431 585
R4798 VSS.n5546 VSS.n5431 585
R4799 VSS.n5427 VSS.n5424 585
R4800 VSS.n5424 VSS.n5423 585
R4801 VSS.n5560 VSS.n5559 585
R4802 VSS.n5559 VSS.n5558 585
R4803 VSS.n5568 VSS.n3688 585
R4804 VSS.n5569 VSS.n5568 585
R4805 VSS.n5413 VSS.n5412 585
R4806 VSS.n5414 VSS.n5413 585
R4807 VSS.n5405 VSS.n5404 585
R4808 VSS.n5404 VSS.n5403 585
R4809 VSS.n3705 VSS.n3704 585
R4810 VSS.n3704 VSS.n3703 585
R4811 VSS.n5387 VSS.n5386 585
R4812 VSS.n5388 VSS.n5387 585
R4813 VSS.n3715 VSS.n3714 585
R4814 VSS.n5377 VSS.n3715 585
R4815 VSS.n5370 VSS.n5369 585
R4816 VSS.n5369 VSS.n5368 585
R4817 VSS.n3726 VSS.n3725 585
R4818 VSS.n3725 VSS.n3724 585
R4819 VSS.n5353 VSS.n5352 585
R4820 VSS.n5354 VSS.n5353 585
R4821 VSS.n3736 VSS.n3735 585
R4822 VSS.n5343 VSS.n3736 585
R4823 VSS.n5335 VSS.n5334 585
R4824 VSS.n5334 VSS.n5333 585
R4825 VSS.n3747 VSS.n3746 585
R4826 VSS.n3746 VSS.n3745 585
R4827 VSS.n5318 VSS.n5317 585
R4828 VSS.n5319 VSS.n5318 585
R4829 VSS.n5128 VSS.n5124 585
R4830 VSS.n5124 VSS.n5123 585
R4831 VSS.n5146 VSS.n5145 585
R4832 VSS.n5145 VSS.n5144 585
R4833 VSS.n5116 VSS.n5112 585
R4834 VSS.n5155 VSS.n5112 585
R4835 VSS.n5108 VSS.n5105 585
R4836 VSS.n5105 VSS.n5104 585
R4837 VSS.n5169 VSS.n5168 585
R4838 VSS.n5168 VSS.n5167 585
R4839 VSS.n5097 VSS.n5093 585
R4840 VSS.n5177 VSS.n5093 585
R4841 VSS.n5089 VSS.n5086 585
R4842 VSS.n5086 VSS.n5085 585
R4843 VSS.n5191 VSS.n5190 585
R4844 VSS.n5190 VSS.n5189 585
R4845 VSS.n5078 VSS.n5074 585
R4846 VSS.n5200 VSS.n5074 585
R4847 VSS.n5070 VSS.n5067 585
R4848 VSS.n5067 VSS.n5066 585
R4849 VSS.n5214 VSS.n5213 585
R4850 VSS.n5213 VSS.n5212 585
R4851 VSS.n5222 VSS.n3829 585
R4852 VSS.n5223 VSS.n5222 585
R4853 VSS.n5056 VSS.n5055 585
R4854 VSS.n5057 VSS.n5056 585
R4855 VSS.n5048 VSS.n5047 585
R4856 VSS.n5047 VSS.n5046 585
R4857 VSS.n3846 VSS.n3845 585
R4858 VSS.n3845 VSS.n3844 585
R4859 VSS.n5030 VSS.n5029 585
R4860 VSS.n5031 VSS.n5030 585
R4861 VSS.n3856 VSS.n3855 585
R4862 VSS.n5020 VSS.n3856 585
R4863 VSS.n5013 VSS.n5012 585
R4864 VSS.n5012 VSS.n5011 585
R4865 VSS.n3867 VSS.n3866 585
R4866 VSS.n3866 VSS.n3865 585
R4867 VSS.n4996 VSS.n4995 585
R4868 VSS.n4997 VSS.n4996 585
R4869 VSS.n3877 VSS.n3876 585
R4870 VSS.n4986 VSS.n3877 585
R4871 VSS.n4978 VSS.n4977 585
R4872 VSS.n4977 VSS.n4976 585
R4873 VSS.n3888 VSS.n3887 585
R4874 VSS.n3887 VSS.n3886 585
R4875 VSS.n4961 VSS.n4960 585
R4876 VSS.n4962 VSS.n4961 585
R4877 VSS.n4771 VSS.n4767 585
R4878 VSS.n4767 VSS.n4766 585
R4879 VSS.n4789 VSS.n4788 585
R4880 VSS.n4788 VSS.n4787 585
R4881 VSS.n4759 VSS.n4755 585
R4882 VSS.n4798 VSS.n4755 585
R4883 VSS.n4751 VSS.n4748 585
R4884 VSS.n4748 VSS.n4747 585
R4885 VSS.n4812 VSS.n4811 585
R4886 VSS.n4811 VSS.n4810 585
R4887 VSS.n4740 VSS.n4736 585
R4888 VSS.n4820 VSS.n4736 585
R4889 VSS.n4732 VSS.n4729 585
R4890 VSS.n4729 VSS.n4728 585
R4891 VSS.n4834 VSS.n4833 585
R4892 VSS.n4833 VSS.n4832 585
R4893 VSS.n4721 VSS.n4717 585
R4894 VSS.n4843 VSS.n4717 585
R4895 VSS.n4713 VSS.n4710 585
R4896 VSS.n4710 VSS.n4709 585
R4897 VSS.n4857 VSS.n4856 585
R4898 VSS.n4856 VSS.n4855 585
R4899 VSS.n4865 VSS.n3970 585
R4900 VSS.n4866 VSS.n4865 585
R4901 VSS.n4699 VSS.n4698 585
R4902 VSS.n4700 VSS.n4699 585
R4903 VSS.n4691 VSS.n4690 585
R4904 VSS.n4690 VSS.n4689 585
R4905 VSS.n3987 VSS.n3986 585
R4906 VSS.n3986 VSS.n3985 585
R4907 VSS.n4673 VSS.n4672 585
R4908 VSS.n4674 VSS.n4673 585
R4909 VSS.n3997 VSS.n3996 585
R4910 VSS.n4663 VSS.n3997 585
R4911 VSS.n4656 VSS.n4655 585
R4912 VSS.n4655 VSS.n4654 585
R4913 VSS.n4008 VSS.n4007 585
R4914 VSS.n4007 VSS.n4006 585
R4915 VSS.n4639 VSS.n4638 585
R4916 VSS.n4640 VSS.n4639 585
R4917 VSS.n4018 VSS.n4017 585
R4918 VSS.n4629 VSS.n4018 585
R4919 VSS.n4621 VSS.n4620 585
R4920 VSS.n4620 VSS.n4619 585
R4921 VSS.n4029 VSS.n4028 585
R4922 VSS.n4028 VSS.n4027 585
R4923 VSS.n4604 VSS.n4603 585
R4924 VSS.n4605 VSS.n4604 585
R4925 VSS.n4414 VSS.n4410 585
R4926 VSS.n4410 VSS.n4409 585
R4927 VSS.n4432 VSS.n4431 585
R4928 VSS.n4431 VSS.n4430 585
R4929 VSS.n4402 VSS.n4398 585
R4930 VSS.n4441 VSS.n4398 585
R4931 VSS.n4394 VSS.n4391 585
R4932 VSS.n4391 VSS.n4390 585
R4933 VSS.n4455 VSS.n4454 585
R4934 VSS.n4454 VSS.n4453 585
R4935 VSS.n4383 VSS.n4379 585
R4936 VSS.n4463 VSS.n4379 585
R4937 VSS.n4375 VSS.n4372 585
R4938 VSS.n4372 VSS.n4371 585
R4939 VSS.n4477 VSS.n4476 585
R4940 VSS.n4476 VSS.n4475 585
R4941 VSS.n4364 VSS.n4360 585
R4942 VSS.n4486 VSS.n4360 585
R4943 VSS.n4356 VSS.n4353 585
R4944 VSS.n4353 VSS.n4352 585
R4945 VSS.n4500 VSS.n4499 585
R4946 VSS.n4499 VSS.n4498 585
R4947 VSS.n4508 VSS.n4111 585
R4948 VSS.n4509 VSS.n4508 585
R4949 VSS.n4342 VSS.n4341 585
R4950 VSS.n4343 VSS.n4342 585
R4951 VSS.n4334 VSS.n4333 585
R4952 VSS.n4333 VSS.n4332 585
R4953 VSS.n4128 VSS.n4127 585
R4954 VSS.n4127 VSS.n4126 585
R4955 VSS.n4316 VSS.n4315 585
R4956 VSS.n4317 VSS.n4316 585
R4957 VSS.n4138 VSS.n4137 585
R4958 VSS.n4306 VSS.n4138 585
R4959 VSS.n4299 VSS.n4298 585
R4960 VSS.n4298 VSS.n4297 585
R4961 VSS.n4149 VSS.n4148 585
R4962 VSS.n4148 VSS.n4147 585
R4963 VSS.n4282 VSS.n4281 585
R4964 VSS.n4283 VSS.n4282 585
R4965 VSS.n4159 VSS.n4158 585
R4966 VSS.n4272 VSS.n4159 585
R4967 VSS.n4264 VSS.n4263 585
R4968 VSS.n4263 VSS.n4262 585
R4969 VSS.n4170 VSS.n4169 585
R4970 VSS.n4169 VSS.n4168 585
R4971 VSS.n4247 VSS.n4246 585
R4972 VSS.n4248 VSS.n4247 585
R4973 VSS.n2882 VSS.n2881 585
R4974 VSS.n2881 VSS.n2880 585
R4975 VSS.n2868 VSS.n2864 585
R4976 VSS.n2891 VSS.n2864 585
R4977 VSS.n2860 VSS.n2857 585
R4978 VSS.n2857 VSS.n2856 585
R4979 VSS.n2905 VSS.n2904 585
R4980 VSS.n2904 VSS.n2903 585
R4981 VSS.n2849 VSS.n2845 585
R4982 VSS.n2914 VSS.n2845 585
R4983 VSS.n2841 VSS.n2838 585
R4984 VSS.n2838 VSS.n2837 585
R4985 VSS.n2927 VSS.n2926 585
R4986 VSS.n2926 VSS.n2925 585
R4987 VSS.n2830 VSS.n2826 585
R4988 VSS.n2936 VSS.n2826 585
R4989 VSS.n2822 VSS.n2819 585
R4990 VSS.n2819 VSS.n2818 585
R4991 VSS.n2950 VSS.n2949 585
R4992 VSS.n2949 VSS.n2948 585
R4993 VSS.n2811 VSS.n2805 585
R4994 VSS.n2959 VSS.n2805 585
R4995 VSS.n2806 VSS.n1312 585
R4996 VSS.n2807 VSS.n2806 585
R4997 VSS.n2792 VSS.n2791 585
R4998 VSS.n2793 VSS.n2792 585
R4999 VSS.n1322 VSS.n1321 585
R5000 VSS.n2782 VSS.n1322 585
R5001 VSS.n2774 VSS.n2773 585
R5002 VSS.n2773 VSS.n2772 585
R5003 VSS.n1333 VSS.n1332 585
R5004 VSS.n1332 VSS.n1331 585
R5005 VSS.n2757 VSS.n2756 585
R5006 VSS.n2758 VSS.n2757 585
R5007 VSS.n1343 VSS.n1342 585
R5008 VSS.n2748 VSS.n1343 585
R5009 VSS.n2740 VSS.n2739 585
R5010 VSS.n2739 VSS.n2738 585
R5011 VSS.n1354 VSS.n1353 585
R5012 VSS.n1353 VSS.n1352 585
R5013 VSS.n2723 VSS.n2722 585
R5014 VSS.n2724 VSS.n2723 585
R5015 VSS.n1364 VSS.n1363 585
R5016 VSS.n2713 VSS.n1364 585
R5017 VSS.n2705 VSS.n2704 585
R5018 VSS.n2704 VSS.n2703 585
R5019 VSS.n1375 VSS.n1374 585
R5020 VSS.n1374 VSS.n1373 585
R5021 VSS.n2688 VSS.n2687 585
R5022 VSS.n2687 VSS.n2686 585
R5023 VSS.n2391 VSS.n2389 585
R5024 VSS.n2399 VSS.n2389 585
R5025 VSS.n2385 VSS.n2382 585
R5026 VSS.n2382 VSS.n2381 585
R5027 VSS.n2413 VSS.n2412 585
R5028 VSS.n2412 VSS.n2411 585
R5029 VSS.n2374 VSS.n2370 585
R5030 VSS.n2422 VSS.n2370 585
R5031 VSS.n2366 VSS.n2363 585
R5032 VSS.n2363 VSS.n2362 585
R5033 VSS.n2435 VSS.n2434 585
R5034 VSS.n2434 VSS.n2433 585
R5035 VSS.n2355 VSS.n2351 585
R5036 VSS.n2444 VSS.n2351 585
R5037 VSS.n2347 VSS.n2344 585
R5038 VSS.n2344 VSS.n2343 585
R5039 VSS.n2458 VSS.n2457 585
R5040 VSS.n2457 VSS.n2456 585
R5041 VSS.n2336 VSS.n2329 585
R5042 VSS.n2467 VSS.n2329 585
R5043 VSS.n2331 VSS.n2330 585
R5044 VSS.n2332 VSS.n2331 585
R5045 VSS.n2482 VSS.n2481 585
R5046 VSS.n2481 VSS.n2480 585
R5047 VSS.n2281 VSS.n2277 585
R5048 VSS.n2491 VSS.n2277 585
R5049 VSS.n2273 VSS.n2270 585
R5050 VSS.n2270 VSS.n2269 585
R5051 VSS.n2505 VSS.n2504 585
R5052 VSS.n2504 VSS.n2503 585
R5053 VSS.n2262 VSS.n2258 585
R5054 VSS.n2514 VSS.n2258 585
R5055 VSS.n2254 VSS.n2251 585
R5056 VSS.n2251 VSS.n2250 585
R5057 VSS.n2527 VSS.n2526 585
R5058 VSS.n2526 VSS.n2525 585
R5059 VSS.n2243 VSS.n2239 585
R5060 VSS.n2536 VSS.n2239 585
R5061 VSS.n2235 VSS.n2232 585
R5062 VSS.n2232 VSS.n2231 585
R5063 VSS.n2550 VSS.n2549 585
R5064 VSS.n2549 VSS.n2548 585
R5065 VSS.n2224 VSS.n2220 585
R5066 VSS.n2559 VSS.n2220 585
R5067 VSS.n2218 VSS.n2217 585
R5068 VSS.n2218 VSS.n1479 585
R5069 VSS.n2211 VSS.n2210 585
R5070 VSS.n2210 VSS.n2209 585
R5071 VSS.n1489 VSS.n1488 585
R5072 VSS.n1488 VSS.n1487 585
R5073 VSS.n2194 VSS.n2193 585
R5074 VSS.n2195 VSS.n2194 585
R5075 VSS.n1499 VSS.n1498 585
R5076 VSS.n2184 VSS.n1499 585
R5077 VSS.n2176 VSS.n2175 585
R5078 VSS.n2175 VSS.n2174 585
R5079 VSS.n1510 VSS.n1509 585
R5080 VSS.n1509 VSS.n1508 585
R5081 VSS.n2160 VSS.n2159 585
R5082 VSS.n2161 VSS.n2160 585
R5083 VSS.n1520 VSS.n1519 585
R5084 VSS.n2150 VSS.n1520 585
R5085 VSS.n2142 VSS.n2141 585
R5086 VSS.n2141 VSS.n2140 585
R5087 VSS.n1531 VSS.n1530 585
R5088 VSS.n1530 VSS.n1529 585
R5089 VSS.n2125 VSS.n2124 585
R5090 VSS.n2126 VSS.n2125 585
R5091 VSS.n1541 VSS.n1540 585
R5092 VSS.n2115 VSS.n1541 585
R5093 VSS.n1787 VSS.n1786 585
R5094 VSS.n1786 VSS.n1785 585
R5095 VSS.n1784 VSS.n1780 585
R5096 VSS.n1798 VSS.n1780 585
R5097 VSS.n1776 VSS.n1773 585
R5098 VSS.n1773 VSS.n1772 585
R5099 VSS.n1812 VSS.n1811 585
R5100 VSS.n1811 VSS.n1810 585
R5101 VSS.n1765 VSS.n1761 585
R5102 VSS.n1821 VSS.n1761 585
R5103 VSS.n1757 VSS.n1754 585
R5104 VSS.n1754 VSS.n1753 585
R5105 VSS.n1834 VSS.n1833 585
R5106 VSS.n1833 VSS.n1832 585
R5107 VSS.n1746 VSS.n1742 585
R5108 VSS.n1843 VSS.n1742 585
R5109 VSS.n1738 VSS.n1735 585
R5110 VSS.n1735 VSS.n1734 585
R5111 VSS.n1857 VSS.n1856 585
R5112 VSS.n1856 VSS.n1855 585
R5113 VSS.n1727 VSS.n1720 585
R5114 VSS.n1866 VSS.n1720 585
R5115 VSS.n1722 VSS.n1721 585
R5116 VSS.n1723 VSS.n1722 585
R5117 VSS.n1881 VSS.n1880 585
R5118 VSS.n1880 VSS.n1879 585
R5119 VSS.n1672 VSS.n1668 585
R5120 VSS.n1890 VSS.n1668 585
R5121 VSS.n1664 VSS.n1661 585
R5122 VSS.n1661 VSS.n1660 585
R5123 VSS.n1904 VSS.n1903 585
R5124 VSS.n1903 VSS.n1902 585
R5125 VSS.n1653 VSS.n1649 585
R5126 VSS.n1913 VSS.n1649 585
R5127 VSS.n1645 VSS.n1642 585
R5128 VSS.n1642 VSS.n1641 585
R5129 VSS.n1926 VSS.n1925 585
R5130 VSS.n1925 VSS.n1924 585
R5131 VSS.n1634 VSS.n1630 585
R5132 VSS.n1935 VSS.n1630 585
R5133 VSS.n1626 VSS.n1623 585
R5134 VSS.n1623 VSS.n1622 585
R5135 VSS.n1949 VSS.n1948 585
R5136 VSS.n1948 VSS.n1947 585
R5137 VSS.n1614 VSS.n1611 585
R5138 VSS.n1958 VSS.n1611 585
R5139 VSS.n1964 VSS.n1963 585
R5140 VSS.n1965 VSS.n1964 585
R5141 VSS.n15945 VSS.n15944 575.163
R5142 VSS.n15919 VSS.n14056 575.163
R5143 VSS.n15414 VSS.n15413 575.163
R5144 VSS.n15389 VSS.n14206 575.163
R5145 VSS.n14811 VSS.n14221 575.163
R5146 VSS.n14836 VSS.n14835 575.163
R5147 VSS.n14775 VSS.n14774 575.163
R5148 VSS.n12160 VSS.n12159 575.163
R5149 VSS.n12437 VSS.n11526 575.163
R5150 VSS.n12464 VSS.n12463 575.163
R5151 VSS.n13370 VSS.n13369 575.163
R5152 VSS.n13345 VSS.n13344 575.163
R5153 VSS.n13121 VSS.n13120 575.163
R5154 VSS.n13096 VSS.n13095 575.163
R5155 VSS.n8825 VSS.n6979 575.163
R5156 VSS.n8800 VSS.n8799 575.163
R5157 VSS.n8603 VSS.n7335 575.163
R5158 VSS.n8578 VSS.n8577 575.163
R5159 VSS.n8245 VSS.n7475 575.163
R5160 VSS.n8220 VSS.n8219 575.163
R5161 VSS.n7887 VSS.n7615 575.163
R5162 VSS.n5609 VSS.n5608 575.163
R5163 VSS.n5288 VSS.n5287 575.163
R5164 VSS.n5263 VSS.n5262 575.163
R5165 VSS.n4931 VSS.n4930 575.163
R5166 VSS.n4906 VSS.n4905 575.163
R5167 VSS.n4574 VSS.n4573 575.163
R5168 VSS.n4549 VSS.n4548 575.163
R5169 VSS.n2993 VSS.n1297 575.163
R5170 VSS.n2655 VSS.n2654 575.163
R5171 VSS.n2630 VSS.n1447 575.163
R5172 VSS.n2052 VSS.n1462 575.163
R5173 VSS.n2077 VSS.n2076 575.163
R5174 VSS.n2016 VSS.n2015 575.163
R5175 VSS.n15678 VSS.n15634 488.888
R5176 VSS.n15566 VSS.n14069 488.888
R5177 VSS.n14144 VSS.n14132 488.888
R5178 VSS.n15091 VSS.n15047 488.888
R5179 VSS.n15331 VSS.n14238 488.888
R5180 VSS.n14874 VSS.n14873 488.888
R5181 VSS.n14482 VSS.n14438 488.888
R5182 VSS.n11992 VSS.n11981 488.888
R5183 VSS.n12406 VSS.n11543 488.888
R5184 VSS.n11808 VSS.n11807 488.888
R5185 VSS.n11673 VSS.n11485 488.888
R5186 VSS.n13306 VSS.n13305 488.888
R5187 VSS.n13152 VSS.n12581 488.888
R5188 VSS.n13057 VSS.n13056 488.888
R5189 VSS.n8856 VSS.n6965 488.888
R5190 VSS.n8772 VSS.n7256 488.888
R5191 VSS.n8635 VSS.n8634 488.888
R5192 VSS.n8550 VSS.n7396 488.888
R5193 VSS.n8277 VSS.n8276 488.888
R5194 VSS.n8192 VSS.n7536 488.888
R5195 VSS.n7919 VSS.n7918 488.888
R5196 VSS.n5570 VSS.n5569 488.888
R5197 VSS.n5319 VSS.n3752 488.888
R5198 VSS.n5224 VSS.n5223 488.888
R5199 VSS.n4962 VSS.n3893 488.888
R5200 VSS.n4867 VSS.n4866 488.888
R5201 VSS.n4605 VSS.n4034 488.888
R5202 VSS.n4510 VSS.n4509 488.888
R5203 VSS.n2807 VSS.n1310 488.888
R5204 VSS.n1385 VSS.n1373 488.888
R5205 VSS.n2332 VSS.n2288 488.888
R5206 VSS.n2572 VSS.n1479 488.888
R5207 VSS.n2115 VSS.n2114 488.888
R5208 VSS.n1723 VSS.n1679 488.888
R5209 VSS.n15667 VSS.n15634 345.098
R5210 VSS.n15894 VSS.n14069 345.098
R5211 VSS.n15439 VSS.n14144 345.098
R5212 VSS.n15080 VSS.n15047 345.098
R5213 VSS.n15332 VSS.n15331 345.098
R5214 VSS.n14873 VSS.n14301 345.098
R5215 VSS.n14471 VSS.n14438 345.098
R5216 VSS.n12102 VSS.n11981 345.098
R5217 VSS.n12407 VSS.n12406 345.098
R5218 VSS.n11807 VSS.n11806 345.098
R5219 VSS.n13395 VSS.n11485 345.098
R5220 VSS.n13306 VSS.n12515 345.098
R5221 VSS.n13146 VSS.n12581 345.098
R5222 VSS.n13057 VSS.n12656 345.098
R5223 VSS.n8856 VSS.n8855 345.098
R5224 VSS.n8773 VSS.n8772 345.098
R5225 VSS.n8634 VSS.n8633 345.098
R5226 VSS.n8551 VSS.n8550 345.098
R5227 VSS.n8276 VSS.n8275 345.098
R5228 VSS.n8193 VSS.n8192 345.098
R5229 VSS.n7918 VSS.n7917 345.098
R5230 VSS.n5570 VSS.n3686 345.098
R5231 VSS.n5313 VSS.n3752 345.098
R5232 VSS.n5224 VSS.n3827 345.098
R5233 VSS.n4956 VSS.n3893 345.098
R5234 VSS.n4867 VSS.n3968 345.098
R5235 VSS.n4599 VSS.n4034 345.098
R5236 VSS.n4510 VSS.n4109 345.098
R5237 VSS.n2968 VSS.n1310 345.098
R5238 VSS.n2680 VSS.n1385 345.098
R5239 VSS.n2321 VSS.n2288 345.098
R5240 VSS.n2573 VSS.n2572 345.098
R5241 VSS.n2114 VSS.n1542 345.098
R5242 VSS.n1712 VSS.n1679 345.098
R5243 VSS.n10436 VSS.n10435 321.976
R5244 VSS.n14725 VSS.n14364 321.258
R5245 VSS.n12790 VSS.n12722 321.258
R5246 VSS.n7840 VSS.n7839 321.258
R5247 VSS.n6828 VSS.n6758 321.258
R5248 VSS.n4243 VSS.n4175 321.258
R5249 VSS.n1966 VSS.n1605 321.258
R5250 VSS.n14728 VSS.n14727 292.5
R5251 VSS.n14727 VSS.n14726 292.5
R5252 VSS.n14351 VSS.n14350 292.5
R5253 VSS.n14749 VSS.n14351 292.5
R5254 VSS.n14747 VSS.n14746 292.5
R5255 VSS.n14748 VSS.n14747 292.5
R5256 VSS.n14745 VSS.n14353 292.5
R5257 VSS.n14353 VSS.n14352 292.5
R5258 VSS.n14744 VSS.n14743 292.5
R5259 VSS.n14743 VSS.n14742 292.5
R5260 VSS.n14355 VSS.n14354 292.5
R5261 VSS.n14741 VSS.n14355 292.5
R5262 VSS.n14739 VSS.n14738 292.5
R5263 VSS.n14740 VSS.n14739 292.5
R5264 VSS.n14737 VSS.n14357 292.5
R5265 VSS.n14357 VSS.n14356 292.5
R5266 VSS.n14736 VSS.n14735 292.5
R5267 VSS.n14735 VSS.n14734 292.5
R5268 VSS.n14359 VSS.n14358 292.5
R5269 VSS.n14733 VSS.n14359 292.5
R5270 VSS.n14731 VSS.n14730 292.5
R5271 VSS.n14732 VSS.n14731 292.5
R5272 VSS.n14729 VSS.n14361 292.5
R5273 VSS.n14361 VSS.n14360 292.5
R5274 VSS.n14010 VSS.n14009 292.5
R5275 VSS.n16006 VSS.n14010 292.5
R5276 VSS.n14014 VSS.n14012 292.5
R5277 VSS.n14012 VSS.n14011 292.5
R5278 VSS.n15674 VSS.n15672 292.5
R5279 VSS.n15679 VSS.n15674 292.5
R5280 VSS.n15791 VSS.n15790 292.5
R5281 VSS.n15792 VSS.n15791 292.5
R5282 VSS.n15688 VSS.n15687 292.5
R5283 VSS.n15781 VSS.n15688 292.5
R5284 VSS.n15696 VSS.n15694 292.5
R5285 VSS.n15698 VSS.n15696 292.5
R5286 VSS.n15768 VSS.n15767 292.5
R5287 VSS.n15769 VSS.n15768 292.5
R5288 VSS.n15707 VSS.n15706 292.5
R5289 VSS.n15758 VSS.n15707 292.5
R5290 VSS.n15715 VSS.n15713 292.5
R5291 VSS.n15717 VSS.n15715 292.5
R5292 VSS.n15746 VSS.n15745 292.5
R5293 VSS.n15747 VSS.n15746 292.5
R5294 VSS.n15726 VSS.n15725 292.5
R5295 VSS.n15736 VSS.n15726 292.5
R5296 VSS.n13999 VSS.n13997 292.5
R5297 VSS.n14001 VSS.n13999 292.5
R5298 VSS.n16016 VSS.n16015 292.5
R5299 VSS.n16017 VSS.n16016 292.5
R5300 VSS.n14016 VSS.n14015 292.5
R5301 VSS.n15994 VSS.n14016 292.5
R5302 VSS.n15992 VSS.n15991 292.5
R5303 VSS.n15993 VSS.n15992 292.5
R5304 VSS.n15990 VSS.n14018 292.5
R5305 VSS.n14018 VSS.n14017 292.5
R5306 VSS.n15989 VSS.n15988 292.5
R5307 VSS.n15988 VSS.n15987 292.5
R5308 VSS.n14020 VSS.n14019 292.5
R5309 VSS.n15986 VSS.n14020 292.5
R5310 VSS.n15984 VSS.n15983 292.5
R5311 VSS.n15985 VSS.n15984 292.5
R5312 VSS.n15982 VSS.n14022 292.5
R5313 VSS.n14022 VSS.n14021 292.5
R5314 VSS.n15981 VSS.n15980 292.5
R5315 VSS.n15980 VSS.n15979 292.5
R5316 VSS.n14024 VSS.n14023 292.5
R5317 VSS.n15978 VSS.n14024 292.5
R5318 VSS.n15976 VSS.n15975 292.5
R5319 VSS.n15977 VSS.n15976 292.5
R5320 VSS.n15974 VSS.n14026 292.5
R5321 VSS.n14026 VSS.n14025 292.5
R5322 VSS.n15997 VSS.n15996 292.5
R5323 VSS.n15996 VSS.n15995 292.5
R5324 VSS.n15950 VSS.n14038 292.5
R5325 VSS.n14038 VSS.n14037 292.5
R5326 VSS.n15952 VSS.n15951 292.5
R5327 VSS.n15953 VSS.n15952 292.5
R5328 VSS.n14036 VSS.n14035 292.5
R5329 VSS.n15954 VSS.n14036 292.5
R5330 VSS.n15957 VSS.n15956 292.5
R5331 VSS.n15956 VSS.n15955 292.5
R5332 VSS.n15958 VSS.n14034 292.5
R5333 VSS.n14034 VSS.n14033 292.5
R5334 VSS.n15960 VSS.n15959 292.5
R5335 VSS.n15961 VSS.n15960 292.5
R5336 VSS.n14032 VSS.n14031 292.5
R5337 VSS.n15962 VSS.n14032 292.5
R5338 VSS.n15965 VSS.n15964 292.5
R5339 VSS.n15964 VSS.n15963 292.5
R5340 VSS.n15966 VSS.n14030 292.5
R5341 VSS.n14030 VSS.n14029 292.5
R5342 VSS.n15968 VSS.n15967 292.5
R5343 VSS.n15969 VSS.n15968 292.5
R5344 VSS.n14028 VSS.n14027 292.5
R5345 VSS.n15970 VSS.n14028 292.5
R5346 VSS.n15973 VSS.n15972 292.5
R5347 VSS.n15972 VSS.n15971 292.5
R5348 VSS.n15922 VSS.n15921 292.5
R5349 VSS.n15921 VSS.n15920 292.5
R5350 VSS.n15923 VSS.n14053 292.5
R5351 VSS.n14053 VSS.n14052 292.5
R5352 VSS.n15925 VSS.n15924 292.5
R5353 VSS.n15926 VSS.n15925 292.5
R5354 VSS.n14051 VSS.n14050 292.5
R5355 VSS.n15927 VSS.n14051 292.5
R5356 VSS.n15930 VSS.n15929 292.5
R5357 VSS.n15929 VSS.n15928 292.5
R5358 VSS.n15931 VSS.n14049 292.5
R5359 VSS.n14049 VSS.n14048 292.5
R5360 VSS.n15933 VSS.n15932 292.5
R5361 VSS.n15934 VSS.n15933 292.5
R5362 VSS.n14047 VSS.n14046 292.5
R5363 VSS.n15935 VSS.n14047 292.5
R5364 VSS.n15939 VSS.n15938 292.5
R5365 VSS.n15938 VSS.n15937 292.5
R5366 VSS.n15940 VSS.n14045 292.5
R5367 VSS.n15936 VSS.n14045 292.5
R5368 VSS.n15942 VSS.n15941 292.5
R5369 VSS.n15942 VSS.n14044 292.5
R5370 VSS.n15943 VSS.n14039 292.5
R5371 VSS.n15944 VSS.n15943 292.5
R5372 VSS.n15633 VSS.n15632 292.5
R5373 VSS.n15805 VSS.n15633 292.5
R5374 VSS.n15815 VSS.n15814 292.5
R5375 VSS.n15816 VSS.n15815 292.5
R5376 VSS.n15622 VSS.n15620 292.5
R5377 VSS.n15624 VSS.n15622 292.5
R5378 VSS.n15614 VSS.n15613 292.5
R5379 VSS.n15828 VSS.n15614 292.5
R5380 VSS.n15838 VSS.n15837 292.5
R5381 VSS.n15839 VSS.n15838 292.5
R5382 VSS.n15603 VSS.n15601 292.5
R5383 VSS.n15605 VSS.n15603 292.5
R5384 VSS.n15595 VSS.n15594 292.5
R5385 VSS.n15850 VSS.n15595 292.5
R5386 VSS.n15860 VSS.n15859 292.5
R5387 VSS.n15861 VSS.n15860 292.5
R5388 VSS.n15584 VSS.n15582 292.5
R5389 VSS.n15586 VSS.n15584 292.5
R5390 VSS.n15576 VSS.n15575 292.5
R5391 VSS.n15873 VSS.n15576 292.5
R5392 VSS.n15883 VSS.n15882 292.5
R5393 VSS.n15884 VSS.n15883 292.5
R5394 VSS.n15563 VSS.n15561 292.5
R5395 VSS.n15567 VSS.n15563 292.5
R5396 VSS.n14075 VSS.n14074 292.5
R5397 VSS.n15553 VSS.n14075 292.5
R5398 VSS.n15544 VSS.n15543 292.5
R5399 VSS.n15543 VSS.n15542 292.5
R5400 VSS.n14084 VSS.n14083 292.5
R5401 VSS.n14083 VSS.n14082 292.5
R5402 VSS.n15528 VSS.n15527 292.5
R5403 VSS.n15529 VSS.n15528 292.5
R5404 VSS.n14096 VSS.n14094 292.5
R5405 VSS.n15518 VSS.n14096 292.5
R5406 VSS.n15510 VSS.n15509 292.5
R5407 VSS.n15509 VSS.n15508 292.5
R5408 VSS.n14105 VSS.n14104 292.5
R5409 VSS.n14104 VSS.n14103 292.5
R5410 VSS.n15494 VSS.n15493 292.5
R5411 VSS.n15495 VSS.n15494 292.5
R5412 VSS.n14117 VSS.n14115 292.5
R5413 VSS.n15484 VSS.n14117 292.5
R5414 VSS.n15475 VSS.n15474 292.5
R5415 VSS.n15474 VSS.n15473 292.5
R5416 VSS.n14126 VSS.n14125 292.5
R5417 VSS.n14125 VSS.n14124 292.5
R5418 VSS.n15459 VSS.n15458 292.5
R5419 VSS.n15460 VSS.n15459 292.5
R5420 VSS.n14192 VSS.n14191 292.5
R5421 VSS.n14193 VSS.n14192 292.5
R5422 VSS.n14190 VSS.n14160 292.5
R5423 VSS.n14160 VSS.n14159 292.5
R5424 VSS.n14189 VSS.n14188 292.5
R5425 VSS.n14188 VSS.n14187 292.5
R5426 VSS.n14162 VSS.n14161 292.5
R5427 VSS.n14186 VSS.n14162 292.5
R5428 VSS.n14184 VSS.n14183 292.5
R5429 VSS.n14185 VSS.n14184 292.5
R5430 VSS.n14182 VSS.n14164 292.5
R5431 VSS.n14164 VSS.n14163 292.5
R5432 VSS.n14181 VSS.n14180 292.5
R5433 VSS.n14180 VSS.n14179 292.5
R5434 VSS.n14166 VSS.n14165 292.5
R5435 VSS.n14178 VSS.n14166 292.5
R5436 VSS.n14176 VSS.n14175 292.5
R5437 VSS.n14177 VSS.n14176 292.5
R5438 VSS.n14174 VSS.n14168 292.5
R5439 VSS.n14168 VSS.n14167 292.5
R5440 VSS.n14173 VSS.n14172 292.5
R5441 VSS.n14172 VSS.n14171 292.5
R5442 VSS.n14170 VSS.n14169 292.5
R5443 VSS.n14170 VSS.n14056 292.5
R5444 VSS.n14205 VSS.n14204 292.5
R5445 VSS.n15390 VSS.n14205 292.5
R5446 VSS.n15393 VSS.n15392 292.5
R5447 VSS.n15392 VSS.n15391 292.5
R5448 VSS.n15394 VSS.n14203 292.5
R5449 VSS.n14203 VSS.n14202 292.5
R5450 VSS.n15396 VSS.n15395 292.5
R5451 VSS.n15397 VSS.n15396 292.5
R5452 VSS.n14201 VSS.n14200 292.5
R5453 VSS.n15398 VSS.n14201 292.5
R5454 VSS.n15401 VSS.n15400 292.5
R5455 VSS.n15400 VSS.n15399 292.5
R5456 VSS.n15402 VSS.n14199 292.5
R5457 VSS.n14199 VSS.n14198 292.5
R5458 VSS.n15404 VSS.n15403 292.5
R5459 VSS.n15405 VSS.n15404 292.5
R5460 VSS.n14197 VSS.n14196 292.5
R5461 VSS.n15406 VSS.n14197 292.5
R5462 VSS.n15409 VSS.n15408 292.5
R5463 VSS.n15408 VSS.n15407 292.5
R5464 VSS.n15410 VSS.n14195 292.5
R5465 VSS.n14195 VSS.n14194 292.5
R5466 VSS.n15412 VSS.n15411 292.5
R5467 VSS.n15413 VSS.n15412 292.5
R5468 VSS.n14142 VSS.n14140 292.5
R5469 VSS.n15444 VSS.n14142 292.5
R5470 VSS.n15156 VSS.n15155 292.5
R5471 VSS.n15157 VSS.n15156 292.5
R5472 VSS.n15147 VSS.n15145 292.5
R5473 VSS.n15149 VSS.n15147 292.5
R5474 VSS.n15139 VSS.n15138 292.5
R5475 VSS.n15169 VSS.n15139 292.5
R5476 VSS.n15179 VSS.n15178 292.5
R5477 VSS.n15180 VSS.n15179 292.5
R5478 VSS.n15128 VSS.n15126 292.5
R5479 VSS.n15130 VSS.n15128 292.5
R5480 VSS.n15120 VSS.n15119 292.5
R5481 VSS.n15191 VSS.n15120 292.5
R5482 VSS.n15201 VSS.n15200 292.5
R5483 VSS.n15202 VSS.n15201 292.5
R5484 VSS.n15109 VSS.n15107 292.5
R5485 VSS.n15111 VSS.n15109 292.5
R5486 VSS.n15101 VSS.n15100 292.5
R5487 VSS.n15214 VSS.n15101 292.5
R5488 VSS.n15224 VSS.n15223 292.5
R5489 VSS.n15225 VSS.n15224 292.5
R5490 VSS.n15087 VSS.n15085 292.5
R5491 VSS.n15092 VSS.n15087 292.5
R5492 VSS.n15046 VSS.n15045 292.5
R5493 VSS.n15238 VSS.n15046 292.5
R5494 VSS.n15248 VSS.n15247 292.5
R5495 VSS.n15249 VSS.n15248 292.5
R5496 VSS.n15035 VSS.n15033 292.5
R5497 VSS.n15037 VSS.n15035 292.5
R5498 VSS.n15027 VSS.n15026 292.5
R5499 VSS.n15261 VSS.n15027 292.5
R5500 VSS.n15271 VSS.n15270 292.5
R5501 VSS.n15272 VSS.n15271 292.5
R5502 VSS.n15016 VSS.n15014 292.5
R5503 VSS.n15018 VSS.n15016 292.5
R5504 VSS.n15008 VSS.n15007 292.5
R5505 VSS.n15283 VSS.n15008 292.5
R5506 VSS.n15293 VSS.n15292 292.5
R5507 VSS.n15294 VSS.n15293 292.5
R5508 VSS.n14997 VSS.n14995 292.5
R5509 VSS.n14999 VSS.n14997 292.5
R5510 VSS.n14989 VSS.n14988 292.5
R5511 VSS.n15306 VSS.n14989 292.5
R5512 VSS.n15316 VSS.n15315 292.5
R5513 VSS.n15317 VSS.n15316 292.5
R5514 VSS.n14978 VSS.n14974 292.5
R5515 VSS.n14980 VSS.n14978 292.5
R5516 VSS.n15361 VSS.n15360 292.5
R5517 VSS.n15362 VSS.n15361 292.5
R5518 VSS.n14220 VSS.n14219 292.5
R5519 VSS.n15363 VSS.n14220 292.5
R5520 VSS.n15366 VSS.n15365 292.5
R5521 VSS.n15365 VSS.n15364 292.5
R5522 VSS.n15367 VSS.n14218 292.5
R5523 VSS.n14218 VSS.n14217 292.5
R5524 VSS.n15369 VSS.n15368 292.5
R5525 VSS.n15370 VSS.n15369 292.5
R5526 VSS.n14216 VSS.n14215 292.5
R5527 VSS.n15371 VSS.n14216 292.5
R5528 VSS.n15374 VSS.n15373 292.5
R5529 VSS.n15373 VSS.n15372 292.5
R5530 VSS.n15375 VSS.n14214 292.5
R5531 VSS.n14214 VSS.n14213 292.5
R5532 VSS.n15378 VSS.n15377 292.5
R5533 VSS.n15379 VSS.n15378 292.5
R5534 VSS.n15376 VSS.n14212 292.5
R5535 VSS.n15380 VSS.n14212 292.5
R5536 VSS.n15382 VSS.n14211 292.5
R5537 VSS.n15382 VSS.n15381 292.5
R5538 VSS.n15384 VSS.n15383 292.5
R5539 VSS.n15383 VSS.n14206 292.5
R5540 VSS.n14833 VSS.n14321 292.5
R5541 VSS.n14834 VSS.n14833 292.5
R5542 VSS.n14832 VSS.n14831 292.5
R5543 VSS.n14832 VSS.n14801 292.5
R5544 VSS.n14830 VSS.n14802 292.5
R5545 VSS.n14805 VSS.n14802 292.5
R5546 VSS.n14829 VSS.n14828 292.5
R5547 VSS.n14828 VSS.n14827 292.5
R5548 VSS.n14804 VSS.n14803 292.5
R5549 VSS.n14826 VSS.n14804 292.5
R5550 VSS.n14824 VSS.n14823 292.5
R5551 VSS.n14825 VSS.n14824 292.5
R5552 VSS.n14822 VSS.n14807 292.5
R5553 VSS.n14807 VSS.n14806 292.5
R5554 VSS.n14821 VSS.n14820 292.5
R5555 VSS.n14820 VSS.n14819 292.5
R5556 VSS.n14809 VSS.n14808 292.5
R5557 VSS.n14818 VSS.n14809 292.5
R5558 VSS.n14816 VSS.n14815 292.5
R5559 VSS.n14817 VSS.n14816 292.5
R5560 VSS.n14814 VSS.n14813 292.5
R5561 VSS.n14813 VSS.n14810 292.5
R5562 VSS.n14812 VSS.n14223 292.5
R5563 VSS.n14812 VSS.n14811 292.5
R5564 VSS.n14241 VSS.n14240 292.5
R5565 VSS.n14240 VSS.n14239 292.5
R5566 VSS.n14965 VSS.n14964 292.5
R5567 VSS.n14966 VSS.n14965 292.5
R5568 VSS.n14252 VSS.n14250 292.5
R5569 VSS.n14955 VSS.n14252 292.5
R5570 VSS.n14946 VSS.n14945 292.5
R5571 VSS.n14945 VSS.n14944 292.5
R5572 VSS.n14261 VSS.n14260 292.5
R5573 VSS.n14260 VSS.n14259 292.5
R5574 VSS.n14930 VSS.n14929 292.5
R5575 VSS.n14931 VSS.n14930 292.5
R5576 VSS.n14273 VSS.n14271 292.5
R5577 VSS.n14921 VSS.n14273 292.5
R5578 VSS.n14912 VSS.n14911 292.5
R5579 VSS.n14911 VSS.n14910 292.5
R5580 VSS.n14282 VSS.n14281 292.5
R5581 VSS.n14281 VSS.n14280 292.5
R5582 VSS.n14896 VSS.n14895 292.5
R5583 VSS.n14897 VSS.n14896 292.5
R5584 VSS.n14294 VSS.n14292 292.5
R5585 VSS.n14886 VSS.n14294 292.5
R5586 VSS.n14877 VSS.n14876 292.5
R5587 VSS.n14876 VSS.n14875 292.5
R5588 VSS.n14305 VSS.n14303 292.5
R5589 VSS.n14303 VSS.n14302 292.5
R5590 VSS.n14555 VSS.n14554 292.5
R5591 VSS.n14556 VSS.n14555 292.5
R5592 VSS.n14538 VSS.n14536 292.5
R5593 VSS.n14540 VSS.n14538 292.5
R5594 VSS.n14530 VSS.n14529 292.5
R5595 VSS.n14568 VSS.n14530 292.5
R5596 VSS.n14578 VSS.n14577 292.5
R5597 VSS.n14579 VSS.n14578 292.5
R5598 VSS.n14519 VSS.n14517 292.5
R5599 VSS.n14521 VSS.n14519 292.5
R5600 VSS.n14511 VSS.n14510 292.5
R5601 VSS.n14590 VSS.n14511 292.5
R5602 VSS.n14600 VSS.n14599 292.5
R5603 VSS.n14601 VSS.n14600 292.5
R5604 VSS.n14500 VSS.n14498 292.5
R5605 VSS.n14502 VSS.n14500 292.5
R5606 VSS.n14492 VSS.n14491 292.5
R5607 VSS.n14613 VSS.n14492 292.5
R5608 VSS.n14623 VSS.n14622 292.5
R5609 VSS.n14624 VSS.n14623 292.5
R5610 VSS.n14478 VSS.n14476 292.5
R5611 VSS.n14483 VSS.n14478 292.5
R5612 VSS.n14780 VSS.n14334 292.5
R5613 VSS.n14334 VSS.n14333 292.5
R5614 VSS.n14782 VSS.n14781 292.5
R5615 VSS.n14783 VSS.n14782 292.5
R5616 VSS.n14332 VSS.n14331 292.5
R5617 VSS.n14784 VSS.n14332 292.5
R5618 VSS.n14787 VSS.n14786 292.5
R5619 VSS.n14786 VSS.n14785 292.5
R5620 VSS.n14788 VSS.n14330 292.5
R5621 VSS.n14330 VSS.n14329 292.5
R5622 VSS.n14790 VSS.n14789 292.5
R5623 VSS.n14791 VSS.n14790 292.5
R5624 VSS.n14328 VSS.n14327 292.5
R5625 VSS.n14792 VSS.n14328 292.5
R5626 VSS.n14795 VSS.n14794 292.5
R5627 VSS.n14794 VSS.n14793 292.5
R5628 VSS.n14796 VSS.n14326 292.5
R5629 VSS.n14326 VSS.n14325 292.5
R5630 VSS.n14798 VSS.n14797 292.5
R5631 VSS.n14799 VSS.n14798 292.5
R5632 VSS.n14323 VSS.n14322 292.5
R5633 VSS.n14800 VSS.n14323 292.5
R5634 VSS.n14838 VSS.n14837 292.5
R5635 VSS.n14837 VSS.n14836 292.5
R5636 VSS.n14753 VSS.n14349 292.5
R5637 VSS.n14349 VSS.n14348 292.5
R5638 VSS.n14755 VSS.n14754 292.5
R5639 VSS.n14756 VSS.n14755 292.5
R5640 VSS.n14347 VSS.n14346 292.5
R5641 VSS.n14757 VSS.n14347 292.5
R5642 VSS.n14760 VSS.n14759 292.5
R5643 VSS.n14759 VSS.n14758 292.5
R5644 VSS.n14761 VSS.n14345 292.5
R5645 VSS.n14345 VSS.n14344 292.5
R5646 VSS.n14763 VSS.n14762 292.5
R5647 VSS.n14764 VSS.n14763 292.5
R5648 VSS.n14343 VSS.n14342 292.5
R5649 VSS.n14765 VSS.n14343 292.5
R5650 VSS.n14769 VSS.n14768 292.5
R5651 VSS.n14768 VSS.n14767 292.5
R5652 VSS.n14770 VSS.n14341 292.5
R5653 VSS.n14766 VSS.n14341 292.5
R5654 VSS.n14772 VSS.n14771 292.5
R5655 VSS.n14772 VSS.n14340 292.5
R5656 VSS.n14773 VSS.n14335 292.5
R5657 VSS.n14774 VSS.n14773 292.5
R5658 VSS.n14752 VSS.n14751 292.5
R5659 VSS.n14751 VSS.n14750 292.5
R5660 VSS.n14437 VSS.n14436 292.5
R5661 VSS.n14637 VSS.n14437 292.5
R5662 VSS.n14647 VSS.n14646 292.5
R5663 VSS.n14648 VSS.n14647 292.5
R5664 VSS.n14426 VSS.n14424 292.5
R5665 VSS.n14428 VSS.n14426 292.5
R5666 VSS.n14418 VSS.n14417 292.5
R5667 VSS.n14660 VSS.n14418 292.5
R5668 VSS.n14670 VSS.n14669 292.5
R5669 VSS.n14671 VSS.n14670 292.5
R5670 VSS.n14407 VSS.n14405 292.5
R5671 VSS.n14409 VSS.n14407 292.5
R5672 VSS.n14399 VSS.n14398 292.5
R5673 VSS.n14682 VSS.n14399 292.5
R5674 VSS.n14692 VSS.n14691 292.5
R5675 VSS.n14693 VSS.n14692 292.5
R5676 VSS.n14388 VSS.n14386 292.5
R5677 VSS.n14390 VSS.n14388 292.5
R5678 VSS.n14380 VSS.n14379 292.5
R5679 VSS.n14705 VSS.n14380 292.5
R5680 VSS.n14715 VSS.n14714 292.5
R5681 VSS.n14716 VSS.n14715 292.5
R5682 VSS.n14721 VSS.n14366 292.5
R5683 VSS.n14366 VSS.n14365 292.5
R5684 VSS.n14364 VSS.n14362 292.5
R5685 VSS.n12789 VSS.n12788 292.5
R5686 VSS.n12788 VSS.n12725 292.5
R5687 VSS.n12767 VSS.n12766 292.5
R5688 VSS.n12768 VSS.n12767 292.5
R5689 VSS.n12735 VSS.n12734 292.5
R5690 VSS.n12769 VSS.n12735 292.5
R5691 VSS.n12772 VSS.n12771 292.5
R5692 VSS.n12771 VSS.n12770 292.5
R5693 VSS.n12773 VSS.n12733 292.5
R5694 VSS.n12733 VSS.n12732 292.5
R5695 VSS.n12775 VSS.n12774 292.5
R5696 VSS.n12776 VSS.n12775 292.5
R5697 VSS.n12731 VSS.n12730 292.5
R5698 VSS.n12777 VSS.n12731 292.5
R5699 VSS.n12780 VSS.n12779 292.5
R5700 VSS.n12779 VSS.n12778 292.5
R5701 VSS.n12781 VSS.n12728 292.5
R5702 VSS.n12728 VSS.n12727 292.5
R5703 VSS.n12783 VSS.n12782 292.5
R5704 VSS.n12784 VSS.n12783 292.5
R5705 VSS.n12729 VSS.n12726 292.5
R5706 VSS.n12785 VSS.n12726 292.5
R5707 VSS.n12787 VSS.n12724 292.5
R5708 VSS.n12787 VSS.n12786 292.5
R5709 VSS.n12059 VSS.n12058 292.5
R5710 VSS.n12221 VSS.n12059 292.5
R5711 VSS.n12063 VSS.n12061 292.5
R5712 VSS.n12061 VSS.n12060 292.5
R5713 VSS.n11988 VSS.n11986 292.5
R5714 VSS.n11993 VSS.n11988 292.5
R5715 VSS.n12299 VSS.n12298 292.5
R5716 VSS.n12300 VSS.n12299 292.5
R5717 VSS.n12002 VSS.n12001 292.5
R5718 VSS.n12289 VSS.n12002 292.5
R5719 VSS.n12010 VSS.n12008 292.5
R5720 VSS.n12012 VSS.n12010 292.5
R5721 VSS.n12276 VSS.n12275 292.5
R5722 VSS.n12277 VSS.n12276 292.5
R5723 VSS.n12021 VSS.n12020 292.5
R5724 VSS.n12266 VSS.n12021 292.5
R5725 VSS.n12029 VSS.n12027 292.5
R5726 VSS.n12031 VSS.n12029 292.5
R5727 VSS.n12254 VSS.n12253 292.5
R5728 VSS.n12255 VSS.n12254 292.5
R5729 VSS.n12040 VSS.n12039 292.5
R5730 VSS.n12244 VSS.n12040 292.5
R5731 VSS.n12048 VSS.n12046 292.5
R5732 VSS.n12050 VSS.n12048 292.5
R5733 VSS.n12231 VSS.n12230 292.5
R5734 VSS.n12232 VSS.n12231 292.5
R5735 VSS.n12065 VSS.n12064 292.5
R5736 VSS.n12209 VSS.n12065 292.5
R5737 VSS.n12207 VSS.n12206 292.5
R5738 VSS.n12208 VSS.n12207 292.5
R5739 VSS.n12205 VSS.n12067 292.5
R5740 VSS.n12067 VSS.n12066 292.5
R5741 VSS.n12204 VSS.n12203 292.5
R5742 VSS.n12203 VSS.n12202 292.5
R5743 VSS.n12069 VSS.n12068 292.5
R5744 VSS.n12201 VSS.n12069 292.5
R5745 VSS.n12199 VSS.n12198 292.5
R5746 VSS.n12200 VSS.n12199 292.5
R5747 VSS.n12197 VSS.n12071 292.5
R5748 VSS.n12071 VSS.n12070 292.5
R5749 VSS.n12196 VSS.n12195 292.5
R5750 VSS.n12195 VSS.n12194 292.5
R5751 VSS.n12073 VSS.n12072 292.5
R5752 VSS.n12193 VSS.n12073 292.5
R5753 VSS.n12191 VSS.n12190 292.5
R5754 VSS.n12192 VSS.n12191 292.5
R5755 VSS.n12189 VSS.n12075 292.5
R5756 VSS.n12075 VSS.n12074 292.5
R5757 VSS.n12212 VSS.n12211 292.5
R5758 VSS.n12211 VSS.n12210 292.5
R5759 VSS.n12165 VSS.n12087 292.5
R5760 VSS.n12087 VSS.n12086 292.5
R5761 VSS.n12167 VSS.n12166 292.5
R5762 VSS.n12168 VSS.n12167 292.5
R5763 VSS.n12085 VSS.n12084 292.5
R5764 VSS.n12169 VSS.n12085 292.5
R5765 VSS.n12172 VSS.n12171 292.5
R5766 VSS.n12171 VSS.n12170 292.5
R5767 VSS.n12173 VSS.n12083 292.5
R5768 VSS.n12083 VSS.n12082 292.5
R5769 VSS.n12175 VSS.n12174 292.5
R5770 VSS.n12176 VSS.n12175 292.5
R5771 VSS.n12081 VSS.n12080 292.5
R5772 VSS.n12177 VSS.n12081 292.5
R5773 VSS.n12180 VSS.n12179 292.5
R5774 VSS.n12179 VSS.n12178 292.5
R5775 VSS.n12181 VSS.n12079 292.5
R5776 VSS.n12079 VSS.n12078 292.5
R5777 VSS.n12183 VSS.n12182 292.5
R5778 VSS.n12184 VSS.n12183 292.5
R5779 VSS.n12077 VSS.n12076 292.5
R5780 VSS.n12185 VSS.n12077 292.5
R5781 VSS.n12188 VSS.n12187 292.5
R5782 VSS.n12187 VSS.n12186 292.5
R5783 VSS.n12136 VSS.n11528 292.5
R5784 VSS.n12136 VSS.n12135 292.5
R5785 VSS.n12138 VSS.n12137 292.5
R5786 VSS.n12137 VSS.n12134 292.5
R5787 VSS.n12140 VSS.n12139 292.5
R5788 VSS.n12141 VSS.n12140 292.5
R5789 VSS.n12133 VSS.n12132 292.5
R5790 VSS.n12142 VSS.n12133 292.5
R5791 VSS.n12145 VSS.n12144 292.5
R5792 VSS.n12144 VSS.n12143 292.5
R5793 VSS.n12146 VSS.n12131 292.5
R5794 VSS.n12131 VSS.n12130 292.5
R5795 VSS.n12148 VSS.n12147 292.5
R5796 VSS.n12149 VSS.n12148 292.5
R5797 VSS.n12129 VSS.n12128 292.5
R5798 VSS.n12150 VSS.n12129 292.5
R5799 VSS.n12154 VSS.n12153 292.5
R5800 VSS.n12153 VSS.n12152 292.5
R5801 VSS.n12155 VSS.n12127 292.5
R5802 VSS.n12151 VSS.n12127 292.5
R5803 VSS.n12157 VSS.n12156 292.5
R5804 VSS.n12157 VSS.n12126 292.5
R5805 VSS.n12158 VSS.n12088 292.5
R5806 VSS.n12159 VSS.n12158 292.5
R5807 VSS.n11980 VSS.n11979 292.5
R5808 VSS.n12313 VSS.n11980 292.5
R5809 VSS.n12323 VSS.n12322 292.5
R5810 VSS.n12324 VSS.n12323 292.5
R5811 VSS.n11969 VSS.n11967 292.5
R5812 VSS.n11971 VSS.n11969 292.5
R5813 VSS.n11961 VSS.n11960 292.5
R5814 VSS.n12336 VSS.n11961 292.5
R5815 VSS.n12346 VSS.n12345 292.5
R5816 VSS.n12347 VSS.n12346 292.5
R5817 VSS.n11950 VSS.n11948 292.5
R5818 VSS.n11952 VSS.n11950 292.5
R5819 VSS.n11942 VSS.n11941 292.5
R5820 VSS.n12358 VSS.n11942 292.5
R5821 VSS.n12368 VSS.n12367 292.5
R5822 VSS.n12369 VSS.n12368 292.5
R5823 VSS.n11931 VSS.n11929 292.5
R5824 VSS.n11933 VSS.n11931 292.5
R5825 VSS.n11923 VSS.n11922 292.5
R5826 VSS.n12381 VSS.n11923 292.5
R5827 VSS.n12391 VSS.n12390 292.5
R5828 VSS.n12392 VSS.n12391 292.5
R5829 VSS.n11912 VSS.n11908 292.5
R5830 VSS.n11914 VSS.n11912 292.5
R5831 VSS.n11546 VSS.n11545 292.5
R5832 VSS.n11545 VSS.n11544 292.5
R5833 VSS.n11899 VSS.n11898 292.5
R5834 VSS.n11900 VSS.n11899 292.5
R5835 VSS.n11557 VSS.n11555 292.5
R5836 VSS.n11889 VSS.n11557 292.5
R5837 VSS.n11880 VSS.n11879 292.5
R5838 VSS.n11879 VSS.n11878 292.5
R5839 VSS.n11566 VSS.n11565 292.5
R5840 VSS.n11565 VSS.n11564 292.5
R5841 VSS.n11864 VSS.n11863 292.5
R5842 VSS.n11865 VSS.n11864 292.5
R5843 VSS.n11578 VSS.n11576 292.5
R5844 VSS.n11855 VSS.n11578 292.5
R5845 VSS.n11846 VSS.n11845 292.5
R5846 VSS.n11845 VSS.n11844 292.5
R5847 VSS.n11587 VSS.n11586 292.5
R5848 VSS.n11586 VSS.n11585 292.5
R5849 VSS.n11830 VSS.n11829 292.5
R5850 VSS.n11831 VSS.n11830 292.5
R5851 VSS.n11599 VSS.n11597 292.5
R5852 VSS.n11820 VSS.n11599 292.5
R5853 VSS.n11811 VSS.n11810 292.5
R5854 VSS.n11810 VSS.n11809 292.5
R5855 VSS.n12458 VSS.n12457 292.5
R5856 VSS.n12457 VSS.n11510 292.5
R5857 VSS.n12456 VSS.n11515 292.5
R5858 VSS.n12456 VSS.n12455 292.5
R5859 VSS.n11519 VSS.n11516 292.5
R5860 VSS.n12454 VSS.n11516 292.5
R5861 VSS.n12452 VSS.n12451 292.5
R5862 VSS.n12453 VSS.n12452 292.5
R5863 VSS.n12450 VSS.n11518 292.5
R5864 VSS.n11518 VSS.n11517 292.5
R5865 VSS.n12449 VSS.n12448 292.5
R5866 VSS.n12448 VSS.n12447 292.5
R5867 VSS.n11521 VSS.n11520 292.5
R5868 VSS.n12446 VSS.n11521 292.5
R5869 VSS.n12444 VSS.n12443 292.5
R5870 VSS.n12445 VSS.n12444 292.5
R5871 VSS.n12442 VSS.n11523 292.5
R5872 VSS.n11523 VSS.n11522 292.5
R5873 VSS.n12441 VSS.n12440 292.5
R5874 VSS.n12440 VSS.n12439 292.5
R5875 VSS.n11525 VSS.n11524 292.5
R5876 VSS.n12438 VSS.n11525 292.5
R5877 VSS.n12436 VSS.n12435 292.5
R5878 VSS.n12437 VSS.n12436 292.5
R5879 VSS.n12486 VSS.n12485 292.5
R5880 VSS.n12487 VSS.n12486 292.5
R5881 VSS.n12484 VSS.n11499 292.5
R5882 VSS.n11499 VSS.n11498 292.5
R5883 VSS.n12483 VSS.n12482 292.5
R5884 VSS.n12482 VSS.n12481 292.5
R5885 VSS.n11501 VSS.n11500 292.5
R5886 VSS.n12480 VSS.n11501 292.5
R5887 VSS.n12478 VSS.n12477 292.5
R5888 VSS.n12479 VSS.n12478 292.5
R5889 VSS.n12476 VSS.n11503 292.5
R5890 VSS.n11503 VSS.n11502 292.5
R5891 VSS.n12475 VSS.n12474 292.5
R5892 VSS.n12474 VSS.n12473 292.5
R5893 VSS.n11505 VSS.n11504 292.5
R5894 VSS.n12472 VSS.n11505 292.5
R5895 VSS.n12470 VSS.n12469 292.5
R5896 VSS.n12471 VSS.n12470 292.5
R5897 VSS.n12468 VSS.n11507 292.5
R5898 VSS.n11507 VSS.n11506 292.5
R5899 VSS.n12467 VSS.n12466 292.5
R5900 VSS.n12466 VSS.n12465 292.5
R5901 VSS.n11509 VSS.n11508 292.5
R5902 VSS.n12464 VSS.n11509 292.5
R5903 VSS.n11768 VSS.n11612 292.5
R5904 VSS.n11768 VSS.n11767 292.5
R5905 VSS.n11616 VSS.n11615 292.5
R5906 VSS.n11615 VSS.n11614 292.5
R5907 VSS.n11753 VSS.n11752 292.5
R5908 VSS.n11754 VSS.n11753 292.5
R5909 VSS.n11629 VSS.n11627 292.5
R5910 VSS.n11743 VSS.n11629 292.5
R5911 VSS.n11734 VSS.n11733 292.5
R5912 VSS.n11733 VSS.n11732 292.5
R5913 VSS.n11638 VSS.n11637 292.5
R5914 VSS.n11637 VSS.n11636 292.5
R5915 VSS.n11719 VSS.n11718 292.5
R5916 VSS.n11720 VSS.n11719 292.5
R5917 VSS.n11650 VSS.n11648 292.5
R5918 VSS.n11709 VSS.n11650 292.5
R5919 VSS.n11700 VSS.n11699 292.5
R5920 VSS.n11699 VSS.n11698 292.5
R5921 VSS.n11659 VSS.n11658 292.5
R5922 VSS.n11658 VSS.n11657 292.5
R5923 VSS.n11684 VSS.n11683 292.5
R5924 VSS.n11685 VSS.n11684 292.5
R5925 VSS.n11671 VSS.n11669 292.5
R5926 VSS.n11674 VSS.n11671 292.5
R5927 VSS.n13405 VSS.n13404 292.5
R5928 VSS.n13406 VSS.n13405 292.5
R5929 VSS.n11471 VSS.n11469 292.5
R5930 VSS.n11473 VSS.n11471 292.5
R5931 VSS.n11463 VSS.n11462 292.5
R5932 VSS.n13418 VSS.n11463 292.5
R5933 VSS.n13428 VSS.n13427 292.5
R5934 VSS.n13429 VSS.n13428 292.5
R5935 VSS.n11452 VSS.n11450 292.5
R5936 VSS.n11454 VSS.n11452 292.5
R5937 VSS.n11444 VSS.n11443 292.5
R5938 VSS.n13440 VSS.n11444 292.5
R5939 VSS.n13450 VSS.n13449 292.5
R5940 VSS.n13451 VSS.n13450 292.5
R5941 VSS.n11433 VSS.n11431 292.5
R5942 VSS.n11435 VSS.n11433 292.5
R5943 VSS.n13280 VSS.n13279 292.5
R5944 VSS.n13281 VSS.n13280 292.5
R5945 VSS.n13263 VSS.n13261 292.5
R5946 VSS.n13265 VSS.n13263 292.5
R5947 VSS.n13254 VSS.n13253 292.5
R5948 VSS.n13293 VSS.n13254 292.5
R5949 VSS.n13303 VSS.n13302 292.5
R5950 VSS.n13303 VSS.n13249 292.5
R5951 VSS.n12499 VSS.n12498 292.5
R5952 VSS.n13346 VSS.n12499 292.5
R5953 VSS.n13349 VSS.n13348 292.5
R5954 VSS.n13348 VSS.n13347 292.5
R5955 VSS.n13350 VSS.n12497 292.5
R5956 VSS.n12497 VSS.n12496 292.5
R5957 VSS.n13352 VSS.n13351 292.5
R5958 VSS.n13353 VSS.n13352 292.5
R5959 VSS.n12495 VSS.n12494 292.5
R5960 VSS.n13354 VSS.n12495 292.5
R5961 VSS.n13357 VSS.n13356 292.5
R5962 VSS.n13356 VSS.n13355 292.5
R5963 VSS.n13358 VSS.n12493 292.5
R5964 VSS.n12493 VSS.n12492 292.5
R5965 VSS.n13360 VSS.n13359 292.5
R5966 VSS.n13361 VSS.n13360 292.5
R5967 VSS.n12491 VSS.n12490 292.5
R5968 VSS.n13362 VSS.n12491 292.5
R5969 VSS.n13365 VSS.n13364 292.5
R5970 VSS.n13364 VSS.n13363 292.5
R5971 VSS.n13366 VSS.n12489 292.5
R5972 VSS.n12489 VSS.n12488 292.5
R5973 VSS.n13368 VSS.n13367 292.5
R5974 VSS.n13369 VSS.n13368 292.5
R5975 VSS.n12627 VSS.n12626 292.5
R5976 VSS.n12628 VSS.n12627 292.5
R5977 VSS.n12625 VSS.n12600 292.5
R5978 VSS.n12600 VSS.n12599 292.5
R5979 VSS.n12624 VSS.n12623 292.5
R5980 VSS.n12623 VSS.n12622 292.5
R5981 VSS.n12602 VSS.n12601 292.5
R5982 VSS.n12621 VSS.n12602 292.5
R5983 VSS.n12619 VSS.n12618 292.5
R5984 VSS.n12620 VSS.n12619 292.5
R5985 VSS.n12617 VSS.n12604 292.5
R5986 VSS.n12604 VSS.n12603 292.5
R5987 VSS.n12616 VSS.n12615 292.5
R5988 VSS.n12615 VSS.n12614 292.5
R5989 VSS.n12606 VSS.n12605 292.5
R5990 VSS.n12613 VSS.n12606 292.5
R5991 VSS.n12611 VSS.n12610 292.5
R5992 VSS.n12612 VSS.n12611 292.5
R5993 VSS.n12609 VSS.n12608 292.5
R5994 VSS.n12608 VSS.n12607 292.5
R5995 VSS.n12504 VSS.n12502 292.5
R5996 VSS.n12502 VSS.n12501 292.5
R5997 VSS.n13343 VSS.n13342 292.5
R5998 VSS.n13344 VSS.n13343 292.5
R5999 VSS.n12522 VSS.n12521 292.5
R6000 VSS.n13248 VSS.n12522 292.5
R6001 VSS.n12531 VSS.n12529 292.5
R6002 VSS.n13235 VSS.n12531 292.5
R6003 VSS.n13232 VSS.n13231 292.5
R6004 VSS.n13233 VSS.n13232 292.5
R6005 VSS.n12538 VSS.n12536 292.5
R6006 VSS.n13222 VSS.n12538 292.5
R6007 VSS.n13213 VSS.n13212 292.5
R6008 VSS.n13212 VSS.n13211 292.5
R6009 VSS.n12547 VSS.n12546 292.5
R6010 VSS.n12546 VSS.n12545 292.5
R6011 VSS.n13198 VSS.n13197 292.5
R6012 VSS.n13199 VSS.n13198 292.5
R6013 VSS.n12559 VSS.n12557 292.5
R6014 VSS.n13188 VSS.n12559 292.5
R6015 VSS.n13179 VSS.n13178 292.5
R6016 VSS.n13178 VSS.n13177 292.5
R6017 VSS.n12568 VSS.n12567 292.5
R6018 VSS.n12567 VSS.n12566 292.5
R6019 VSS.n13163 VSS.n13162 292.5
R6020 VSS.n13164 VSS.n13163 292.5
R6021 VSS.n12580 VSS.n12578 292.5
R6022 VSS.n13153 VSS.n12580 292.5
R6023 VSS.n12964 VSS.n12962 292.5
R6024 VSS.n12965 VSS.n12964 292.5
R6025 VSS.n12955 VSS.n12954 292.5
R6026 VSS.n12976 VSS.n12955 292.5
R6027 VSS.n12986 VSS.n12985 292.5
R6028 VSS.n12987 VSS.n12986 292.5
R6029 VSS.n12944 VSS.n12942 292.5
R6030 VSS.n12946 VSS.n12944 292.5
R6031 VSS.n12936 VSS.n12935 292.5
R6032 VSS.n12999 VSS.n12936 292.5
R6033 VSS.n13008 VSS.n13007 292.5
R6034 VSS.n13009 VSS.n13008 292.5
R6035 VSS.n12925 VSS.n12923 292.5
R6036 VSS.n12927 VSS.n12925 292.5
R6037 VSS.n12917 VSS.n12916 292.5
R6038 VSS.n13021 VSS.n12917 292.5
R6039 VSS.n13031 VSS.n13030 292.5
R6040 VSS.n13032 VSS.n13031 292.5
R6041 VSS.n12906 VSS.n12904 292.5
R6042 VSS.n12908 VSS.n12906 292.5
R6043 VSS.n12897 VSS.n12896 292.5
R6044 VSS.n13044 VSS.n12897 292.5
R6045 VSS.n13054 VSS.n13053 292.5
R6046 VSS.n13054 VSS.n12892 292.5
R6047 VSS.n12640 VSS.n12639 292.5
R6048 VSS.n13097 VSS.n12640 292.5
R6049 VSS.n13100 VSS.n13099 292.5
R6050 VSS.n13099 VSS.n13098 292.5
R6051 VSS.n13101 VSS.n12638 292.5
R6052 VSS.n12638 VSS.n12637 292.5
R6053 VSS.n13103 VSS.n13102 292.5
R6054 VSS.n13104 VSS.n13103 292.5
R6055 VSS.n12636 VSS.n12635 292.5
R6056 VSS.n13105 VSS.n12636 292.5
R6057 VSS.n13108 VSS.n13107 292.5
R6058 VSS.n13107 VSS.n13106 292.5
R6059 VSS.n13109 VSS.n12634 292.5
R6060 VSS.n12634 VSS.n12633 292.5
R6061 VSS.n13111 VSS.n13110 292.5
R6062 VSS.n13112 VSS.n13111 292.5
R6063 VSS.n12632 VSS.n12631 292.5
R6064 VSS.n13113 VSS.n12632 292.5
R6065 VSS.n13116 VSS.n13115 292.5
R6066 VSS.n13115 VSS.n13114 292.5
R6067 VSS.n13117 VSS.n12630 292.5
R6068 VSS.n12630 VSS.n12629 292.5
R6069 VSS.n13119 VSS.n13118 292.5
R6070 VSS.n13120 VSS.n13119 292.5
R6071 VSS.n12764 VSS.n12763 292.5
R6072 VSS.n12763 VSS.n12762 292.5
R6073 VSS.n12739 VSS.n12738 292.5
R6074 VSS.n12761 VSS.n12739 292.5
R6075 VSS.n12759 VSS.n12758 292.5
R6076 VSS.n12760 VSS.n12759 292.5
R6077 VSS.n12757 VSS.n12741 292.5
R6078 VSS.n12741 VSS.n12740 292.5
R6079 VSS.n12756 VSS.n12755 292.5
R6080 VSS.n12755 VSS.n12754 292.5
R6081 VSS.n12743 VSS.n12742 292.5
R6082 VSS.n12753 VSS.n12743 292.5
R6083 VSS.n12751 VSS.n12750 292.5
R6084 VSS.n12752 VSS.n12751 292.5
R6085 VSS.n12749 VSS.n12745 292.5
R6086 VSS.n12745 VSS.n12744 292.5
R6087 VSS.n12748 VSS.n12747 292.5
R6088 VSS.n12747 VSS.n12746 292.5
R6089 VSS.n12645 VSS.n12643 292.5
R6090 VSS.n12643 VSS.n12642 292.5
R6091 VSS.n13094 VSS.n13093 292.5
R6092 VSS.n13095 VSS.n13094 292.5
R6093 VSS.n12765 VSS.n12737 292.5
R6094 VSS.n12737 VSS.n12736 292.5
R6095 VSS.n12663 VSS.n12662 292.5
R6096 VSS.n12891 VSS.n12663 292.5
R6097 VSS.n12672 VSS.n12670 292.5
R6098 VSS.n12878 VSS.n12672 292.5
R6099 VSS.n12875 VSS.n12874 292.5
R6100 VSS.n12876 VSS.n12875 292.5
R6101 VSS.n12679 VSS.n12677 292.5
R6102 VSS.n12865 VSS.n12679 292.5
R6103 VSS.n12856 VSS.n12855 292.5
R6104 VSS.n12855 VSS.n12854 292.5
R6105 VSS.n12688 VSS.n12687 292.5
R6106 VSS.n12687 VSS.n12686 292.5
R6107 VSS.n12841 VSS.n12840 292.5
R6108 VSS.n12842 VSS.n12841 292.5
R6109 VSS.n12700 VSS.n12698 292.5
R6110 VSS.n12831 VSS.n12700 292.5
R6111 VSS.n12822 VSS.n12821 292.5
R6112 VSS.n12821 VSS.n12820 292.5
R6113 VSS.n12709 VSS.n12708 292.5
R6114 VSS.n12708 VSS.n12707 292.5
R6115 VSS.n12806 VSS.n12805 292.5
R6116 VSS.n12807 VSS.n12806 292.5
R6117 VSS.n12721 VSS.n12719 292.5
R6118 VSS.n12796 VSS.n12721 292.5
R6119 VSS.n12791 VSS.n12790 292.5
R6120 VSS.n7842 VSS.n7670 292.5
R6121 VSS.n7670 VSS.n7669 292.5
R6122 VSS.n7865 VSS.n7864 292.5
R6123 VSS.n7864 VSS.n7863 292.5
R6124 VSS.n7660 VSS.n7659 292.5
R6125 VSS.n7862 VSS.n7660 292.5
R6126 VSS.n7860 VSS.n7859 292.5
R6127 VSS.n7861 VSS.n7860 292.5
R6128 VSS.n7858 VSS.n7662 292.5
R6129 VSS.n7662 VSS.n7661 292.5
R6130 VSS.n7857 VSS.n7856 292.5
R6131 VSS.n7856 VSS.n7855 292.5
R6132 VSS.n7664 VSS.n7663 292.5
R6133 VSS.n7854 VSS.n7664 292.5
R6134 VSS.n7852 VSS.n7851 292.5
R6135 VSS.n7853 VSS.n7852 292.5
R6136 VSS.n7850 VSS.n7666 292.5
R6137 VSS.n7666 VSS.n7665 292.5
R6138 VSS.n7849 VSS.n7848 292.5
R6139 VSS.n7848 VSS.n7847 292.5
R6140 VSS.n7668 VSS.n7667 292.5
R6141 VSS.n7846 VSS.n7668 292.5
R6142 VSS.n7844 VSS.n7843 292.5
R6143 VSS.n7845 VSS.n7844 292.5
R6144 VSS.n7009 VSS.n7007 292.5
R6145 VSS.n7169 VSS.n7009 292.5
R6146 VSS.n7010 VSS.n7005 292.5
R6147 VSS.n7170 VSS.n7010 292.5
R6148 VSS.n7075 VSS.n7074 292.5
R6149 VSS.n7076 VSS.n7075 292.5
R6150 VSS.n7061 VSS.n7060 292.5
R6151 VSS.n7060 VSS.n7059 292.5
R6152 VSS.n7091 VSS.n7090 292.5
R6153 VSS.n7090 VSS.n7089 292.5
R6154 VSS.n7052 VSS.n7050 292.5
R6155 VSS.n7100 VSS.n7052 292.5
R6156 VSS.n7110 VSS.n7109 292.5
R6157 VSS.n7111 VSS.n7110 292.5
R6158 VSS.n7040 VSS.n7039 292.5
R6159 VSS.n7039 VSS.n7038 292.5
R6160 VSS.n7126 VSS.n7125 292.5
R6161 VSS.n7125 VSS.n7124 292.5
R6162 VSS.n7031 VSS.n7029 292.5
R6163 VSS.n7134 VSS.n7031 292.5
R6164 VSS.n7144 VSS.n7143 292.5
R6165 VSS.n7145 VSS.n7144 292.5
R6166 VSS.n7019 VSS.n7018 292.5
R6167 VSS.n7018 VSS.n7017 292.5
R6168 VSS.n7160 VSS.n7159 292.5
R6169 VSS.n7159 VSS.n7158 292.5
R6170 VSS.n7181 VSS.n7180 292.5
R6171 VSS.n7182 VSS.n7181 292.5
R6172 VSS.n7002 VSS.n7001 292.5
R6173 VSS.n7183 VSS.n7002 292.5
R6174 VSS.n7186 VSS.n7185 292.5
R6175 VSS.n7185 VSS.n7184 292.5
R6176 VSS.n7187 VSS.n7000 292.5
R6177 VSS.n7000 VSS.n6999 292.5
R6178 VSS.n7189 VSS.n7188 292.5
R6179 VSS.n7190 VSS.n7189 292.5
R6180 VSS.n6998 VSS.n6997 292.5
R6181 VSS.n7191 VSS.n6998 292.5
R6182 VSS.n7194 VSS.n7193 292.5
R6183 VSS.n7193 VSS.n7192 292.5
R6184 VSS.n7195 VSS.n6996 292.5
R6185 VSS.n6996 VSS.n6995 292.5
R6186 VSS.n7197 VSS.n7196 292.5
R6187 VSS.n7198 VSS.n7197 292.5
R6188 VSS.n6994 VSS.n6993 292.5
R6189 VSS.n7199 VSS.n6994 292.5
R6190 VSS.n7202 VSS.n7201 292.5
R6191 VSS.n7201 VSS.n7200 292.5
R6192 VSS.n7179 VSS.n7004 292.5
R6193 VSS.n7004 VSS.n7003 292.5
R6194 VSS.n7226 VSS.n7225 292.5
R6195 VSS.n7225 VSS.n7224 292.5
R6196 VSS.n6982 VSS.n6981 292.5
R6197 VSS.n7223 VSS.n6982 292.5
R6198 VSS.n7221 VSS.n7220 292.5
R6199 VSS.n7222 VSS.n7221 292.5
R6200 VSS.n7219 VSS.n6984 292.5
R6201 VSS.n6984 VSS.n6983 292.5
R6202 VSS.n7218 VSS.n7217 292.5
R6203 VSS.n7217 VSS.n7216 292.5
R6204 VSS.n6986 VSS.n6985 292.5
R6205 VSS.n7215 VSS.n6986 292.5
R6206 VSS.n7213 VSS.n7212 292.5
R6207 VSS.n7214 VSS.n7213 292.5
R6208 VSS.n7211 VSS.n6988 292.5
R6209 VSS.n6988 VSS.n6987 292.5
R6210 VSS.n7210 VSS.n7209 292.5
R6211 VSS.n7209 VSS.n7208 292.5
R6212 VSS.n6990 VSS.n6989 292.5
R6213 VSS.n7207 VSS.n6990 292.5
R6214 VSS.n7205 VSS.n7204 292.5
R6215 VSS.n7206 VSS.n7205 292.5
R6216 VSS.n7203 VSS.n6992 292.5
R6217 VSS.n6992 VSS.n6991 292.5
R6218 VSS.n8804 VSS.n7238 292.5
R6219 VSS.n7238 VSS.n7237 292.5
R6220 VSS.n8806 VSS.n8805 292.5
R6221 VSS.n8807 VSS.n8806 292.5
R6222 VSS.n7236 VSS.n7235 292.5
R6223 VSS.n8808 VSS.n7236 292.5
R6224 VSS.n8811 VSS.n8810 292.5
R6225 VSS.n8810 VSS.n8809 292.5
R6226 VSS.n8812 VSS.n7234 292.5
R6227 VSS.n7234 VSS.n7233 292.5
R6228 VSS.n8814 VSS.n8813 292.5
R6229 VSS.n8815 VSS.n8814 292.5
R6230 VSS.n7232 VSS.n7231 292.5
R6231 VSS.n8816 VSS.n7232 292.5
R6232 VSS.n8819 VSS.n8818 292.5
R6233 VSS.n8818 VSS.n8817 292.5
R6234 VSS.n8820 VSS.n7230 292.5
R6235 VSS.n7230 VSS.n7229 292.5
R6236 VSS.n8822 VSS.n8821 292.5
R6237 VSS.n8823 VSS.n8822 292.5
R6238 VSS.n7228 VSS.n7227 292.5
R6239 VSS.n8824 VSS.n7228 292.5
R6240 VSS.n8827 VSS.n8826 292.5
R6241 VSS.n8826 VSS.n8825 292.5
R6242 VSS.n6962 VSS.n6960 292.5
R6243 VSS.n6964 VSS.n6962 292.5
R6244 VSS.n6954 VSS.n6953 292.5
R6245 VSS.n8867 VSS.n6954 292.5
R6246 VSS.n8877 VSS.n8876 292.5
R6247 VSS.n8878 VSS.n8877 292.5
R6248 VSS.n6943 VSS.n6941 292.5
R6249 VSS.n6945 VSS.n6943 292.5
R6250 VSS.n6935 VSS.n6934 292.5
R6251 VSS.n8890 VSS.n6935 292.5
R6252 VSS.n8899 VSS.n8898 292.5
R6253 VSS.n8900 VSS.n8899 292.5
R6254 VSS.n6924 VSS.n6922 292.5
R6255 VSS.n6926 VSS.n6924 292.5
R6256 VSS.n6916 VSS.n6915 292.5
R6257 VSS.n8912 VSS.n6916 292.5
R6258 VSS.n8922 VSS.n8921 292.5
R6259 VSS.n8923 VSS.n8922 292.5
R6260 VSS.n6905 VSS.n6903 292.5
R6261 VSS.n6907 VSS.n6905 292.5
R6262 VSS.n8755 VSS.n8738 292.5
R6263 VSS.n8738 VSS.n8737 292.5
R6264 VSS.n8761 VSS.n8735 292.5
R6265 VSS.n8761 VSS.n8760 292.5
R6266 VSS.n7260 VSS.n7258 292.5
R6267 VSS.n7258 VSS.n7257 292.5
R6268 VSS.n8726 VSS.n8725 292.5
R6269 VSS.n8727 VSS.n8726 292.5
R6270 VSS.n7271 VSS.n7269 292.5
R6271 VSS.n8716 VSS.n7271 292.5
R6272 VSS.n8707 VSS.n8706 292.5
R6273 VSS.n8706 VSS.n8705 292.5
R6274 VSS.n7280 VSS.n7279 292.5
R6275 VSS.n7279 VSS.n7278 292.5
R6276 VSS.n8691 VSS.n8690 292.5
R6277 VSS.n8692 VSS.n8691 292.5
R6278 VSS.n7292 VSS.n7290 292.5
R6279 VSS.n8682 VSS.n7292 292.5
R6280 VSS.n8673 VSS.n8672 292.5
R6281 VSS.n8672 VSS.n8671 292.5
R6282 VSS.n7301 VSS.n7300 292.5
R6283 VSS.n7300 VSS.n7299 292.5
R6284 VSS.n8657 VSS.n8656 292.5
R6285 VSS.n8658 VSS.n8657 292.5
R6286 VSS.n7313 VSS.n7311 292.5
R6287 VSS.n8647 VSS.n7313 292.5
R6288 VSS.n8638 VSS.n8637 292.5
R6289 VSS.n8637 VSS.n8636 292.5
R6290 VSS.n7366 VSS.n7365 292.5
R6291 VSS.n7365 VSS.n7364 292.5
R6292 VSS.n7338 VSS.n7337 292.5
R6293 VSS.n7363 VSS.n7338 292.5
R6294 VSS.n7361 VSS.n7360 292.5
R6295 VSS.n7362 VSS.n7361 292.5
R6296 VSS.n7359 VSS.n7340 292.5
R6297 VSS.n7340 VSS.n7339 292.5
R6298 VSS.n7358 VSS.n7357 292.5
R6299 VSS.n7357 VSS.n7356 292.5
R6300 VSS.n7342 VSS.n7341 292.5
R6301 VSS.n7355 VSS.n7342 292.5
R6302 VSS.n7353 VSS.n7352 292.5
R6303 VSS.n7354 VSS.n7353 292.5
R6304 VSS.n7351 VSS.n7344 292.5
R6305 VSS.n7344 VSS.n7343 292.5
R6306 VSS.n7350 VSS.n7349 292.5
R6307 VSS.n7349 VSS.n7348 292.5
R6308 VSS.n7346 VSS.n7345 292.5
R6309 VSS.n7347 VSS.n7346 292.5
R6310 VSS.n7241 VSS.n7240 292.5
R6311 VSS.n7243 VSS.n7241 292.5
R6312 VSS.n8802 VSS.n8801 292.5
R6313 VSS.n8801 VSS.n8800 292.5
R6314 VSS.n8582 VSS.n7378 292.5
R6315 VSS.n7378 VSS.n7377 292.5
R6316 VSS.n8584 VSS.n8583 292.5
R6317 VSS.n8585 VSS.n8584 292.5
R6318 VSS.n7376 VSS.n7375 292.5
R6319 VSS.n8586 VSS.n7376 292.5
R6320 VSS.n8589 VSS.n8588 292.5
R6321 VSS.n8588 VSS.n8587 292.5
R6322 VSS.n8590 VSS.n7374 292.5
R6323 VSS.n7374 VSS.n7373 292.5
R6324 VSS.n8592 VSS.n8591 292.5
R6325 VSS.n8593 VSS.n8592 292.5
R6326 VSS.n7372 VSS.n7371 292.5
R6327 VSS.n8594 VSS.n7372 292.5
R6328 VSS.n8597 VSS.n8596 292.5
R6329 VSS.n8596 VSS.n8595 292.5
R6330 VSS.n8598 VSS.n7370 292.5
R6331 VSS.n7370 VSS.n7369 292.5
R6332 VSS.n8600 VSS.n8599 292.5
R6333 VSS.n8601 VSS.n8600 292.5
R6334 VSS.n7368 VSS.n7367 292.5
R6335 VSS.n8602 VSS.n7368 292.5
R6336 VSS.n8605 VSS.n8604 292.5
R6337 VSS.n8604 VSS.n8603 292.5
R6338 VSS.n8459 VSS.n8458 292.5
R6339 VSS.n8460 VSS.n8459 292.5
R6340 VSS.n8445 VSS.n8443 292.5
R6341 VSS.n8447 VSS.n8445 292.5
R6342 VSS.n8437 VSS.n8436 292.5
R6343 VSS.n8472 VSS.n8437 292.5
R6344 VSS.n8482 VSS.n8481 292.5
R6345 VSS.n8483 VSS.n8482 292.5
R6346 VSS.n8426 VSS.n8424 292.5
R6347 VSS.n8428 VSS.n8426 292.5
R6348 VSS.n8418 VSS.n8417 292.5
R6349 VSS.n8494 VSS.n8418 292.5
R6350 VSS.n8504 VSS.n8503 292.5
R6351 VSS.n8505 VSS.n8504 292.5
R6352 VSS.n8407 VSS.n8405 292.5
R6353 VSS.n8409 VSS.n8407 292.5
R6354 VSS.n8399 VSS.n8398 292.5
R6355 VSS.n8517 VSS.n8399 292.5
R6356 VSS.n8527 VSS.n8526 292.5
R6357 VSS.n8528 VSS.n8527 292.5
R6358 VSS.n8533 VSS.n8380 292.5
R6359 VSS.n8380 VSS.n8379 292.5
R6360 VSS.n8539 VSS.n8377 292.5
R6361 VSS.n8539 VSS.n8538 292.5
R6362 VSS.n7400 VSS.n7398 292.5
R6363 VSS.n7398 VSS.n7397 292.5
R6364 VSS.n8368 VSS.n8367 292.5
R6365 VSS.n8369 VSS.n8368 292.5
R6366 VSS.n7411 VSS.n7409 292.5
R6367 VSS.n8358 VSS.n7411 292.5
R6368 VSS.n8349 VSS.n8348 292.5
R6369 VSS.n8348 VSS.n8347 292.5
R6370 VSS.n7420 VSS.n7419 292.5
R6371 VSS.n7419 VSS.n7418 292.5
R6372 VSS.n8333 VSS.n8332 292.5
R6373 VSS.n8334 VSS.n8333 292.5
R6374 VSS.n7432 VSS.n7430 292.5
R6375 VSS.n8324 VSS.n7432 292.5
R6376 VSS.n8315 VSS.n8314 292.5
R6377 VSS.n8314 VSS.n8313 292.5
R6378 VSS.n7441 VSS.n7440 292.5
R6379 VSS.n7440 VSS.n7439 292.5
R6380 VSS.n8299 VSS.n8298 292.5
R6381 VSS.n8300 VSS.n8299 292.5
R6382 VSS.n7453 VSS.n7451 292.5
R6383 VSS.n8289 VSS.n7453 292.5
R6384 VSS.n8280 VSS.n8279 292.5
R6385 VSS.n8279 VSS.n8278 292.5
R6386 VSS.n7506 VSS.n7505 292.5
R6387 VSS.n7505 VSS.n7504 292.5
R6388 VSS.n7478 VSS.n7477 292.5
R6389 VSS.n7503 VSS.n7478 292.5
R6390 VSS.n7501 VSS.n7500 292.5
R6391 VSS.n7502 VSS.n7501 292.5
R6392 VSS.n7499 VSS.n7480 292.5
R6393 VSS.n7480 VSS.n7479 292.5
R6394 VSS.n7498 VSS.n7497 292.5
R6395 VSS.n7497 VSS.n7496 292.5
R6396 VSS.n7482 VSS.n7481 292.5
R6397 VSS.n7495 VSS.n7482 292.5
R6398 VSS.n7493 VSS.n7492 292.5
R6399 VSS.n7494 VSS.n7493 292.5
R6400 VSS.n7491 VSS.n7484 292.5
R6401 VSS.n7484 VSS.n7483 292.5
R6402 VSS.n7490 VSS.n7489 292.5
R6403 VSS.n7489 VSS.n7488 292.5
R6404 VSS.n7486 VSS.n7485 292.5
R6405 VSS.n7487 VSS.n7486 292.5
R6406 VSS.n7381 VSS.n7380 292.5
R6407 VSS.n7383 VSS.n7381 292.5
R6408 VSS.n8580 VSS.n8579 292.5
R6409 VSS.n8579 VSS.n8578 292.5
R6410 VSS.n8224 VSS.n7518 292.5
R6411 VSS.n7518 VSS.n7517 292.5
R6412 VSS.n8226 VSS.n8225 292.5
R6413 VSS.n8227 VSS.n8226 292.5
R6414 VSS.n7516 VSS.n7515 292.5
R6415 VSS.n8228 VSS.n7516 292.5
R6416 VSS.n8231 VSS.n8230 292.5
R6417 VSS.n8230 VSS.n8229 292.5
R6418 VSS.n8232 VSS.n7514 292.5
R6419 VSS.n7514 VSS.n7513 292.5
R6420 VSS.n8234 VSS.n8233 292.5
R6421 VSS.n8235 VSS.n8234 292.5
R6422 VSS.n7512 VSS.n7511 292.5
R6423 VSS.n8236 VSS.n7512 292.5
R6424 VSS.n8239 VSS.n8238 292.5
R6425 VSS.n8238 VSS.n8237 292.5
R6426 VSS.n8240 VSS.n7510 292.5
R6427 VSS.n7510 VSS.n7509 292.5
R6428 VSS.n8242 VSS.n8241 292.5
R6429 VSS.n8243 VSS.n8242 292.5
R6430 VSS.n7508 VSS.n7507 292.5
R6431 VSS.n8244 VSS.n7508 292.5
R6432 VSS.n8247 VSS.n8246 292.5
R6433 VSS.n8246 VSS.n8245 292.5
R6434 VSS.n8101 VSS.n8100 292.5
R6435 VSS.n8102 VSS.n8101 292.5
R6436 VSS.n8087 VSS.n8085 292.5
R6437 VSS.n8089 VSS.n8087 292.5
R6438 VSS.n8079 VSS.n8078 292.5
R6439 VSS.n8114 VSS.n8079 292.5
R6440 VSS.n8124 VSS.n8123 292.5
R6441 VSS.n8125 VSS.n8124 292.5
R6442 VSS.n8068 VSS.n8066 292.5
R6443 VSS.n8070 VSS.n8068 292.5
R6444 VSS.n8060 VSS.n8059 292.5
R6445 VSS.n8136 VSS.n8060 292.5
R6446 VSS.n8146 VSS.n8145 292.5
R6447 VSS.n8147 VSS.n8146 292.5
R6448 VSS.n8049 VSS.n8047 292.5
R6449 VSS.n8051 VSS.n8049 292.5
R6450 VSS.n8041 VSS.n8040 292.5
R6451 VSS.n8159 VSS.n8041 292.5
R6452 VSS.n8169 VSS.n8168 292.5
R6453 VSS.n8170 VSS.n8169 292.5
R6454 VSS.n8175 VSS.n8022 292.5
R6455 VSS.n8022 VSS.n8021 292.5
R6456 VSS.n8181 VSS.n8019 292.5
R6457 VSS.n8181 VSS.n8180 292.5
R6458 VSS.n7540 VSS.n7538 292.5
R6459 VSS.n7538 VSS.n7537 292.5
R6460 VSS.n8010 VSS.n8009 292.5
R6461 VSS.n8011 VSS.n8010 292.5
R6462 VSS.n7551 VSS.n7549 292.5
R6463 VSS.n8000 VSS.n7551 292.5
R6464 VSS.n7991 VSS.n7990 292.5
R6465 VSS.n7990 VSS.n7989 292.5
R6466 VSS.n7560 VSS.n7559 292.5
R6467 VSS.n7559 VSS.n7558 292.5
R6468 VSS.n7975 VSS.n7974 292.5
R6469 VSS.n7976 VSS.n7975 292.5
R6470 VSS.n7572 VSS.n7570 292.5
R6471 VSS.n7966 VSS.n7572 292.5
R6472 VSS.n7957 VSS.n7956 292.5
R6473 VSS.n7956 VSS.n7955 292.5
R6474 VSS.n7581 VSS.n7580 292.5
R6475 VSS.n7580 VSS.n7579 292.5
R6476 VSS.n7941 VSS.n7940 292.5
R6477 VSS.n7942 VSS.n7941 292.5
R6478 VSS.n7593 VSS.n7591 292.5
R6479 VSS.n7931 VSS.n7593 292.5
R6480 VSS.n7922 VSS.n7921 292.5
R6481 VSS.n7921 VSS.n7920 292.5
R6482 VSS.n7646 VSS.n7645 292.5
R6483 VSS.n7645 VSS.n7644 292.5
R6484 VSS.n7618 VSS.n7617 292.5
R6485 VSS.n7643 VSS.n7618 292.5
R6486 VSS.n7641 VSS.n7640 292.5
R6487 VSS.n7642 VSS.n7641 292.5
R6488 VSS.n7639 VSS.n7620 292.5
R6489 VSS.n7620 VSS.n7619 292.5
R6490 VSS.n7638 VSS.n7637 292.5
R6491 VSS.n7637 VSS.n7636 292.5
R6492 VSS.n7622 VSS.n7621 292.5
R6493 VSS.n7635 VSS.n7622 292.5
R6494 VSS.n7633 VSS.n7632 292.5
R6495 VSS.n7634 VSS.n7633 292.5
R6496 VSS.n7631 VSS.n7624 292.5
R6497 VSS.n7624 VSS.n7623 292.5
R6498 VSS.n7630 VSS.n7629 292.5
R6499 VSS.n7629 VSS.n7628 292.5
R6500 VSS.n7626 VSS.n7625 292.5
R6501 VSS.n7627 VSS.n7626 292.5
R6502 VSS.n7521 VSS.n7520 292.5
R6503 VSS.n7523 VSS.n7521 292.5
R6504 VSS.n8222 VSS.n8221 292.5
R6505 VSS.n8221 VSS.n8220 292.5
R6506 VSS.n7868 VSS.n7867 292.5
R6507 VSS.n7869 VSS.n7868 292.5
R6508 VSS.n7656 VSS.n7655 292.5
R6509 VSS.n7870 VSS.n7656 292.5
R6510 VSS.n7873 VSS.n7872 292.5
R6511 VSS.n7872 VSS.n7871 292.5
R6512 VSS.n7874 VSS.n7654 292.5
R6513 VSS.n7654 VSS.n7653 292.5
R6514 VSS.n7876 VSS.n7875 292.5
R6515 VSS.n7877 VSS.n7876 292.5
R6516 VSS.n7652 VSS.n7651 292.5
R6517 VSS.n7878 VSS.n7652 292.5
R6518 VSS.n7881 VSS.n7880 292.5
R6519 VSS.n7880 VSS.n7879 292.5
R6520 VSS.n7882 VSS.n7650 292.5
R6521 VSS.n7650 VSS.n7649 292.5
R6522 VSS.n7884 VSS.n7883 292.5
R6523 VSS.n7885 VSS.n7884 292.5
R6524 VSS.n7648 VSS.n7647 292.5
R6525 VSS.n7886 VSS.n7648 292.5
R6526 VSS.n7889 VSS.n7888 292.5
R6527 VSS.n7888 VSS.n7887 292.5
R6528 VSS.n7866 VSS.n7658 292.5
R6529 VSS.n7658 VSS.n7657 292.5
R6530 VSS.n7750 VSS.n7743 292.5
R6531 VSS.n7751 VSS.n7750 292.5
R6532 VSS.n7761 VSS.n7760 292.5
R6533 VSS.n7762 VSS.n7761 292.5
R6534 VSS.n7733 VSS.n7731 292.5
R6535 VSS.n7735 VSS.n7733 292.5
R6536 VSS.n7725 VSS.n7724 292.5
R6537 VSS.n7774 VSS.n7725 292.5
R6538 VSS.n7784 VSS.n7783 292.5
R6539 VSS.n7785 VSS.n7784 292.5
R6540 VSS.n7714 VSS.n7712 292.5
R6541 VSS.n7716 VSS.n7714 292.5
R6542 VSS.n7706 VSS.n7705 292.5
R6543 VSS.n7796 VSS.n7706 292.5
R6544 VSS.n7806 VSS.n7805 292.5
R6545 VSS.n7807 VSS.n7806 292.5
R6546 VSS.n7695 VSS.n7693 292.5
R6547 VSS.n7697 VSS.n7695 292.5
R6548 VSS.n7687 VSS.n7686 292.5
R6549 VSS.n7819 VSS.n7687 292.5
R6550 VSS.n7829 VSS.n7828 292.5
R6551 VSS.n7830 VSS.n7829 292.5
R6552 VSS.n7835 VSS.n7674 292.5
R6553 VSS.n7674 VSS.n7673 292.5
R6554 VSS.n7841 VSS.n7840 292.5
R6555 VSS.n6831 VSS.n6830 292.5
R6556 VSS.n6830 VSS.n6829 292.5
R6557 VSS.n6850 VSS.n6849 292.5
R6558 VSS.n6851 VSS.n6850 292.5
R6559 VSS.n6848 VSS.n6747 292.5
R6560 VSS.n6747 VSS.n6746 292.5
R6561 VSS.n6847 VSS.n6846 292.5
R6562 VSS.n6846 VSS.n6845 292.5
R6563 VSS.n6749 VSS.n6748 292.5
R6564 VSS.n6844 VSS.n6749 292.5
R6565 VSS.n6842 VSS.n6841 292.5
R6566 VSS.n6843 VSS.n6842 292.5
R6567 VSS.n6840 VSS.n6751 292.5
R6568 VSS.n6751 VSS.n6750 292.5
R6569 VSS.n6839 VSS.n6838 292.5
R6570 VSS.n6838 VSS.n6837 292.5
R6571 VSS.n6753 VSS.n6752 292.5
R6572 VSS.n6836 VSS.n6753 292.5
R6573 VSS.n6834 VSS.n6833 292.5
R6574 VSS.n6835 VSS.n6834 292.5
R6575 VSS.n6832 VSS.n6755 292.5
R6576 VSS.n6755 VSS.n6754 292.5
R6577 VSS.n6745 VSS.n6744 292.5
R6578 VSS.n6852 VSS.n6745 292.5
R6579 VSS.n6758 VSS.n6756 292.5
R6580 VSS.n6802 VSS.n6801 292.5
R6581 VSS.n6803 VSS.n6802 292.5
R6582 VSS.n6826 VSS.n6825 292.5
R6583 VSS.n6827 VSS.n6826 292.5
R6584 VSS.n6824 VSS.n6760 292.5
R6585 VSS.n6760 VSS.n6759 292.5
R6586 VSS.n6823 VSS.n6822 292.5
R6587 VSS.n6822 VSS.n6821 292.5
R6588 VSS.n6762 VSS.n6761 292.5
R6589 VSS.n6820 VSS.n6762 292.5
R6590 VSS.n6818 VSS.n6817 292.5
R6591 VSS.n6819 VSS.n6818 292.5
R6592 VSS.n6816 VSS.n6764 292.5
R6593 VSS.n6764 VSS.n6763 292.5
R6594 VSS.n6815 VSS.n6814 292.5
R6595 VSS.n6814 VSS.n6813 292.5
R6596 VSS.n6768 VSS.n6765 292.5
R6597 VSS.n6812 VSS.n6765 292.5
R6598 VSS.n6810 VSS.n6809 292.5
R6599 VSS.n6811 VSS.n6810 292.5
R6600 VSS.n6808 VSS.n6767 292.5
R6601 VSS.n6767 VSS.n6766 292.5
R6602 VSS.n6807 VSS.n6806 292.5
R6603 VSS.n6806 VSS.n6805 292.5
R6604 VSS.n6770 VSS.n6769 292.5
R6605 VSS.n6804 VSS.n6770 292.5
R6606 VSS.n6800 VSS.n6772 292.5
R6607 VSS.n6772 VSS.n6771 292.5
R6608 VSS.n6799 VSS.n6798 292.5
R6609 VSS.n6798 VSS.n6797 292.5
R6610 VSS.n6774 VSS.n6773 292.5
R6611 VSS.n6796 VSS.n6774 292.5
R6612 VSS.n6794 VSS.n6793 292.5
R6613 VSS.n6795 VSS.n6794 292.5
R6614 VSS.n6792 VSS.n6776 292.5
R6615 VSS.n6776 VSS.n6775 292.5
R6616 VSS.n6791 VSS.n6790 292.5
R6617 VSS.n6790 VSS.n6789 292.5
R6618 VSS.n6778 VSS.n6777 292.5
R6619 VSS.n6788 VSS.n6778 292.5
R6620 VSS.n6786 VSS.n6785 292.5
R6621 VSS.n6787 VSS.n6786 292.5
R6622 VSS.n6784 VSS.n6780 292.5
R6623 VSS.n6780 VSS.n6779 292.5
R6624 VSS.n6783 VSS.n6782 292.5
R6625 VSS.n6782 VSS.n6781 292.5
R6626 VSS.n6731 VSS.n6730 292.5
R6627 VSS.n6733 VSS.n6731 292.5
R6628 VSS.n6879 VSS.n6878 292.5
R6629 VSS.n6878 VSS.n6877 292.5
R6630 VSS.n6855 VSS.n6854 292.5
R6631 VSS.n6854 VSS.n6853 292.5
R6632 VSS.n6856 VSS.n6743 292.5
R6633 VSS.n6743 VSS.n6742 292.5
R6634 VSS.n6858 VSS.n6857 292.5
R6635 VSS.n6859 VSS.n6858 292.5
R6636 VSS.n6741 VSS.n6740 292.5
R6637 VSS.n6860 VSS.n6741 292.5
R6638 VSS.n6863 VSS.n6862 292.5
R6639 VSS.n6862 VSS.n6861 292.5
R6640 VSS.n6864 VSS.n6739 292.5
R6641 VSS.n6739 VSS.n6738 292.5
R6642 VSS.n6866 VSS.n6865 292.5
R6643 VSS.n6867 VSS.n6866 292.5
R6644 VSS.n6737 VSS.n6736 292.5
R6645 VSS.n6868 VSS.n6737 292.5
R6646 VSS.n6871 VSS.n6870 292.5
R6647 VSS.n6870 VSS.n6869 292.5
R6648 VSS.n6872 VSS.n6735 292.5
R6649 VSS.n6735 VSS.n6734 292.5
R6650 VSS.n6874 VSS.n6873 292.5
R6651 VSS.n6875 VSS.n6874 292.5
R6652 VSS.n6732 VSS.n6729 292.5
R6653 VSS.n6876 VSS.n6732 292.5
R6654 VSS.n4242 VSS.n4241 292.5
R6655 VSS.n4241 VSS.n4178 292.5
R6656 VSS.n4220 VSS.n4219 292.5
R6657 VSS.n4221 VSS.n4220 292.5
R6658 VSS.n4188 VSS.n4187 292.5
R6659 VSS.n4222 VSS.n4188 292.5
R6660 VSS.n4225 VSS.n4224 292.5
R6661 VSS.n4224 VSS.n4223 292.5
R6662 VSS.n4226 VSS.n4186 292.5
R6663 VSS.n4186 VSS.n4185 292.5
R6664 VSS.n4228 VSS.n4227 292.5
R6665 VSS.n4229 VSS.n4228 292.5
R6666 VSS.n4184 VSS.n4183 292.5
R6667 VSS.n4230 VSS.n4184 292.5
R6668 VSS.n4233 VSS.n4232 292.5
R6669 VSS.n4232 VSS.n4231 292.5
R6670 VSS.n4234 VSS.n4181 292.5
R6671 VSS.n4181 VSS.n4180 292.5
R6672 VSS.n4236 VSS.n4235 292.5
R6673 VSS.n4237 VSS.n4236 292.5
R6674 VSS.n4182 VSS.n4179 292.5
R6675 VSS.n4238 VSS.n4179 292.5
R6676 VSS.n4240 VSS.n4177 292.5
R6677 VSS.n4240 VSS.n4239 292.5
R6678 VSS.n3639 VSS.n3637 292.5
R6679 VSS.n3641 VSS.n3639 292.5
R6680 VSS.n3644 VSS.n3640 292.5
R6681 VSS.n5658 VSS.n3640 292.5
R6682 VSS.n5567 VSS.n5566 292.5
R6683 VSS.n5567 VSS.n5416 292.5
R6684 VSS.n5421 VSS.n5420 292.5
R6685 VSS.n5557 VSS.n5421 292.5
R6686 VSS.n5430 VSS.n5428 292.5
R6687 VSS.n5432 VSS.n5430 292.5
R6688 VSS.n5544 VSS.n5543 292.5
R6689 VSS.n5545 VSS.n5544 292.5
R6690 VSS.n5441 VSS.n5440 292.5
R6691 VSS.n5534 VSS.n5441 292.5
R6692 VSS.n5449 VSS.n5447 292.5
R6693 VSS.n5451 VSS.n5449 292.5
R6694 VSS.n5521 VSS.n5520 292.5
R6695 VSS.n5522 VSS.n5521 292.5
R6696 VSS.n5460 VSS.n5459 292.5
R6697 VSS.n5512 VSS.n5460 292.5
R6698 VSS.n5468 VSS.n5466 292.5
R6699 VSS.n5470 VSS.n5468 292.5
R6700 VSS.n5499 VSS.n5498 292.5
R6701 VSS.n5500 VSS.n5499 292.5
R6702 VSS.n5479 VSS.n5478 292.5
R6703 VSS.n5489 VSS.n5479 292.5
R6704 VSS.n5654 VSS.n3643 292.5
R6705 VSS.n3643 VSS.n3642 292.5
R6706 VSS.n5653 VSS.n5652 292.5
R6707 VSS.n5652 VSS.n5651 292.5
R6708 VSS.n3650 VSS.n3649 292.5
R6709 VSS.n5650 VSS.n3650 292.5
R6710 VSS.n5648 VSS.n5647 292.5
R6711 VSS.n5649 VSS.n5648 292.5
R6712 VSS.n5646 VSS.n3652 292.5
R6713 VSS.n3652 VSS.n3651 292.5
R6714 VSS.n5645 VSS.n5644 292.5
R6715 VSS.n5644 VSS.n5643 292.5
R6716 VSS.n3654 VSS.n3653 292.5
R6717 VSS.n5642 VSS.n3654 292.5
R6718 VSS.n5640 VSS.n5639 292.5
R6719 VSS.n5641 VSS.n5640 292.5
R6720 VSS.n5638 VSS.n3656 292.5
R6721 VSS.n3656 VSS.n3655 292.5
R6722 VSS.n5637 VSS.n5636 292.5
R6723 VSS.n5636 VSS.n5635 292.5
R6724 VSS.n3658 VSS.n3657 292.5
R6725 VSS.n5634 VSS.n3658 292.5
R6726 VSS.n5656 VSS.n5655 292.5
R6727 VSS.n5657 VSS.n5656 292.5
R6728 VSS.n3670 VSS.n3669 292.5
R6729 VSS.n5610 VSS.n3670 292.5
R6730 VSS.n5613 VSS.n5612 292.5
R6731 VSS.n5612 VSS.n5611 292.5
R6732 VSS.n5614 VSS.n3668 292.5
R6733 VSS.n3668 VSS.n3667 292.5
R6734 VSS.n5616 VSS.n5615 292.5
R6735 VSS.n5617 VSS.n5616 292.5
R6736 VSS.n3666 VSS.n3665 292.5
R6737 VSS.n5618 VSS.n3666 292.5
R6738 VSS.n5621 VSS.n5620 292.5
R6739 VSS.n5620 VSS.n5619 292.5
R6740 VSS.n5622 VSS.n3664 292.5
R6741 VSS.n3664 VSS.n3663 292.5
R6742 VSS.n5624 VSS.n5623 292.5
R6743 VSS.n5625 VSS.n5624 292.5
R6744 VSS.n3662 VSS.n3661 292.5
R6745 VSS.n5626 VSS.n3662 292.5
R6746 VSS.n5629 VSS.n5628 292.5
R6747 VSS.n5628 VSS.n5627 292.5
R6748 VSS.n5630 VSS.n3660 292.5
R6749 VSS.n3660 VSS.n3659 292.5
R6750 VSS.n5632 VSS.n5631 292.5
R6751 VSS.n5633 VSS.n5632 292.5
R6752 VSS.n3798 VSS.n3797 292.5
R6753 VSS.n3799 VSS.n3798 292.5
R6754 VSS.n3796 VSS.n3771 292.5
R6755 VSS.n3771 VSS.n3770 292.5
R6756 VSS.n3795 VSS.n3794 292.5
R6757 VSS.n3794 VSS.n3793 292.5
R6758 VSS.n3773 VSS.n3772 292.5
R6759 VSS.n3792 VSS.n3773 292.5
R6760 VSS.n3790 VSS.n3789 292.5
R6761 VSS.n3791 VSS.n3790 292.5
R6762 VSS.n3788 VSS.n3775 292.5
R6763 VSS.n3775 VSS.n3774 292.5
R6764 VSS.n3787 VSS.n3786 292.5
R6765 VSS.n3786 VSS.n3785 292.5
R6766 VSS.n3777 VSS.n3776 292.5
R6767 VSS.n3784 VSS.n3777 292.5
R6768 VSS.n3782 VSS.n3781 292.5
R6769 VSS.n3783 VSS.n3782 292.5
R6770 VSS.n3780 VSS.n3779 292.5
R6771 VSS.n3779 VSS.n3778 292.5
R6772 VSS.n3675 VSS.n3673 292.5
R6773 VSS.n3673 VSS.n3672 292.5
R6774 VSS.n5607 VSS.n5606 292.5
R6775 VSS.n5608 VSS.n5607 292.5
R6776 VSS.n3693 VSS.n3692 292.5
R6777 VSS.n5415 VSS.n3693 292.5
R6778 VSS.n3702 VSS.n3700 292.5
R6779 VSS.n5402 VSS.n3702 292.5
R6780 VSS.n5399 VSS.n5398 292.5
R6781 VSS.n5400 VSS.n5399 292.5
R6782 VSS.n3709 VSS.n3707 292.5
R6783 VSS.n5389 VSS.n3709 292.5
R6784 VSS.n5380 VSS.n5379 292.5
R6785 VSS.n5379 VSS.n5378 292.5
R6786 VSS.n3718 VSS.n3717 292.5
R6787 VSS.n3717 VSS.n3716 292.5
R6788 VSS.n5365 VSS.n5364 292.5
R6789 VSS.n5366 VSS.n5365 292.5
R6790 VSS.n3730 VSS.n3728 292.5
R6791 VSS.n5355 VSS.n3730 292.5
R6792 VSS.n5346 VSS.n5345 292.5
R6793 VSS.n5345 VSS.n5344 292.5
R6794 VSS.n3739 VSS.n3738 292.5
R6795 VSS.n3738 VSS.n3737 292.5
R6796 VSS.n5330 VSS.n5329 292.5
R6797 VSS.n5331 VSS.n5330 292.5
R6798 VSS.n3751 VSS.n3749 292.5
R6799 VSS.n5320 VSS.n3751 292.5
R6800 VSS.n5131 VSS.n5129 292.5
R6801 VSS.n5132 VSS.n5131 292.5
R6802 VSS.n5122 VSS.n5121 292.5
R6803 VSS.n5143 VSS.n5122 292.5
R6804 VSS.n5153 VSS.n5152 292.5
R6805 VSS.n5154 VSS.n5153 292.5
R6806 VSS.n5111 VSS.n5109 292.5
R6807 VSS.n5113 VSS.n5111 292.5
R6808 VSS.n5103 VSS.n5102 292.5
R6809 VSS.n5166 VSS.n5103 292.5
R6810 VSS.n5175 VSS.n5174 292.5
R6811 VSS.n5176 VSS.n5175 292.5
R6812 VSS.n5092 VSS.n5090 292.5
R6813 VSS.n5094 VSS.n5092 292.5
R6814 VSS.n5084 VSS.n5083 292.5
R6815 VSS.n5188 VSS.n5084 292.5
R6816 VSS.n5198 VSS.n5197 292.5
R6817 VSS.n5199 VSS.n5198 292.5
R6818 VSS.n5073 VSS.n5071 292.5
R6819 VSS.n5075 VSS.n5073 292.5
R6820 VSS.n5064 VSS.n5063 292.5
R6821 VSS.n5211 VSS.n5064 292.5
R6822 VSS.n5221 VSS.n5220 292.5
R6823 VSS.n5221 VSS.n5059 292.5
R6824 VSS.n3811 VSS.n3810 292.5
R6825 VSS.n5264 VSS.n3811 292.5
R6826 VSS.n5267 VSS.n5266 292.5
R6827 VSS.n5266 VSS.n5265 292.5
R6828 VSS.n5268 VSS.n3809 292.5
R6829 VSS.n3809 VSS.n3808 292.5
R6830 VSS.n5270 VSS.n5269 292.5
R6831 VSS.n5271 VSS.n5270 292.5
R6832 VSS.n3807 VSS.n3806 292.5
R6833 VSS.n5272 VSS.n3807 292.5
R6834 VSS.n5275 VSS.n5274 292.5
R6835 VSS.n5274 VSS.n5273 292.5
R6836 VSS.n5276 VSS.n3805 292.5
R6837 VSS.n3805 VSS.n3804 292.5
R6838 VSS.n5278 VSS.n5277 292.5
R6839 VSS.n5279 VSS.n5278 292.5
R6840 VSS.n3803 VSS.n3802 292.5
R6841 VSS.n5280 VSS.n3803 292.5
R6842 VSS.n5283 VSS.n5282 292.5
R6843 VSS.n5282 VSS.n5281 292.5
R6844 VSS.n5284 VSS.n3801 292.5
R6845 VSS.n3801 VSS.n3800 292.5
R6846 VSS.n5286 VSS.n5285 292.5
R6847 VSS.n5287 VSS.n5286 292.5
R6848 VSS.n3939 VSS.n3938 292.5
R6849 VSS.n3940 VSS.n3939 292.5
R6850 VSS.n3937 VSS.n3912 292.5
R6851 VSS.n3912 VSS.n3911 292.5
R6852 VSS.n3936 VSS.n3935 292.5
R6853 VSS.n3935 VSS.n3934 292.5
R6854 VSS.n3914 VSS.n3913 292.5
R6855 VSS.n3933 VSS.n3914 292.5
R6856 VSS.n3931 VSS.n3930 292.5
R6857 VSS.n3932 VSS.n3931 292.5
R6858 VSS.n3929 VSS.n3916 292.5
R6859 VSS.n3916 VSS.n3915 292.5
R6860 VSS.n3928 VSS.n3927 292.5
R6861 VSS.n3927 VSS.n3926 292.5
R6862 VSS.n3918 VSS.n3917 292.5
R6863 VSS.n3925 VSS.n3918 292.5
R6864 VSS.n3923 VSS.n3922 292.5
R6865 VSS.n3924 VSS.n3923 292.5
R6866 VSS.n3921 VSS.n3920 292.5
R6867 VSS.n3920 VSS.n3919 292.5
R6868 VSS.n3816 VSS.n3814 292.5
R6869 VSS.n3814 VSS.n3813 292.5
R6870 VSS.n5261 VSS.n5260 292.5
R6871 VSS.n5262 VSS.n5261 292.5
R6872 VSS.n3834 VSS.n3833 292.5
R6873 VSS.n5058 VSS.n3834 292.5
R6874 VSS.n3843 VSS.n3841 292.5
R6875 VSS.n5045 VSS.n3843 292.5
R6876 VSS.n5042 VSS.n5041 292.5
R6877 VSS.n5043 VSS.n5042 292.5
R6878 VSS.n3850 VSS.n3848 292.5
R6879 VSS.n5032 VSS.n3850 292.5
R6880 VSS.n5023 VSS.n5022 292.5
R6881 VSS.n5022 VSS.n5021 292.5
R6882 VSS.n3859 VSS.n3858 292.5
R6883 VSS.n3858 VSS.n3857 292.5
R6884 VSS.n5008 VSS.n5007 292.5
R6885 VSS.n5009 VSS.n5008 292.5
R6886 VSS.n3871 VSS.n3869 292.5
R6887 VSS.n4998 VSS.n3871 292.5
R6888 VSS.n4989 VSS.n4988 292.5
R6889 VSS.n4988 VSS.n4987 292.5
R6890 VSS.n3880 VSS.n3879 292.5
R6891 VSS.n3879 VSS.n3878 292.5
R6892 VSS.n4973 VSS.n4972 292.5
R6893 VSS.n4974 VSS.n4973 292.5
R6894 VSS.n3892 VSS.n3890 292.5
R6895 VSS.n4963 VSS.n3892 292.5
R6896 VSS.n4774 VSS.n4772 292.5
R6897 VSS.n4775 VSS.n4774 292.5
R6898 VSS.n4765 VSS.n4764 292.5
R6899 VSS.n4786 VSS.n4765 292.5
R6900 VSS.n4796 VSS.n4795 292.5
R6901 VSS.n4797 VSS.n4796 292.5
R6902 VSS.n4754 VSS.n4752 292.5
R6903 VSS.n4756 VSS.n4754 292.5
R6904 VSS.n4746 VSS.n4745 292.5
R6905 VSS.n4809 VSS.n4746 292.5
R6906 VSS.n4818 VSS.n4817 292.5
R6907 VSS.n4819 VSS.n4818 292.5
R6908 VSS.n4735 VSS.n4733 292.5
R6909 VSS.n4737 VSS.n4735 292.5
R6910 VSS.n4727 VSS.n4726 292.5
R6911 VSS.n4831 VSS.n4727 292.5
R6912 VSS.n4841 VSS.n4840 292.5
R6913 VSS.n4842 VSS.n4841 292.5
R6914 VSS.n4716 VSS.n4714 292.5
R6915 VSS.n4718 VSS.n4716 292.5
R6916 VSS.n4707 VSS.n4706 292.5
R6917 VSS.n4854 VSS.n4707 292.5
R6918 VSS.n4864 VSS.n4863 292.5
R6919 VSS.n4864 VSS.n4702 292.5
R6920 VSS.n3952 VSS.n3951 292.5
R6921 VSS.n4907 VSS.n3952 292.5
R6922 VSS.n4910 VSS.n4909 292.5
R6923 VSS.n4909 VSS.n4908 292.5
R6924 VSS.n4911 VSS.n3950 292.5
R6925 VSS.n3950 VSS.n3949 292.5
R6926 VSS.n4913 VSS.n4912 292.5
R6927 VSS.n4914 VSS.n4913 292.5
R6928 VSS.n3948 VSS.n3947 292.5
R6929 VSS.n4915 VSS.n3948 292.5
R6930 VSS.n4918 VSS.n4917 292.5
R6931 VSS.n4917 VSS.n4916 292.5
R6932 VSS.n4919 VSS.n3946 292.5
R6933 VSS.n3946 VSS.n3945 292.5
R6934 VSS.n4921 VSS.n4920 292.5
R6935 VSS.n4922 VSS.n4921 292.5
R6936 VSS.n3944 VSS.n3943 292.5
R6937 VSS.n4923 VSS.n3944 292.5
R6938 VSS.n4926 VSS.n4925 292.5
R6939 VSS.n4925 VSS.n4924 292.5
R6940 VSS.n4927 VSS.n3942 292.5
R6941 VSS.n3942 VSS.n3941 292.5
R6942 VSS.n4929 VSS.n4928 292.5
R6943 VSS.n4930 VSS.n4929 292.5
R6944 VSS.n4080 VSS.n4079 292.5
R6945 VSS.n4081 VSS.n4080 292.5
R6946 VSS.n4078 VSS.n4053 292.5
R6947 VSS.n4053 VSS.n4052 292.5
R6948 VSS.n4077 VSS.n4076 292.5
R6949 VSS.n4076 VSS.n4075 292.5
R6950 VSS.n4055 VSS.n4054 292.5
R6951 VSS.n4074 VSS.n4055 292.5
R6952 VSS.n4072 VSS.n4071 292.5
R6953 VSS.n4073 VSS.n4072 292.5
R6954 VSS.n4070 VSS.n4057 292.5
R6955 VSS.n4057 VSS.n4056 292.5
R6956 VSS.n4069 VSS.n4068 292.5
R6957 VSS.n4068 VSS.n4067 292.5
R6958 VSS.n4059 VSS.n4058 292.5
R6959 VSS.n4066 VSS.n4059 292.5
R6960 VSS.n4064 VSS.n4063 292.5
R6961 VSS.n4065 VSS.n4064 292.5
R6962 VSS.n4062 VSS.n4061 292.5
R6963 VSS.n4061 VSS.n4060 292.5
R6964 VSS.n3957 VSS.n3955 292.5
R6965 VSS.n3955 VSS.n3954 292.5
R6966 VSS.n4904 VSS.n4903 292.5
R6967 VSS.n4905 VSS.n4904 292.5
R6968 VSS.n3975 VSS.n3974 292.5
R6969 VSS.n4701 VSS.n3975 292.5
R6970 VSS.n3984 VSS.n3982 292.5
R6971 VSS.n4688 VSS.n3984 292.5
R6972 VSS.n4685 VSS.n4684 292.5
R6973 VSS.n4686 VSS.n4685 292.5
R6974 VSS.n3991 VSS.n3989 292.5
R6975 VSS.n4675 VSS.n3991 292.5
R6976 VSS.n4666 VSS.n4665 292.5
R6977 VSS.n4665 VSS.n4664 292.5
R6978 VSS.n4000 VSS.n3999 292.5
R6979 VSS.n3999 VSS.n3998 292.5
R6980 VSS.n4651 VSS.n4650 292.5
R6981 VSS.n4652 VSS.n4651 292.5
R6982 VSS.n4012 VSS.n4010 292.5
R6983 VSS.n4641 VSS.n4012 292.5
R6984 VSS.n4632 VSS.n4631 292.5
R6985 VSS.n4631 VSS.n4630 292.5
R6986 VSS.n4021 VSS.n4020 292.5
R6987 VSS.n4020 VSS.n4019 292.5
R6988 VSS.n4616 VSS.n4615 292.5
R6989 VSS.n4617 VSS.n4616 292.5
R6990 VSS.n4033 VSS.n4031 292.5
R6991 VSS.n4606 VSS.n4033 292.5
R6992 VSS.n4417 VSS.n4415 292.5
R6993 VSS.n4418 VSS.n4417 292.5
R6994 VSS.n4408 VSS.n4407 292.5
R6995 VSS.n4429 VSS.n4408 292.5
R6996 VSS.n4439 VSS.n4438 292.5
R6997 VSS.n4440 VSS.n4439 292.5
R6998 VSS.n4397 VSS.n4395 292.5
R6999 VSS.n4399 VSS.n4397 292.5
R7000 VSS.n4389 VSS.n4388 292.5
R7001 VSS.n4452 VSS.n4389 292.5
R7002 VSS.n4461 VSS.n4460 292.5
R7003 VSS.n4462 VSS.n4461 292.5
R7004 VSS.n4378 VSS.n4376 292.5
R7005 VSS.n4380 VSS.n4378 292.5
R7006 VSS.n4370 VSS.n4369 292.5
R7007 VSS.n4474 VSS.n4370 292.5
R7008 VSS.n4484 VSS.n4483 292.5
R7009 VSS.n4485 VSS.n4484 292.5
R7010 VSS.n4359 VSS.n4357 292.5
R7011 VSS.n4361 VSS.n4359 292.5
R7012 VSS.n4350 VSS.n4349 292.5
R7013 VSS.n4497 VSS.n4350 292.5
R7014 VSS.n4507 VSS.n4506 292.5
R7015 VSS.n4507 VSS.n4345 292.5
R7016 VSS.n4093 VSS.n4092 292.5
R7017 VSS.n4550 VSS.n4093 292.5
R7018 VSS.n4553 VSS.n4552 292.5
R7019 VSS.n4552 VSS.n4551 292.5
R7020 VSS.n4554 VSS.n4091 292.5
R7021 VSS.n4091 VSS.n4090 292.5
R7022 VSS.n4556 VSS.n4555 292.5
R7023 VSS.n4557 VSS.n4556 292.5
R7024 VSS.n4089 VSS.n4088 292.5
R7025 VSS.n4558 VSS.n4089 292.5
R7026 VSS.n4561 VSS.n4560 292.5
R7027 VSS.n4560 VSS.n4559 292.5
R7028 VSS.n4562 VSS.n4087 292.5
R7029 VSS.n4087 VSS.n4086 292.5
R7030 VSS.n4564 VSS.n4563 292.5
R7031 VSS.n4565 VSS.n4564 292.5
R7032 VSS.n4085 VSS.n4084 292.5
R7033 VSS.n4566 VSS.n4085 292.5
R7034 VSS.n4569 VSS.n4568 292.5
R7035 VSS.n4568 VSS.n4567 292.5
R7036 VSS.n4570 VSS.n4083 292.5
R7037 VSS.n4083 VSS.n4082 292.5
R7038 VSS.n4572 VSS.n4571 292.5
R7039 VSS.n4573 VSS.n4572 292.5
R7040 VSS.n4217 VSS.n4216 292.5
R7041 VSS.n4216 VSS.n4215 292.5
R7042 VSS.n4192 VSS.n4191 292.5
R7043 VSS.n4214 VSS.n4192 292.5
R7044 VSS.n4212 VSS.n4211 292.5
R7045 VSS.n4213 VSS.n4212 292.5
R7046 VSS.n4210 VSS.n4194 292.5
R7047 VSS.n4194 VSS.n4193 292.5
R7048 VSS.n4209 VSS.n4208 292.5
R7049 VSS.n4208 VSS.n4207 292.5
R7050 VSS.n4196 VSS.n4195 292.5
R7051 VSS.n4206 VSS.n4196 292.5
R7052 VSS.n4204 VSS.n4203 292.5
R7053 VSS.n4205 VSS.n4204 292.5
R7054 VSS.n4202 VSS.n4198 292.5
R7055 VSS.n4198 VSS.n4197 292.5
R7056 VSS.n4201 VSS.n4200 292.5
R7057 VSS.n4200 VSS.n4199 292.5
R7058 VSS.n4098 VSS.n4096 292.5
R7059 VSS.n4096 VSS.n4095 292.5
R7060 VSS.n4547 VSS.n4546 292.5
R7061 VSS.n4548 VSS.n4547 292.5
R7062 VSS.n4218 VSS.n4190 292.5
R7063 VSS.n4190 VSS.n4189 292.5
R7064 VSS.n4116 VSS.n4115 292.5
R7065 VSS.n4344 VSS.n4116 292.5
R7066 VSS.n4125 VSS.n4123 292.5
R7067 VSS.n4331 VSS.n4125 292.5
R7068 VSS.n4328 VSS.n4327 292.5
R7069 VSS.n4329 VSS.n4328 292.5
R7070 VSS.n4132 VSS.n4130 292.5
R7071 VSS.n4318 VSS.n4132 292.5
R7072 VSS.n4309 VSS.n4308 292.5
R7073 VSS.n4308 VSS.n4307 292.5
R7074 VSS.n4141 VSS.n4140 292.5
R7075 VSS.n4140 VSS.n4139 292.5
R7076 VSS.n4294 VSS.n4293 292.5
R7077 VSS.n4295 VSS.n4294 292.5
R7078 VSS.n4153 VSS.n4151 292.5
R7079 VSS.n4284 VSS.n4153 292.5
R7080 VSS.n4275 VSS.n4274 292.5
R7081 VSS.n4274 VSS.n4273 292.5
R7082 VSS.n4162 VSS.n4161 292.5
R7083 VSS.n4161 VSS.n4160 292.5
R7084 VSS.n4259 VSS.n4258 292.5
R7085 VSS.n4260 VSS.n4259 292.5
R7086 VSS.n4174 VSS.n4172 292.5
R7087 VSS.n4249 VSS.n4174 292.5
R7088 VSS.n4244 VSS.n4243 292.5
R7089 VSS.n1969 VSS.n1968 292.5
R7090 VSS.n1968 VSS.n1967 292.5
R7091 VSS.n1592 VSS.n1591 292.5
R7092 VSS.n1990 VSS.n1592 292.5
R7093 VSS.n1988 VSS.n1987 292.5
R7094 VSS.n1989 VSS.n1988 292.5
R7095 VSS.n1986 VSS.n1594 292.5
R7096 VSS.n1594 VSS.n1593 292.5
R7097 VSS.n1985 VSS.n1984 292.5
R7098 VSS.n1984 VSS.n1983 292.5
R7099 VSS.n1596 VSS.n1595 292.5
R7100 VSS.n1982 VSS.n1596 292.5
R7101 VSS.n1980 VSS.n1979 292.5
R7102 VSS.n1981 VSS.n1980 292.5
R7103 VSS.n1978 VSS.n1598 292.5
R7104 VSS.n1598 VSS.n1597 292.5
R7105 VSS.n1977 VSS.n1976 292.5
R7106 VSS.n1976 VSS.n1975 292.5
R7107 VSS.n1600 VSS.n1599 292.5
R7108 VSS.n1974 VSS.n1600 292.5
R7109 VSS.n1972 VSS.n1971 292.5
R7110 VSS.n1973 VSS.n1972 292.5
R7111 VSS.n1970 VSS.n1602 292.5
R7112 VSS.n1602 VSS.n1601 292.5
R7113 VSS.n1284 VSS.n1283 292.5
R7114 VSS.n3017 VSS.n1284 292.5
R7115 VSS.n2996 VSS.n2995 292.5
R7116 VSS.n2995 VSS.n2994 292.5
R7117 VSS.n2997 VSS.n1294 292.5
R7118 VSS.n1294 VSS.n1293 292.5
R7119 VSS.n2999 VSS.n2998 292.5
R7120 VSS.n3000 VSS.n2999 292.5
R7121 VSS.n1292 VSS.n1291 292.5
R7122 VSS.n3001 VSS.n1292 292.5
R7123 VSS.n3004 VSS.n3003 292.5
R7124 VSS.n3003 VSS.n3002 292.5
R7125 VSS.n3005 VSS.n1290 292.5
R7126 VSS.n1290 VSS.n1289 292.5
R7127 VSS.n3007 VSS.n3006 292.5
R7128 VSS.n3008 VSS.n3007 292.5
R7129 VSS.n1288 VSS.n1287 292.5
R7130 VSS.n3009 VSS.n1288 292.5
R7131 VSS.n3012 VSS.n3011 292.5
R7132 VSS.n3011 VSS.n3010 292.5
R7133 VSS.n3013 VSS.n1286 292.5
R7134 VSS.n1286 VSS.n1285 292.5
R7135 VSS.n3015 VSS.n3014 292.5
R7136 VSS.n3016 VSS.n3015 292.5
R7137 VSS.n3039 VSS.n3038 292.5
R7138 VSS.n3040 VSS.n3039 292.5
R7139 VSS.n3037 VSS.n1274 292.5
R7140 VSS.n1274 VSS.n1273 292.5
R7141 VSS.n3036 VSS.n3035 292.5
R7142 VSS.n3035 VSS.n3034 292.5
R7143 VSS.n1276 VSS.n1275 292.5
R7144 VSS.n3033 VSS.n1276 292.5
R7145 VSS.n3031 VSS.n3030 292.5
R7146 VSS.n3032 VSS.n3031 292.5
R7147 VSS.n3029 VSS.n1278 292.5
R7148 VSS.n1278 VSS.n1277 292.5
R7149 VSS.n3028 VSS.n3027 292.5
R7150 VSS.n3027 VSS.n3026 292.5
R7151 VSS.n1280 VSS.n1279 292.5
R7152 VSS.n3025 VSS.n1280 292.5
R7153 VSS.n3023 VSS.n3022 292.5
R7154 VSS.n3024 VSS.n3023 292.5
R7155 VSS.n3021 VSS.n1282 292.5
R7156 VSS.n1282 VSS.n1281 292.5
R7157 VSS.n3020 VSS.n3019 292.5
R7158 VSS.n3019 VSS.n3018 292.5
R7159 VSS.n1271 VSS.n1268 292.5
R7160 VSS.n3041 VSS.n1271 292.5
R7161 VSS.n3044 VSS.n3043 292.5
R7162 VSS.n3043 VSS.n3042 292.5
R7163 VSS.n2804 VSS.n2802 292.5
R7164 VSS.n2808 VSS.n2804 292.5
R7165 VSS.n2957 VSS.n2956 292.5
R7166 VSS.n2958 VSS.n2957 292.5
R7167 VSS.n2817 VSS.n2816 292.5
R7168 VSS.n2947 VSS.n2817 292.5
R7169 VSS.n2825 VSS.n2823 292.5
R7170 VSS.n2827 VSS.n2825 292.5
R7171 VSS.n2934 VSS.n2933 292.5
R7172 VSS.n2935 VSS.n2934 292.5
R7173 VSS.n2836 VSS.n2835 292.5
R7174 VSS.n2924 VSS.n2836 292.5
R7175 VSS.n2844 VSS.n2842 292.5
R7176 VSS.n2846 VSS.n2844 292.5
R7177 VSS.n2912 VSS.n2911 292.5
R7178 VSS.n2913 VSS.n2912 292.5
R7179 VSS.n2855 VSS.n2854 292.5
R7180 VSS.n2902 VSS.n2855 292.5
R7181 VSS.n2863 VSS.n2861 292.5
R7182 VSS.n2865 VSS.n2863 292.5
R7183 VSS.n2889 VSS.n2888 292.5
R7184 VSS.n2890 VSS.n2889 292.5
R7185 VSS.n2878 VSS.n2877 292.5
R7186 VSS.n2879 VSS.n2878 292.5
R7187 VSS.n1316 VSS.n1315 292.5
R7188 VSS.n2794 VSS.n1316 292.5
R7189 VSS.n2785 VSS.n2784 292.5
R7190 VSS.n2784 VSS.n2783 292.5
R7191 VSS.n1325 VSS.n1324 292.5
R7192 VSS.n1324 VSS.n1323 292.5
R7193 VSS.n2769 VSS.n2768 292.5
R7194 VSS.n2770 VSS.n2769 292.5
R7195 VSS.n1337 VSS.n1335 292.5
R7196 VSS.n2759 VSS.n1337 292.5
R7197 VSS.n2751 VSS.n2750 292.5
R7198 VSS.n2750 VSS.n2749 292.5
R7199 VSS.n1346 VSS.n1345 292.5
R7200 VSS.n1345 VSS.n1344 292.5
R7201 VSS.n2735 VSS.n2734 292.5
R7202 VSS.n2736 VSS.n2735 292.5
R7203 VSS.n1358 VSS.n1356 292.5
R7204 VSS.n2725 VSS.n1358 292.5
R7205 VSS.n2716 VSS.n2715 292.5
R7206 VSS.n2715 VSS.n2714 292.5
R7207 VSS.n1367 VSS.n1366 292.5
R7208 VSS.n1366 VSS.n1365 292.5
R7209 VSS.n2700 VSS.n2699 292.5
R7210 VSS.n2701 VSS.n2700 292.5
R7211 VSS.n1433 VSS.n1432 292.5
R7212 VSS.n1434 VSS.n1433 292.5
R7213 VSS.n1431 VSS.n1401 292.5
R7214 VSS.n1401 VSS.n1400 292.5
R7215 VSS.n1430 VSS.n1429 292.5
R7216 VSS.n1429 VSS.n1428 292.5
R7217 VSS.n1403 VSS.n1402 292.5
R7218 VSS.n1427 VSS.n1403 292.5
R7219 VSS.n1425 VSS.n1424 292.5
R7220 VSS.n1426 VSS.n1425 292.5
R7221 VSS.n1423 VSS.n1405 292.5
R7222 VSS.n1405 VSS.n1404 292.5
R7223 VSS.n1422 VSS.n1421 292.5
R7224 VSS.n1421 VSS.n1420 292.5
R7225 VSS.n1407 VSS.n1406 292.5
R7226 VSS.n1419 VSS.n1407 292.5
R7227 VSS.n1417 VSS.n1416 292.5
R7228 VSS.n1418 VSS.n1417 292.5
R7229 VSS.n1415 VSS.n1409 292.5
R7230 VSS.n1409 VSS.n1408 292.5
R7231 VSS.n1414 VSS.n1413 292.5
R7232 VSS.n1413 VSS.n1412 292.5
R7233 VSS.n1411 VSS.n1410 292.5
R7234 VSS.n1411 VSS.n1297 292.5
R7235 VSS.n1446 VSS.n1445 292.5
R7236 VSS.n2631 VSS.n1446 292.5
R7237 VSS.n2634 VSS.n2633 292.5
R7238 VSS.n2633 VSS.n2632 292.5
R7239 VSS.n2635 VSS.n1444 292.5
R7240 VSS.n1444 VSS.n1443 292.5
R7241 VSS.n2637 VSS.n2636 292.5
R7242 VSS.n2638 VSS.n2637 292.5
R7243 VSS.n1442 VSS.n1441 292.5
R7244 VSS.n2639 VSS.n1442 292.5
R7245 VSS.n2642 VSS.n2641 292.5
R7246 VSS.n2641 VSS.n2640 292.5
R7247 VSS.n2643 VSS.n1440 292.5
R7248 VSS.n1440 VSS.n1439 292.5
R7249 VSS.n2645 VSS.n2644 292.5
R7250 VSS.n2646 VSS.n2645 292.5
R7251 VSS.n1438 VSS.n1437 292.5
R7252 VSS.n2647 VSS.n1438 292.5
R7253 VSS.n2650 VSS.n2649 292.5
R7254 VSS.n2649 VSS.n2648 292.5
R7255 VSS.n2651 VSS.n1436 292.5
R7256 VSS.n1436 VSS.n1435 292.5
R7257 VSS.n2653 VSS.n2652 292.5
R7258 VSS.n2654 VSS.n2653 292.5
R7259 VSS.n1383 VSS.n1381 292.5
R7260 VSS.n2685 VSS.n1383 292.5
R7261 VSS.n2397 VSS.n2396 292.5
R7262 VSS.n2398 VSS.n2397 292.5
R7263 VSS.n2388 VSS.n2386 292.5
R7264 VSS.n2390 VSS.n2388 292.5
R7265 VSS.n2380 VSS.n2379 292.5
R7266 VSS.n2410 VSS.n2380 292.5
R7267 VSS.n2420 VSS.n2419 292.5
R7268 VSS.n2421 VSS.n2420 292.5
R7269 VSS.n2369 VSS.n2367 292.5
R7270 VSS.n2371 VSS.n2369 292.5
R7271 VSS.n2361 VSS.n2360 292.5
R7272 VSS.n2432 VSS.n2361 292.5
R7273 VSS.n2442 VSS.n2441 292.5
R7274 VSS.n2443 VSS.n2442 292.5
R7275 VSS.n2350 VSS.n2348 292.5
R7276 VSS.n2352 VSS.n2350 292.5
R7277 VSS.n2342 VSS.n2341 292.5
R7278 VSS.n2455 VSS.n2342 292.5
R7279 VSS.n2465 VSS.n2464 292.5
R7280 VSS.n2466 VSS.n2465 292.5
R7281 VSS.n2328 VSS.n2326 292.5
R7282 VSS.n2333 VSS.n2328 292.5
R7283 VSS.n2287 VSS.n2286 292.5
R7284 VSS.n2479 VSS.n2287 292.5
R7285 VSS.n2489 VSS.n2488 292.5
R7286 VSS.n2490 VSS.n2489 292.5
R7287 VSS.n2276 VSS.n2274 292.5
R7288 VSS.n2278 VSS.n2276 292.5
R7289 VSS.n2268 VSS.n2267 292.5
R7290 VSS.n2502 VSS.n2268 292.5
R7291 VSS.n2512 VSS.n2511 292.5
R7292 VSS.n2513 VSS.n2512 292.5
R7293 VSS.n2257 VSS.n2255 292.5
R7294 VSS.n2259 VSS.n2257 292.5
R7295 VSS.n2249 VSS.n2248 292.5
R7296 VSS.n2524 VSS.n2249 292.5
R7297 VSS.n2534 VSS.n2533 292.5
R7298 VSS.n2535 VSS.n2534 292.5
R7299 VSS.n2238 VSS.n2236 292.5
R7300 VSS.n2240 VSS.n2238 292.5
R7301 VSS.n2230 VSS.n2229 292.5
R7302 VSS.n2547 VSS.n2230 292.5
R7303 VSS.n2557 VSS.n2556 292.5
R7304 VSS.n2558 VSS.n2557 292.5
R7305 VSS.n2219 VSS.n2215 292.5
R7306 VSS.n2221 VSS.n2219 292.5
R7307 VSS.n2602 VSS.n2601 292.5
R7308 VSS.n2603 VSS.n2602 292.5
R7309 VSS.n1461 VSS.n1460 292.5
R7310 VSS.n2604 VSS.n1461 292.5
R7311 VSS.n2607 VSS.n2606 292.5
R7312 VSS.n2606 VSS.n2605 292.5
R7313 VSS.n2608 VSS.n1459 292.5
R7314 VSS.n1459 VSS.n1458 292.5
R7315 VSS.n2610 VSS.n2609 292.5
R7316 VSS.n2611 VSS.n2610 292.5
R7317 VSS.n1457 VSS.n1456 292.5
R7318 VSS.n2612 VSS.n1457 292.5
R7319 VSS.n2615 VSS.n2614 292.5
R7320 VSS.n2614 VSS.n2613 292.5
R7321 VSS.n2616 VSS.n1455 292.5
R7322 VSS.n1455 VSS.n1454 292.5
R7323 VSS.n2619 VSS.n2618 292.5
R7324 VSS.n2620 VSS.n2619 292.5
R7325 VSS.n2617 VSS.n1453 292.5
R7326 VSS.n2621 VSS.n1453 292.5
R7327 VSS.n2623 VSS.n1452 292.5
R7328 VSS.n2623 VSS.n2622 292.5
R7329 VSS.n2625 VSS.n2624 292.5
R7330 VSS.n2624 VSS.n1447 292.5
R7331 VSS.n2074 VSS.n1562 292.5
R7332 VSS.n2075 VSS.n2074 292.5
R7333 VSS.n2073 VSS.n2072 292.5
R7334 VSS.n2073 VSS.n2042 292.5
R7335 VSS.n2071 VSS.n2043 292.5
R7336 VSS.n2046 VSS.n2043 292.5
R7337 VSS.n2070 VSS.n2069 292.5
R7338 VSS.n2069 VSS.n2068 292.5
R7339 VSS.n2045 VSS.n2044 292.5
R7340 VSS.n2067 VSS.n2045 292.5
R7341 VSS.n2065 VSS.n2064 292.5
R7342 VSS.n2066 VSS.n2065 292.5
R7343 VSS.n2063 VSS.n2048 292.5
R7344 VSS.n2048 VSS.n2047 292.5
R7345 VSS.n2062 VSS.n2061 292.5
R7346 VSS.n2061 VSS.n2060 292.5
R7347 VSS.n2050 VSS.n2049 292.5
R7348 VSS.n2059 VSS.n2050 292.5
R7349 VSS.n2057 VSS.n2056 292.5
R7350 VSS.n2058 VSS.n2057 292.5
R7351 VSS.n2055 VSS.n2054 292.5
R7352 VSS.n2054 VSS.n2051 292.5
R7353 VSS.n2053 VSS.n1464 292.5
R7354 VSS.n2053 VSS.n2052 292.5
R7355 VSS.n1482 VSS.n1481 292.5
R7356 VSS.n1481 VSS.n1480 292.5
R7357 VSS.n2206 VSS.n2205 292.5
R7358 VSS.n2207 VSS.n2206 292.5
R7359 VSS.n1493 VSS.n1491 292.5
R7360 VSS.n2196 VSS.n1493 292.5
R7361 VSS.n2187 VSS.n2186 292.5
R7362 VSS.n2186 VSS.n2185 292.5
R7363 VSS.n1502 VSS.n1501 292.5
R7364 VSS.n1501 VSS.n1500 292.5
R7365 VSS.n2171 VSS.n2170 292.5
R7366 VSS.n2172 VSS.n2171 292.5
R7367 VSS.n1514 VSS.n1512 292.5
R7368 VSS.n2162 VSS.n1514 292.5
R7369 VSS.n2153 VSS.n2152 292.5
R7370 VSS.n2152 VSS.n2151 292.5
R7371 VSS.n1523 VSS.n1522 292.5
R7372 VSS.n1522 VSS.n1521 292.5
R7373 VSS.n2137 VSS.n2136 292.5
R7374 VSS.n2138 VSS.n2137 292.5
R7375 VSS.n1535 VSS.n1533 292.5
R7376 VSS.n2127 VSS.n1535 292.5
R7377 VSS.n2118 VSS.n2117 292.5
R7378 VSS.n2117 VSS.n2116 292.5
R7379 VSS.n1546 VSS.n1544 292.5
R7380 VSS.n1544 VSS.n1543 292.5
R7381 VSS.n1796 VSS.n1795 292.5
R7382 VSS.n1797 VSS.n1796 292.5
R7383 VSS.n1779 VSS.n1777 292.5
R7384 VSS.n1781 VSS.n1779 292.5
R7385 VSS.n1771 VSS.n1770 292.5
R7386 VSS.n1809 VSS.n1771 292.5
R7387 VSS.n1819 VSS.n1818 292.5
R7388 VSS.n1820 VSS.n1819 292.5
R7389 VSS.n1760 VSS.n1758 292.5
R7390 VSS.n1762 VSS.n1760 292.5
R7391 VSS.n1752 VSS.n1751 292.5
R7392 VSS.n1831 VSS.n1752 292.5
R7393 VSS.n1841 VSS.n1840 292.5
R7394 VSS.n1842 VSS.n1841 292.5
R7395 VSS.n1741 VSS.n1739 292.5
R7396 VSS.n1743 VSS.n1741 292.5
R7397 VSS.n1733 VSS.n1732 292.5
R7398 VSS.n1854 VSS.n1733 292.5
R7399 VSS.n1864 VSS.n1863 292.5
R7400 VSS.n1865 VSS.n1864 292.5
R7401 VSS.n1719 VSS.n1717 292.5
R7402 VSS.n1724 VSS.n1719 292.5
R7403 VSS.n2021 VSS.n1575 292.5
R7404 VSS.n1575 VSS.n1574 292.5
R7405 VSS.n2023 VSS.n2022 292.5
R7406 VSS.n2024 VSS.n2023 292.5
R7407 VSS.n1573 VSS.n1572 292.5
R7408 VSS.n2025 VSS.n1573 292.5
R7409 VSS.n2028 VSS.n2027 292.5
R7410 VSS.n2027 VSS.n2026 292.5
R7411 VSS.n2029 VSS.n1571 292.5
R7412 VSS.n1571 VSS.n1570 292.5
R7413 VSS.n2031 VSS.n2030 292.5
R7414 VSS.n2032 VSS.n2031 292.5
R7415 VSS.n1569 VSS.n1568 292.5
R7416 VSS.n2033 VSS.n1569 292.5
R7417 VSS.n2036 VSS.n2035 292.5
R7418 VSS.n2035 VSS.n2034 292.5
R7419 VSS.n2037 VSS.n1567 292.5
R7420 VSS.n1567 VSS.n1566 292.5
R7421 VSS.n2039 VSS.n2038 292.5
R7422 VSS.n2040 VSS.n2039 292.5
R7423 VSS.n1564 VSS.n1563 292.5
R7424 VSS.n2041 VSS.n1564 292.5
R7425 VSS.n2079 VSS.n2078 292.5
R7426 VSS.n2078 VSS.n2077 292.5
R7427 VSS.n1994 VSS.n1590 292.5
R7428 VSS.n1590 VSS.n1589 292.5
R7429 VSS.n1996 VSS.n1995 292.5
R7430 VSS.n1997 VSS.n1996 292.5
R7431 VSS.n1588 VSS.n1587 292.5
R7432 VSS.n1998 VSS.n1588 292.5
R7433 VSS.n2001 VSS.n2000 292.5
R7434 VSS.n2000 VSS.n1999 292.5
R7435 VSS.n2002 VSS.n1586 292.5
R7436 VSS.n1586 VSS.n1585 292.5
R7437 VSS.n2004 VSS.n2003 292.5
R7438 VSS.n2005 VSS.n2004 292.5
R7439 VSS.n1584 VSS.n1583 292.5
R7440 VSS.n2006 VSS.n1584 292.5
R7441 VSS.n2010 VSS.n2009 292.5
R7442 VSS.n2009 VSS.n2008 292.5
R7443 VSS.n2011 VSS.n1582 292.5
R7444 VSS.n2007 VSS.n1582 292.5
R7445 VSS.n2013 VSS.n2012 292.5
R7446 VSS.n2013 VSS.n1581 292.5
R7447 VSS.n2014 VSS.n1576 292.5
R7448 VSS.n2015 VSS.n2014 292.5
R7449 VSS.n1993 VSS.n1992 292.5
R7450 VSS.n1992 VSS.n1991 292.5
R7451 VSS.n1678 VSS.n1677 292.5
R7452 VSS.n1878 VSS.n1678 292.5
R7453 VSS.n1888 VSS.n1887 292.5
R7454 VSS.n1889 VSS.n1888 292.5
R7455 VSS.n1667 VSS.n1665 292.5
R7456 VSS.n1669 VSS.n1667 292.5
R7457 VSS.n1659 VSS.n1658 292.5
R7458 VSS.n1901 VSS.n1659 292.5
R7459 VSS.n1911 VSS.n1910 292.5
R7460 VSS.n1912 VSS.n1911 292.5
R7461 VSS.n1648 VSS.n1646 292.5
R7462 VSS.n1650 VSS.n1648 292.5
R7463 VSS.n1640 VSS.n1639 292.5
R7464 VSS.n1923 VSS.n1640 292.5
R7465 VSS.n1933 VSS.n1932 292.5
R7466 VSS.n1934 VSS.n1933 292.5
R7467 VSS.n1629 VSS.n1627 292.5
R7468 VSS.n1631 VSS.n1629 292.5
R7469 VSS.n1621 VSS.n1620 292.5
R7470 VSS.n1946 VSS.n1621 292.5
R7471 VSS.n1956 VSS.n1955 292.5
R7472 VSS.n1957 VSS.n1956 292.5
R7473 VSS.n1962 VSS.n1607 292.5
R7474 VSS.n1607 VSS.n1606 292.5
R7475 VSS.n1605 VSS.n1603 292.5
R7476 VSS.n15794 VSS.n15679 287.581
R7477 VSS.n15792 VSS.n15680 287.581
R7478 VSS.n15781 VSS.n15780 287.581
R7479 VSS.n15771 VSS.n15698 287.581
R7480 VSS.n15769 VSS.n15699 287.581
R7481 VSS.n15758 VSS.n15757 287.581
R7482 VSS.n15749 VSS.n15717 287.581
R7483 VSS.n15747 VSS.n15718 287.581
R7484 VSS.n15736 VSS.n15735 287.581
R7485 VSS.n16019 VSS.n14001 287.581
R7486 VSS.n16017 VSS.n14002 287.581
R7487 VSS.n16006 VSS.n16005 287.581
R7488 VSS.n15886 VSS.n15567 287.581
R7489 VSS.n15884 VSS.n15568 287.581
R7490 VSS.n15873 VSS.n15872 287.581
R7491 VSS.n15863 VSS.n15586 287.581
R7492 VSS.n15861 VSS.n15587 287.581
R7493 VSS.n15850 VSS.n15849 287.581
R7494 VSS.n15841 VSS.n15605 287.581
R7495 VSS.n15839 VSS.n15606 287.581
R7496 VSS.n15828 VSS.n15827 287.581
R7497 VSS.n15818 VSS.n15624 287.581
R7498 VSS.n15816 VSS.n15625 287.581
R7499 VSS.n15805 VSS.n15804 287.581
R7500 VSS.n15804 VSS.n15634 287.581
R7501 VSS.n15461 VSS.n15460 287.581
R7502 VSS.n15471 VSS.n14124 287.581
R7503 VSS.n15473 VSS.n14118 287.581
R7504 VSS.n15485 VSS.n15484 287.581
R7505 VSS.n15496 VSS.n15495 287.581
R7506 VSS.n15506 VSS.n14103 287.581
R7507 VSS.n15508 VSS.n14097 287.581
R7508 VSS.n15519 VSS.n15518 287.581
R7509 VSS.n15530 VSS.n15529 287.581
R7510 VSS.n15540 VSS.n14082 287.581
R7511 VSS.n15542 VSS.n14076 287.581
R7512 VSS.n15554 VSS.n15553 287.581
R7513 VSS.n15554 VSS.n14069 287.581
R7514 VSS.n15227 VSS.n15092 287.581
R7515 VSS.n15225 VSS.n15093 287.581
R7516 VSS.n15214 VSS.n15213 287.581
R7517 VSS.n15204 VSS.n15111 287.581
R7518 VSS.n15202 VSS.n15112 287.581
R7519 VSS.n15191 VSS.n15190 287.581
R7520 VSS.n15182 VSS.n15130 287.581
R7521 VSS.n15180 VSS.n15131 287.581
R7522 VSS.n15169 VSS.n15168 287.581
R7523 VSS.n15159 VSS.n15149 287.581
R7524 VSS.n15157 VSS.n14143 287.581
R7525 VSS.n15444 VSS.n15443 287.581
R7526 VSS.n15443 VSS.n14144 287.581
R7527 VSS.n15319 VSS.n14980 287.581
R7528 VSS.n15317 VSS.n14981 287.581
R7529 VSS.n15306 VSS.n15305 287.581
R7530 VSS.n15296 VSS.n14999 287.581
R7531 VSS.n15294 VSS.n15000 287.581
R7532 VSS.n15283 VSS.n15282 287.581
R7533 VSS.n15274 VSS.n15018 287.581
R7534 VSS.n15272 VSS.n15019 287.581
R7535 VSS.n15261 VSS.n15260 287.581
R7536 VSS.n15251 VSS.n15037 287.581
R7537 VSS.n15249 VSS.n15038 287.581
R7538 VSS.n15238 VSS.n15237 287.581
R7539 VSS.n15237 VSS.n15047 287.581
R7540 VSS.n14875 VSS.n14295 287.581
R7541 VSS.n14887 VSS.n14886 287.581
R7542 VSS.n14898 VSS.n14897 287.581
R7543 VSS.n14908 VSS.n14280 287.581
R7544 VSS.n14910 VSS.n14274 287.581
R7545 VSS.n14922 VSS.n14921 287.581
R7546 VSS.n14932 VSS.n14931 287.581
R7547 VSS.n14942 VSS.n14259 287.581
R7548 VSS.n14944 VSS.n14253 287.581
R7549 VSS.n14956 VSS.n14955 287.581
R7550 VSS.n14967 VSS.n14966 287.581
R7551 VSS.n15330 VSS.n14239 287.581
R7552 VSS.n15331 VSS.n15330 287.581
R7553 VSS.n14626 VSS.n14483 287.581
R7554 VSS.n14624 VSS.n14484 287.581
R7555 VSS.n14613 VSS.n14612 287.581
R7556 VSS.n14603 VSS.n14502 287.581
R7557 VSS.n14601 VSS.n14503 287.581
R7558 VSS.n14590 VSS.n14589 287.581
R7559 VSS.n14581 VSS.n14521 287.581
R7560 VSS.n14579 VSS.n14522 287.581
R7561 VSS.n14568 VSS.n14567 287.581
R7562 VSS.n14558 VSS.n14540 287.581
R7563 VSS.n14556 VSS.n14541 287.581
R7564 VSS.n14872 VSS.n14302 287.581
R7565 VSS.n14873 VSS.n14872 287.581
R7566 VSS.n14718 VSS.n14365 287.581
R7567 VSS.n14716 VSS.n14371 287.581
R7568 VSS.n14705 VSS.n14704 287.581
R7569 VSS.n14695 VSS.n14390 287.581
R7570 VSS.n14693 VSS.n14391 287.581
R7571 VSS.n14682 VSS.n14681 287.581
R7572 VSS.n14673 VSS.n14409 287.581
R7573 VSS.n14671 VSS.n14410 287.581
R7574 VSS.n14660 VSS.n14659 287.581
R7575 VSS.n14650 VSS.n14428 287.581
R7576 VSS.n14648 VSS.n14429 287.581
R7577 VSS.n14637 VSS.n14636 287.581
R7578 VSS.n14636 VSS.n14438 287.581
R7579 VSS.n12302 VSS.n11993 287.581
R7580 VSS.n12300 VSS.n11994 287.581
R7581 VSS.n12289 VSS.n12288 287.581
R7582 VSS.n12279 VSS.n12012 287.581
R7583 VSS.n12277 VSS.n12013 287.581
R7584 VSS.n12266 VSS.n12265 287.581
R7585 VSS.n12257 VSS.n12031 287.581
R7586 VSS.n12255 VSS.n12032 287.581
R7587 VSS.n12244 VSS.n12243 287.581
R7588 VSS.n12234 VSS.n12050 287.581
R7589 VSS.n12232 VSS.n12051 287.581
R7590 VSS.n12221 VSS.n12220 287.581
R7591 VSS.n12394 VSS.n11914 287.581
R7592 VSS.n12392 VSS.n11915 287.581
R7593 VSS.n12381 VSS.n12380 287.581
R7594 VSS.n12371 VSS.n11933 287.581
R7595 VSS.n12369 VSS.n11934 287.581
R7596 VSS.n12358 VSS.n12357 287.581
R7597 VSS.n12349 VSS.n11952 287.581
R7598 VSS.n12347 VSS.n11953 287.581
R7599 VSS.n12336 VSS.n12335 287.581
R7600 VSS.n12326 VSS.n11971 287.581
R7601 VSS.n12324 VSS.n11972 287.581
R7602 VSS.n12313 VSS.n12312 287.581
R7603 VSS.n12312 VSS.n11981 287.581
R7604 VSS.n11809 VSS.n11600 287.581
R7605 VSS.n11821 VSS.n11820 287.581
R7606 VSS.n11832 VSS.n11831 287.581
R7607 VSS.n11842 VSS.n11585 287.581
R7608 VSS.n11844 VSS.n11579 287.581
R7609 VSS.n11856 VSS.n11855 287.581
R7610 VSS.n11866 VSS.n11865 287.581
R7611 VSS.n11876 VSS.n11564 287.581
R7612 VSS.n11878 VSS.n11558 287.581
R7613 VSS.n11890 VSS.n11889 287.581
R7614 VSS.n11901 VSS.n11900 287.581
R7615 VSS.n12405 VSS.n11544 287.581
R7616 VSS.n12406 VSS.n12405 287.581
R7617 VSS.n11675 VSS.n11674 287.581
R7618 VSS.n11686 VSS.n11685 287.581
R7619 VSS.n11696 VSS.n11657 287.581
R7620 VSS.n11698 VSS.n11651 287.581
R7621 VSS.n11710 VSS.n11709 287.581
R7622 VSS.n11721 VSS.n11720 287.581
R7623 VSS.n11730 VSS.n11636 287.581
R7624 VSS.n11732 VSS.n11630 287.581
R7625 VSS.n11744 VSS.n11743 287.581
R7626 VSS.n11755 VSS.n11754 287.581
R7627 VSS.n11765 VSS.n11614 287.581
R7628 VSS.n11767 VSS.n11606 287.581
R7629 VSS.n11807 VSS.n11606 287.581
R7630 VSS.n13255 VSS.n13249 287.581
R7631 VSS.n13293 VSS.n13292 287.581
R7632 VSS.n13283 VSS.n13265 287.581
R7633 VSS.n13281 VSS.n13266 287.581
R7634 VSS.n13453 VSS.n11435 287.581
R7635 VSS.n13451 VSS.n11436 287.581
R7636 VSS.n13440 VSS.n13439 287.581
R7637 VSS.n13431 VSS.n11454 287.581
R7638 VSS.n13429 VSS.n11455 287.581
R7639 VSS.n13418 VSS.n13417 287.581
R7640 VSS.n13408 VSS.n11473 287.581
R7641 VSS.n13406 VSS.n11474 287.581
R7642 VSS.n11485 VSS.n11474 287.581
R7643 VSS.n13154 VSS.n13153 287.581
R7644 VSS.n13165 VSS.n13164 287.581
R7645 VSS.n13175 VSS.n12566 287.581
R7646 VSS.n13177 VSS.n12560 287.581
R7647 VSS.n13189 VSS.n13188 287.581
R7648 VSS.n13200 VSS.n13199 287.581
R7649 VSS.n13209 VSS.n12545 287.581
R7650 VSS.n13211 VSS.n12539 287.581
R7651 VSS.n13223 VSS.n13222 287.581
R7652 VSS.n13234 VSS.n13233 287.581
R7653 VSS.n13235 VSS.n12524 287.581
R7654 VSS.n13307 VSS.n13248 287.581
R7655 VSS.n13307 VSS.n13306 287.581
R7656 VSS.n12898 VSS.n12892 287.581
R7657 VSS.n13044 VSS.n13043 287.581
R7658 VSS.n13034 VSS.n12908 287.581
R7659 VSS.n13032 VSS.n12909 287.581
R7660 VSS.n13021 VSS.n13020 287.581
R7661 VSS.n13011 VSS.n12927 287.581
R7662 VSS.n13009 VSS.n12928 287.581
R7663 VSS.n12999 VSS.n12998 287.581
R7664 VSS.n12989 VSS.n12946 287.581
R7665 VSS.n12987 VSS.n12947 287.581
R7666 VSS.n12976 VSS.n12975 287.581
R7667 VSS.n12966 VSS.n12965 287.581
R7668 VSS.n12966 VSS.n12581 287.581
R7669 VSS.n12797 VSS.n12796 287.581
R7670 VSS.n12808 VSS.n12807 287.581
R7671 VSS.n12818 VSS.n12707 287.581
R7672 VSS.n12820 VSS.n12701 287.581
R7673 VSS.n12832 VSS.n12831 287.581
R7674 VSS.n12843 VSS.n12842 287.581
R7675 VSS.n12852 VSS.n12686 287.581
R7676 VSS.n12854 VSS.n12680 287.581
R7677 VSS.n12866 VSS.n12865 287.581
R7678 VSS.n12877 VSS.n12876 287.581
R7679 VSS.n12878 VSS.n12665 287.581
R7680 VSS.n13058 VSS.n12891 287.581
R7681 VSS.n13058 VSS.n13057 287.581
R7682 VSS.n7077 VSS.n7076 287.581
R7683 VSS.n7087 VSS.n7059 287.581
R7684 VSS.n7089 VSS.n7053 287.581
R7685 VSS.n7101 VSS.n7100 287.581
R7686 VSS.n7112 VSS.n7111 287.581
R7687 VSS.n7122 VSS.n7038 287.581
R7688 VSS.n7124 VSS.n7032 287.581
R7689 VSS.n7135 VSS.n7134 287.581
R7690 VSS.n7146 VSS.n7145 287.581
R7691 VSS.n7156 VSS.n7017 287.581
R7692 VSS.n7158 VSS.n7011 287.581
R7693 VSS.n7171 VSS.n7169 287.581
R7694 VSS.n8760 VSS.n8759 287.581
R7695 VSS.n8752 VSS.n8737 287.581
R7696 VSS.n8925 VSS.n6907 287.581
R7697 VSS.n8923 VSS.n6908 287.581
R7698 VSS.n8912 VSS.n8911 287.581
R7699 VSS.n8902 VSS.n6926 287.581
R7700 VSS.n8900 VSS.n6927 287.581
R7701 VSS.n8890 VSS.n8889 287.581
R7702 VSS.n8880 VSS.n6945 287.581
R7703 VSS.n8878 VSS.n6946 287.581
R7704 VSS.n8867 VSS.n8866 287.581
R7705 VSS.n8857 VSS.n6964 287.581
R7706 VSS.n8857 VSS.n8856 287.581
R7707 VSS.n8636 VSS.n7314 287.581
R7708 VSS.n8648 VSS.n8647 287.581
R7709 VSS.n8659 VSS.n8658 287.581
R7710 VSS.n8669 VSS.n7299 287.581
R7711 VSS.n8671 VSS.n7293 287.581
R7712 VSS.n8683 VSS.n8682 287.581
R7713 VSS.n8693 VSS.n8692 287.581
R7714 VSS.n8703 VSS.n7278 287.581
R7715 VSS.n8705 VSS.n7272 287.581
R7716 VSS.n8717 VSS.n8716 287.581
R7717 VSS.n8728 VSS.n8727 287.581
R7718 VSS.n8771 VSS.n7257 287.581
R7719 VSS.n8772 VSS.n8771 287.581
R7720 VSS.n8538 VSS.n8537 287.581
R7721 VSS.n8530 VSS.n8379 287.581
R7722 VSS.n8528 VSS.n8390 287.581
R7723 VSS.n8517 VSS.n8516 287.581
R7724 VSS.n8507 VSS.n8409 287.581
R7725 VSS.n8505 VSS.n8410 287.581
R7726 VSS.n8494 VSS.n8493 287.581
R7727 VSS.n8485 VSS.n8428 287.581
R7728 VSS.n8483 VSS.n8429 287.581
R7729 VSS.n8472 VSS.n8471 287.581
R7730 VSS.n8462 VSS.n8447 287.581
R7731 VSS.n8460 VSS.n7320 287.581
R7732 VSS.n8634 VSS.n7320 287.581
R7733 VSS.n8278 VSS.n7454 287.581
R7734 VSS.n8290 VSS.n8289 287.581
R7735 VSS.n8301 VSS.n8300 287.581
R7736 VSS.n8311 VSS.n7439 287.581
R7737 VSS.n8313 VSS.n7433 287.581
R7738 VSS.n8325 VSS.n8324 287.581
R7739 VSS.n8335 VSS.n8334 287.581
R7740 VSS.n8345 VSS.n7418 287.581
R7741 VSS.n8347 VSS.n7412 287.581
R7742 VSS.n8359 VSS.n8358 287.581
R7743 VSS.n8370 VSS.n8369 287.581
R7744 VSS.n8549 VSS.n7397 287.581
R7745 VSS.n8550 VSS.n8549 287.581
R7746 VSS.n8180 VSS.n8179 287.581
R7747 VSS.n8172 VSS.n8021 287.581
R7748 VSS.n8170 VSS.n8032 287.581
R7749 VSS.n8159 VSS.n8158 287.581
R7750 VSS.n8149 VSS.n8051 287.581
R7751 VSS.n8147 VSS.n8052 287.581
R7752 VSS.n8136 VSS.n8135 287.581
R7753 VSS.n8127 VSS.n8070 287.581
R7754 VSS.n8125 VSS.n8071 287.581
R7755 VSS.n8114 VSS.n8113 287.581
R7756 VSS.n8104 VSS.n8089 287.581
R7757 VSS.n8102 VSS.n7460 287.581
R7758 VSS.n8276 VSS.n7460 287.581
R7759 VSS.n7920 VSS.n7594 287.581
R7760 VSS.n7932 VSS.n7931 287.581
R7761 VSS.n7943 VSS.n7942 287.581
R7762 VSS.n7953 VSS.n7579 287.581
R7763 VSS.n7955 VSS.n7573 287.581
R7764 VSS.n7967 VSS.n7966 287.581
R7765 VSS.n7977 VSS.n7976 287.581
R7766 VSS.n7987 VSS.n7558 287.581
R7767 VSS.n7989 VSS.n7552 287.581
R7768 VSS.n8001 VSS.n8000 287.581
R7769 VSS.n8012 VSS.n8011 287.581
R7770 VSS.n8191 VSS.n7537 287.581
R7771 VSS.n8192 VSS.n8191 287.581
R7772 VSS.n7832 VSS.n7673 287.581
R7773 VSS.n7830 VSS.n7678 287.581
R7774 VSS.n7819 VSS.n7818 287.581
R7775 VSS.n7809 VSS.n7697 287.581
R7776 VSS.n7807 VSS.n7698 287.581
R7777 VSS.n7796 VSS.n7795 287.581
R7778 VSS.n7787 VSS.n7716 287.581
R7779 VSS.n7785 VSS.n7717 287.581
R7780 VSS.n7774 VSS.n7773 287.581
R7781 VSS.n7764 VSS.n7735 287.581
R7782 VSS.n7762 VSS.n7736 287.581
R7783 VSS.n7751 VSS.n7600 287.581
R7784 VSS.n7918 VSS.n7600 287.581
R7785 VSS.n5422 VSS.n5416 287.581
R7786 VSS.n5557 VSS.n5556 287.581
R7787 VSS.n5547 VSS.n5432 287.581
R7788 VSS.n5545 VSS.n5433 287.581
R7789 VSS.n5534 VSS.n5533 287.581
R7790 VSS.n5524 VSS.n5451 287.581
R7791 VSS.n5522 VSS.n5452 287.581
R7792 VSS.n5512 VSS.n5511 287.581
R7793 VSS.n5502 VSS.n5470 287.581
R7794 VSS.n5500 VSS.n5471 287.581
R7795 VSS.n5489 VSS.n5488 287.581
R7796 VSS.n5659 VSS.n3641 287.581
R7797 VSS.n5321 VSS.n5320 287.581
R7798 VSS.n5332 VSS.n5331 287.581
R7799 VSS.n5342 VSS.n3737 287.581
R7800 VSS.n5344 VSS.n3731 287.581
R7801 VSS.n5356 VSS.n5355 287.581
R7802 VSS.n5367 VSS.n5366 287.581
R7803 VSS.n5376 VSS.n3716 287.581
R7804 VSS.n5378 VSS.n3710 287.581
R7805 VSS.n5390 VSS.n5389 287.581
R7806 VSS.n5401 VSS.n5400 287.581
R7807 VSS.n5402 VSS.n3695 287.581
R7808 VSS.n5571 VSS.n5415 287.581
R7809 VSS.n5571 VSS.n5570 287.581
R7810 VSS.n5065 VSS.n5059 287.581
R7811 VSS.n5211 VSS.n5210 287.581
R7812 VSS.n5201 VSS.n5075 287.581
R7813 VSS.n5199 VSS.n5076 287.581
R7814 VSS.n5188 VSS.n5187 287.581
R7815 VSS.n5178 VSS.n5094 287.581
R7816 VSS.n5176 VSS.n5095 287.581
R7817 VSS.n5166 VSS.n5165 287.581
R7818 VSS.n5156 VSS.n5113 287.581
R7819 VSS.n5154 VSS.n5114 287.581
R7820 VSS.n5143 VSS.n5142 287.581
R7821 VSS.n5133 VSS.n5132 287.581
R7822 VSS.n5133 VSS.n3752 287.581
R7823 VSS.n4964 VSS.n4963 287.581
R7824 VSS.n4975 VSS.n4974 287.581
R7825 VSS.n4985 VSS.n3878 287.581
R7826 VSS.n4987 VSS.n3872 287.581
R7827 VSS.n4999 VSS.n4998 287.581
R7828 VSS.n5010 VSS.n5009 287.581
R7829 VSS.n5019 VSS.n3857 287.581
R7830 VSS.n5021 VSS.n3851 287.581
R7831 VSS.n5033 VSS.n5032 287.581
R7832 VSS.n5044 VSS.n5043 287.581
R7833 VSS.n5045 VSS.n3836 287.581
R7834 VSS.n5225 VSS.n5058 287.581
R7835 VSS.n5225 VSS.n5224 287.581
R7836 VSS.n4708 VSS.n4702 287.581
R7837 VSS.n4854 VSS.n4853 287.581
R7838 VSS.n4844 VSS.n4718 287.581
R7839 VSS.n4842 VSS.n4719 287.581
R7840 VSS.n4831 VSS.n4830 287.581
R7841 VSS.n4821 VSS.n4737 287.581
R7842 VSS.n4819 VSS.n4738 287.581
R7843 VSS.n4809 VSS.n4808 287.581
R7844 VSS.n4799 VSS.n4756 287.581
R7845 VSS.n4797 VSS.n4757 287.581
R7846 VSS.n4786 VSS.n4785 287.581
R7847 VSS.n4776 VSS.n4775 287.581
R7848 VSS.n4776 VSS.n3893 287.581
R7849 VSS.n4607 VSS.n4606 287.581
R7850 VSS.n4618 VSS.n4617 287.581
R7851 VSS.n4628 VSS.n4019 287.581
R7852 VSS.n4630 VSS.n4013 287.581
R7853 VSS.n4642 VSS.n4641 287.581
R7854 VSS.n4653 VSS.n4652 287.581
R7855 VSS.n4662 VSS.n3998 287.581
R7856 VSS.n4664 VSS.n3992 287.581
R7857 VSS.n4676 VSS.n4675 287.581
R7858 VSS.n4687 VSS.n4686 287.581
R7859 VSS.n4688 VSS.n3977 287.581
R7860 VSS.n4868 VSS.n4701 287.581
R7861 VSS.n4868 VSS.n4867 287.581
R7862 VSS.n4351 VSS.n4345 287.581
R7863 VSS.n4497 VSS.n4496 287.581
R7864 VSS.n4487 VSS.n4361 287.581
R7865 VSS.n4485 VSS.n4362 287.581
R7866 VSS.n4474 VSS.n4473 287.581
R7867 VSS.n4464 VSS.n4380 287.581
R7868 VSS.n4462 VSS.n4381 287.581
R7869 VSS.n4452 VSS.n4451 287.581
R7870 VSS.n4442 VSS.n4399 287.581
R7871 VSS.n4440 VSS.n4400 287.581
R7872 VSS.n4429 VSS.n4428 287.581
R7873 VSS.n4419 VSS.n4418 287.581
R7874 VSS.n4419 VSS.n4034 287.581
R7875 VSS.n4250 VSS.n4249 287.581
R7876 VSS.n4261 VSS.n4260 287.581
R7877 VSS.n4271 VSS.n4160 287.581
R7878 VSS.n4273 VSS.n4154 287.581
R7879 VSS.n4285 VSS.n4284 287.581
R7880 VSS.n4296 VSS.n4295 287.581
R7881 VSS.n4305 VSS.n4139 287.581
R7882 VSS.n4307 VSS.n4133 287.581
R7883 VSS.n4319 VSS.n4318 287.581
R7884 VSS.n4330 VSS.n4329 287.581
R7885 VSS.n4331 VSS.n4118 287.581
R7886 VSS.n4511 VSS.n4344 287.581
R7887 VSS.n4511 VSS.n4510 287.581
R7888 VSS.n2960 VSS.n2808 287.581
R7889 VSS.n2958 VSS.n2809 287.581
R7890 VSS.n2947 VSS.n2946 287.581
R7891 VSS.n2937 VSS.n2827 287.581
R7892 VSS.n2935 VSS.n2828 287.581
R7893 VSS.n2924 VSS.n2923 287.581
R7894 VSS.n2915 VSS.n2846 287.581
R7895 VSS.n2913 VSS.n2847 287.581
R7896 VSS.n2902 VSS.n2901 287.581
R7897 VSS.n2892 VSS.n2865 287.581
R7898 VSS.n2890 VSS.n2866 287.581
R7899 VSS.n2879 VSS.n1272 287.581
R7900 VSS.n2702 VSS.n2701 287.581
R7901 VSS.n2712 VSS.n1365 287.581
R7902 VSS.n2714 VSS.n1359 287.581
R7903 VSS.n2726 VSS.n2725 287.581
R7904 VSS.n2737 VSS.n2736 287.581
R7905 VSS.n2747 VSS.n1344 287.581
R7906 VSS.n2749 VSS.n1338 287.581
R7907 VSS.n2760 VSS.n2759 287.581
R7908 VSS.n2771 VSS.n2770 287.581
R7909 VSS.n2781 VSS.n1323 287.581
R7910 VSS.n2783 VSS.n1317 287.581
R7911 VSS.n2795 VSS.n2794 287.581
R7912 VSS.n2795 VSS.n1310 287.581
R7913 VSS.n2468 VSS.n2333 287.581
R7914 VSS.n2466 VSS.n2334 287.581
R7915 VSS.n2455 VSS.n2454 287.581
R7916 VSS.n2445 VSS.n2352 287.581
R7917 VSS.n2443 VSS.n2353 287.581
R7918 VSS.n2432 VSS.n2431 287.581
R7919 VSS.n2423 VSS.n2371 287.581
R7920 VSS.n2421 VSS.n2372 287.581
R7921 VSS.n2410 VSS.n2409 287.581
R7922 VSS.n2400 VSS.n2390 287.581
R7923 VSS.n2398 VSS.n1384 287.581
R7924 VSS.n2685 VSS.n2684 287.581
R7925 VSS.n2684 VSS.n1385 287.581
R7926 VSS.n2560 VSS.n2221 287.581
R7927 VSS.n2558 VSS.n2222 287.581
R7928 VSS.n2547 VSS.n2546 287.581
R7929 VSS.n2537 VSS.n2240 287.581
R7930 VSS.n2535 VSS.n2241 287.581
R7931 VSS.n2524 VSS.n2523 287.581
R7932 VSS.n2515 VSS.n2259 287.581
R7933 VSS.n2513 VSS.n2260 287.581
R7934 VSS.n2502 VSS.n2501 287.581
R7935 VSS.n2492 VSS.n2278 287.581
R7936 VSS.n2490 VSS.n2279 287.581
R7937 VSS.n2479 VSS.n2478 287.581
R7938 VSS.n2478 VSS.n2288 287.581
R7939 VSS.n2116 VSS.n1536 287.581
R7940 VSS.n2128 VSS.n2127 287.581
R7941 VSS.n2139 VSS.n2138 287.581
R7942 VSS.n2149 VSS.n1521 287.581
R7943 VSS.n2151 VSS.n1515 287.581
R7944 VSS.n2163 VSS.n2162 287.581
R7945 VSS.n2173 VSS.n2172 287.581
R7946 VSS.n2183 VSS.n1500 287.581
R7947 VSS.n2185 VSS.n1494 287.581
R7948 VSS.n2197 VSS.n2196 287.581
R7949 VSS.n2208 VSS.n2207 287.581
R7950 VSS.n2571 VSS.n1480 287.581
R7951 VSS.n2572 VSS.n2571 287.581
R7952 VSS.n1867 VSS.n1724 287.581
R7953 VSS.n1865 VSS.n1725 287.581
R7954 VSS.n1854 VSS.n1853 287.581
R7955 VSS.n1844 VSS.n1743 287.581
R7956 VSS.n1842 VSS.n1744 287.581
R7957 VSS.n1831 VSS.n1830 287.581
R7958 VSS.n1822 VSS.n1762 287.581
R7959 VSS.n1820 VSS.n1763 287.581
R7960 VSS.n1809 VSS.n1808 287.581
R7961 VSS.n1799 VSS.n1781 287.581
R7962 VSS.n1797 VSS.n1782 287.581
R7963 VSS.n2113 VSS.n1543 287.581
R7964 VSS.n2114 VSS.n2113 287.581
R7965 VSS.n1959 VSS.n1606 287.581
R7966 VSS.n1957 VSS.n1612 287.581
R7967 VSS.n1946 VSS.n1945 287.581
R7968 VSS.n1936 VSS.n1631 287.581
R7969 VSS.n1934 VSS.n1632 287.581
R7970 VSS.n1923 VSS.n1922 287.581
R7971 VSS.n1914 VSS.n1650 287.581
R7972 VSS.n1912 VSS.n1651 287.581
R7973 VSS.n1901 VSS.n1900 287.581
R7974 VSS.n1891 VSS.n1669 287.581
R7975 VSS.n1889 VSS.n1670 287.581
R7976 VSS.n1878 VSS.n1877 287.581
R7977 VSS.n1877 VSS.n1679 287.581
R7978 VSS.n17350 VSS.n17321 258.333
R7979 VSS.n16106 VSS.n16065 258.333
R7980 VSS.n16196 VSS.n16155 258.333
R7981 VSS.n16286 VSS.n16245 258.333
R7982 VSS.n16376 VSS.n16335 258.333
R7983 VSS.n16466 VSS.n16425 258.333
R7984 VSS.n16556 VSS.n16515 258.333
R7985 VSS.n16646 VSS.n16605 258.333
R7986 VSS.n11113 VSS.n11072 258.333
R7987 VSS.n11023 VSS.n10982 258.333
R7988 VSS.n10933 VSS.n10892 258.333
R7989 VSS.n10843 VSS.n10802 258.333
R7990 VSS.n10753 VSS.n10712 258.333
R7991 VSS.n10663 VSS.n10622 258.333
R7992 VSS.n10573 VSS.n10532 258.333
R7993 VSS.n13850 VSS.n13818 258.333
R7994 VSS.n9241 VSS.n9200 258.333
R7995 VSS.n9331 VSS.n9290 258.333
R7996 VSS.n9421 VSS.n9380 258.333
R7997 VSS.n9511 VSS.n9470 258.333
R7998 VSS.n9601 VSS.n9560 258.333
R7999 VSS.n9691 VSS.n9650 258.333
R8000 VSS.n6726 VSS.n6725 258.333
R8001 VSS.n5698 VSS.n5678 258.333
R8002 VSS.n5820 VSS.n5800 258.333
R8003 VSS.n5942 VSS.n5922 258.333
R8004 VSS.n6064 VSS.n6044 258.333
R8005 VSS.n6186 VSS.n6166 258.333
R8006 VSS.n6308 VSS.n6288 258.333
R8007 VSS.n6430 VSS.n6410 258.333
R8008 VSS.n6573 VSS.n6525 258.333
R8009 VSS.n59 VSS.n17 258.333
R8010 VSS.n149 VSS.n108 258.333
R8011 VSS.n239 VSS.n198 258.333
R8012 VSS.n329 VSS.n288 258.333
R8013 VSS.n419 VSS.n378 258.333
R8014 VSS.n509 VSS.n468 258.333
R8015 VSS.n599 VSS.n558 258.333
R8016 VSS.n14751 VSS.n14351 257.464
R8017 VSS.n12767 VSS.n12737 257.464
R8018 VSS.n7864 VSS.n7658 257.464
R8019 VSS.n6854 VSS.n6745 257.464
R8020 VSS.n4220 VSS.n4190 257.464
R8021 VSS.n1992 VSS.n1592 257.464
R8022 VSS.n15972 VSS.n14026 251.613
R8023 VSS.n12187 VSS.n12075 251.613
R8024 VSS.n7201 VSS.n6992 251.613
R8025 VSS.n6878 VSS.n6732 251.613
R8026 VSS.n5632 VSS.n3658 251.613
R8027 VSS.n3019 VSS.n1284 251.613
R8028 VSS.n17369 VSS.n17368 249.999
R8029 VSS.n16125 VSS.n16124 249.999
R8030 VSS.n16215 VSS.n16214 249.999
R8031 VSS.n16305 VSS.n16304 249.999
R8032 VSS.n16395 VSS.n16394 249.999
R8033 VSS.n16485 VSS.n16484 249.999
R8034 VSS.n16575 VSS.n16574 249.999
R8035 VSS.n16665 VSS.n16664 249.999
R8036 VSS.n11132 VSS.n11131 249.999
R8037 VSS.n11042 VSS.n11041 249.999
R8038 VSS.n10952 VSS.n10951 249.999
R8039 VSS.n10862 VSS.n10861 249.999
R8040 VSS.n10772 VSS.n10771 249.999
R8041 VSS.n10682 VSS.n10681 249.999
R8042 VSS.n10592 VSS.n10591 249.999
R8043 VSS.n13869 VSS.n13868 249.999
R8044 VSS.n9113 VSS.n8993 249.999
R8045 VSS.n9260 VSS.n9259 249.999
R8046 VSS.n9350 VSS.n9349 249.999
R8047 VSS.n9440 VSS.n9439 249.999
R8048 VSS.n9530 VSS.n9529 249.999
R8049 VSS.n9620 VSS.n9619 249.999
R8050 VSS.n9710 VSS.n9709 249.999
R8051 VSS.n10297 VSS.n9165 249.999
R8052 VSS.n5717 VSS.n5716 249.999
R8053 VSS.n5839 VSS.n5838 249.999
R8054 VSS.n5961 VSS.n5960 249.999
R8055 VSS.n6083 VSS.n6082 249.999
R8056 VSS.n6205 VSS.n6204 249.999
R8057 VSS.n6327 VSS.n6326 249.999
R8058 VSS.n6449 VSS.n6448 249.999
R8059 VSS.n6558 VSS.n6556 249.999
R8060 VSS.n78 VSS.n77 249.999
R8061 VSS.n168 VSS.n167 249.999
R8062 VSS.n258 VSS.n257 249.999
R8063 VSS.n348 VSS.n347 249.999
R8064 VSS.n438 VSS.n437 249.999
R8065 VSS.n528 VSS.n527 249.999
R8066 VSS.n618 VSS.n617 249.999
R8067 VSS.n6710 VSS.n6709 221.666
R8068 VSS.n17461 VSS.n16030 205
R8069 VSS.n17307 VSS.n16055 205
R8070 VSS.n17217 VSS.n16145 205
R8071 VSS.n17127 VSS.n16235 205
R8072 VSS.n17037 VSS.n16325 205
R8073 VSS.n16947 VSS.n16415 205
R8074 VSS.n16857 VSS.n16505 205
R8075 VSS.n16767 VSS.n16595 205
R8076 VSS.n11234 VSS.n11062 205
R8077 VSS.n11324 VSS.n10972 205
R8078 VSS.n11414 VSS.n10882 205
R8079 VSS.n13534 VSS.n10792 205
R8080 VSS.n13624 VSS.n10702 205
R8081 VSS.n13714 VSS.n10612 205
R8082 VSS.n13804 VSS.n10522 205
R8083 VSS.n13953 VSS.n10497 205
R8084 VSS.n9154 VSS.n9016 205
R8085 VSS.n10262 VSS.n9190 205
R8086 VSS.n10172 VSS.n9280 205
R8087 VSS.n10082 VSS.n9370 205
R8088 VSS.n9992 VSS.n9460 205
R8089 VSS.n9902 VSS.n9550 205
R8090 VSS.n9812 VSS.n9640 205
R8091 VSS.n10326 VSS.n10325 205
R8092 VSS.n5735 VSS.n5734 205
R8093 VSS.n5857 VSS.n5856 205
R8094 VSS.n5979 VSS.n5978 205
R8095 VSS.n6101 VSS.n6100 205
R8096 VSS.n6223 VSS.n6222 205
R8097 VSS.n6345 VSS.n6344 205
R8098 VSS.n6467 VSS.n6466 205
R8099 VSS.n6596 VSS.n3158 205
R8100 VSS.n1255 VSS.n1254 205
R8101 VSS.n1170 VSS.n98 205
R8102 VSS.n1080 VSS.n188 205
R8103 VSS.n990 VSS.n278 205
R8104 VSS.n900 VSS.n368 205
R8105 VSS.n810 VSS.n458 205
R8106 VSS.n720 VSS.n548 205
R8107 VSS.n15679 VSS.n15678 201.307
R8108 VSS.n15793 VSS.n15792 201.307
R8109 VSS.n15782 VSS.n15781 201.307
R8110 VSS.n15698 VSS.n15689 201.307
R8111 VSS.n15770 VSS.n15769 201.307
R8112 VSS.n15759 VSS.n15758 201.307
R8113 VSS.n15717 VSS.n15708 201.307
R8114 VSS.n15748 VSS.n15747 201.307
R8115 VSS.n15737 VSS.n15736 201.307
R8116 VSS.n15727 VSS.n14001 201.307
R8117 VSS.n16018 VSS.n16017 201.307
R8118 VSS.n16007 VSS.n16006 201.307
R8119 VSS.n15567 VSS.n15566 201.307
R8120 VSS.n15885 VSS.n15884 201.307
R8121 VSS.n15874 VSS.n15873 201.307
R8122 VSS.n15586 VSS.n15577 201.307
R8123 VSS.n15862 VSS.n15861 201.307
R8124 VSS.n15851 VSS.n15850 201.307
R8125 VSS.n15605 VSS.n15596 201.307
R8126 VSS.n15840 VSS.n15839 201.307
R8127 VSS.n15829 VSS.n15828 201.307
R8128 VSS.n15624 VSS.n15615 201.307
R8129 VSS.n15817 VSS.n15816 201.307
R8130 VSS.n15806 VSS.n15805 201.307
R8131 VSS.n15460 VSS.n14132 201.307
R8132 VSS.n15462 VSS.n14124 201.307
R8133 VSS.n15473 VSS.n15472 201.307
R8134 VSS.n15484 VSS.n15483 201.307
R8135 VSS.n15495 VSS.n14111 201.307
R8136 VSS.n15497 VSS.n14103 201.307
R8137 VSS.n15508 VSS.n15507 201.307
R8138 VSS.n15518 VSS.n15517 201.307
R8139 VSS.n15529 VSS.n14090 201.307
R8140 VSS.n15531 VSS.n14082 201.307
R8141 VSS.n15542 VSS.n15541 201.307
R8142 VSS.n15553 VSS.n15552 201.307
R8143 VSS.n15092 VSS.n15091 201.307
R8144 VSS.n15226 VSS.n15225 201.307
R8145 VSS.n15215 VSS.n15214 201.307
R8146 VSS.n15111 VSS.n15102 201.307
R8147 VSS.n15203 VSS.n15202 201.307
R8148 VSS.n15192 VSS.n15191 201.307
R8149 VSS.n15130 VSS.n15121 201.307
R8150 VSS.n15181 VSS.n15180 201.307
R8151 VSS.n15170 VSS.n15169 201.307
R8152 VSS.n15149 VSS.n15140 201.307
R8153 VSS.n15158 VSS.n15157 201.307
R8154 VSS.n15445 VSS.n15444 201.307
R8155 VSS.n14980 VSS.n14238 201.307
R8156 VSS.n15318 VSS.n15317 201.307
R8157 VSS.n15307 VSS.n15306 201.307
R8158 VSS.n14999 VSS.n14990 201.307
R8159 VSS.n15295 VSS.n15294 201.307
R8160 VSS.n15284 VSS.n15283 201.307
R8161 VSS.n15018 VSS.n15009 201.307
R8162 VSS.n15273 VSS.n15272 201.307
R8163 VSS.n15262 VSS.n15261 201.307
R8164 VSS.n15037 VSS.n15028 201.307
R8165 VSS.n15250 VSS.n15249 201.307
R8166 VSS.n15239 VSS.n15238 201.307
R8167 VSS.n14875 VSS.n14874 201.307
R8168 VSS.n14886 VSS.n14885 201.307
R8169 VSS.n14897 VSS.n14288 201.307
R8170 VSS.n14899 VSS.n14280 201.307
R8171 VSS.n14910 VSS.n14909 201.307
R8172 VSS.n14921 VSS.n14920 201.307
R8173 VSS.n14931 VSS.n14267 201.307
R8174 VSS.n14933 VSS.n14259 201.307
R8175 VSS.n14944 VSS.n14943 201.307
R8176 VSS.n14955 VSS.n14954 201.307
R8177 VSS.n14966 VSS.n14246 201.307
R8178 VSS.n14968 VSS.n14239 201.307
R8179 VSS.n14483 VSS.n14482 201.307
R8180 VSS.n14625 VSS.n14624 201.307
R8181 VSS.n14614 VSS.n14613 201.307
R8182 VSS.n14502 VSS.n14493 201.307
R8183 VSS.n14602 VSS.n14601 201.307
R8184 VSS.n14591 VSS.n14590 201.307
R8185 VSS.n14521 VSS.n14512 201.307
R8186 VSS.n14580 VSS.n14579 201.307
R8187 VSS.n14569 VSS.n14568 201.307
R8188 VSS.n14540 VSS.n14531 201.307
R8189 VSS.n14557 VSS.n14556 201.307
R8190 VSS.n14544 VSS.n14302 201.307
R8191 VSS.n14724 VSS.n14365 201.307
R8192 VSS.n14717 VSS.n14716 201.307
R8193 VSS.n14706 VSS.n14705 201.307
R8194 VSS.n14390 VSS.n14381 201.307
R8195 VSS.n14694 VSS.n14693 201.307
R8196 VSS.n14683 VSS.n14682 201.307
R8197 VSS.n14409 VSS.n14400 201.307
R8198 VSS.n14672 VSS.n14671 201.307
R8199 VSS.n14661 VSS.n14660 201.307
R8200 VSS.n14428 VSS.n14419 201.307
R8201 VSS.n14649 VSS.n14648 201.307
R8202 VSS.n14638 VSS.n14637 201.307
R8203 VSS.n11993 VSS.n11992 201.307
R8204 VSS.n12301 VSS.n12300 201.307
R8205 VSS.n12290 VSS.n12289 201.307
R8206 VSS.n12012 VSS.n12003 201.307
R8207 VSS.n12278 VSS.n12277 201.307
R8208 VSS.n12267 VSS.n12266 201.307
R8209 VSS.n12031 VSS.n12022 201.307
R8210 VSS.n12256 VSS.n12255 201.307
R8211 VSS.n12245 VSS.n12244 201.307
R8212 VSS.n12050 VSS.n12041 201.307
R8213 VSS.n12233 VSS.n12232 201.307
R8214 VSS.n12222 VSS.n12221 201.307
R8215 VSS.n11914 VSS.n11543 201.307
R8216 VSS.n12393 VSS.n12392 201.307
R8217 VSS.n12382 VSS.n12381 201.307
R8218 VSS.n11933 VSS.n11924 201.307
R8219 VSS.n12370 VSS.n12369 201.307
R8220 VSS.n12359 VSS.n12358 201.307
R8221 VSS.n11952 VSS.n11943 201.307
R8222 VSS.n12348 VSS.n12347 201.307
R8223 VSS.n12337 VSS.n12336 201.307
R8224 VSS.n11971 VSS.n11962 201.307
R8225 VSS.n12325 VSS.n12324 201.307
R8226 VSS.n12314 VSS.n12313 201.307
R8227 VSS.n11809 VSS.n11808 201.307
R8228 VSS.n11820 VSS.n11819 201.307
R8229 VSS.n11831 VSS.n11593 201.307
R8230 VSS.n11833 VSS.n11585 201.307
R8231 VSS.n11844 VSS.n11843 201.307
R8232 VSS.n11855 VSS.n11854 201.307
R8233 VSS.n11865 VSS.n11572 201.307
R8234 VSS.n11867 VSS.n11564 201.307
R8235 VSS.n11878 VSS.n11877 201.307
R8236 VSS.n11889 VSS.n11888 201.307
R8237 VSS.n11900 VSS.n11551 201.307
R8238 VSS.n11902 VSS.n11544 201.307
R8239 VSS.n11674 VSS.n11673 201.307
R8240 VSS.n11685 VSS.n11665 201.307
R8241 VSS.n11687 VSS.n11657 201.307
R8242 VSS.n11698 VSS.n11697 201.307
R8243 VSS.n11709 VSS.n11708 201.307
R8244 VSS.n11720 VSS.n11644 201.307
R8245 VSS.n11722 VSS.n11636 201.307
R8246 VSS.n11732 VSS.n11731 201.307
R8247 VSS.n11743 VSS.n11742 201.307
R8248 VSS.n11754 VSS.n11623 201.307
R8249 VSS.n11756 VSS.n11614 201.307
R8250 VSS.n11767 VSS.n11766 201.307
R8251 VSS.n13305 VSS.n13249 201.307
R8252 VSS.n13294 VSS.n13293 201.307
R8253 VSS.n13265 VSS.n13256 201.307
R8254 VSS.n13282 VSS.n13281 201.307
R8255 VSS.n13269 VSS.n11435 201.307
R8256 VSS.n13452 VSS.n13451 201.307
R8257 VSS.n13441 VSS.n13440 201.307
R8258 VSS.n11454 VSS.n11445 201.307
R8259 VSS.n13430 VSS.n13429 201.307
R8260 VSS.n13419 VSS.n13418 201.307
R8261 VSS.n11473 VSS.n11464 201.307
R8262 VSS.n13407 VSS.n13406 201.307
R8263 VSS.n13153 VSS.n13152 201.307
R8264 VSS.n13164 VSS.n12574 201.307
R8265 VSS.n13166 VSS.n12566 201.307
R8266 VSS.n13177 VSS.n13176 201.307
R8267 VSS.n13188 VSS.n13187 201.307
R8268 VSS.n13199 VSS.n12553 201.307
R8269 VSS.n13201 VSS.n12545 201.307
R8270 VSS.n13211 VSS.n13210 201.307
R8271 VSS.n13222 VSS.n13221 201.307
R8272 VSS.n13233 VSS.n12532 201.307
R8273 VSS.n13236 VSS.n13235 201.307
R8274 VSS.n13248 VSS.n13247 201.307
R8275 VSS.n13056 VSS.n12892 201.307
R8276 VSS.n13045 VSS.n13044 201.307
R8277 VSS.n12908 VSS.n12899 201.307
R8278 VSS.n13033 VSS.n13032 201.307
R8279 VSS.n13022 VSS.n13021 201.307
R8280 VSS.n12927 VSS.n12918 201.307
R8281 VSS.n13010 VSS.n13009 201.307
R8282 VSS.n13000 VSS.n12999 201.307
R8283 VSS.n12946 VSS.n12937 201.307
R8284 VSS.n12988 VSS.n12987 201.307
R8285 VSS.n12977 VSS.n12976 201.307
R8286 VSS.n12965 VSS.n12956 201.307
R8287 VSS.n12796 VSS.n12795 201.307
R8288 VSS.n12807 VSS.n12715 201.307
R8289 VSS.n12809 VSS.n12707 201.307
R8290 VSS.n12820 VSS.n12819 201.307
R8291 VSS.n12831 VSS.n12830 201.307
R8292 VSS.n12842 VSS.n12694 201.307
R8293 VSS.n12844 VSS.n12686 201.307
R8294 VSS.n12854 VSS.n12853 201.307
R8295 VSS.n12865 VSS.n12864 201.307
R8296 VSS.n12876 VSS.n12673 201.307
R8297 VSS.n12879 VSS.n12878 201.307
R8298 VSS.n12891 VSS.n12890 201.307
R8299 VSS.n7076 VSS.n6965 201.307
R8300 VSS.n7078 VSS.n7059 201.307
R8301 VSS.n7089 VSS.n7088 201.307
R8302 VSS.n7100 VSS.n7099 201.307
R8303 VSS.n7111 VSS.n7046 201.307
R8304 VSS.n7113 VSS.n7038 201.307
R8305 VSS.n7124 VSS.n7123 201.307
R8306 VSS.n7134 VSS.n7133 201.307
R8307 VSS.n7145 VSS.n7025 201.307
R8308 VSS.n7147 VSS.n7017 201.307
R8309 VSS.n7158 VSS.n7157 201.307
R8310 VSS.n7169 VSS.n7168 201.307
R8311 VSS.n8760 VSS.n7256 201.307
R8312 VSS.n8758 VSS.n8737 201.307
R8313 VSS.n8751 VSS.n6907 201.307
R8314 VSS.n8924 VSS.n8923 201.307
R8315 VSS.n8913 VSS.n8912 201.307
R8316 VSS.n6926 VSS.n6917 201.307
R8317 VSS.n8901 VSS.n8900 201.307
R8318 VSS.n8891 VSS.n8890 201.307
R8319 VSS.n6945 VSS.n6936 201.307
R8320 VSS.n8879 VSS.n8878 201.307
R8321 VSS.n8868 VSS.n8867 201.307
R8322 VSS.n6964 VSS.n6955 201.307
R8323 VSS.n8636 VSS.n8635 201.307
R8324 VSS.n8647 VSS.n8646 201.307
R8325 VSS.n8658 VSS.n7307 201.307
R8326 VSS.n8660 VSS.n7299 201.307
R8327 VSS.n8671 VSS.n8670 201.307
R8328 VSS.n8682 VSS.n8681 201.307
R8329 VSS.n8692 VSS.n7286 201.307
R8330 VSS.n8694 VSS.n7278 201.307
R8331 VSS.n8705 VSS.n8704 201.307
R8332 VSS.n8716 VSS.n8715 201.307
R8333 VSS.n8727 VSS.n7265 201.307
R8334 VSS.n8729 VSS.n7257 201.307
R8335 VSS.n8538 VSS.n7396 201.307
R8336 VSS.n8536 VSS.n8379 201.307
R8337 VSS.n8529 VSS.n8528 201.307
R8338 VSS.n8518 VSS.n8517 201.307
R8339 VSS.n8409 VSS.n8400 201.307
R8340 VSS.n8506 VSS.n8505 201.307
R8341 VSS.n8495 VSS.n8494 201.307
R8342 VSS.n8428 VSS.n8419 201.307
R8343 VSS.n8484 VSS.n8483 201.307
R8344 VSS.n8473 VSS.n8472 201.307
R8345 VSS.n8447 VSS.n8438 201.307
R8346 VSS.n8461 VSS.n8460 201.307
R8347 VSS.n8278 VSS.n8277 201.307
R8348 VSS.n8289 VSS.n8288 201.307
R8349 VSS.n8300 VSS.n7447 201.307
R8350 VSS.n8302 VSS.n7439 201.307
R8351 VSS.n8313 VSS.n8312 201.307
R8352 VSS.n8324 VSS.n8323 201.307
R8353 VSS.n8334 VSS.n7426 201.307
R8354 VSS.n8336 VSS.n7418 201.307
R8355 VSS.n8347 VSS.n8346 201.307
R8356 VSS.n8358 VSS.n8357 201.307
R8357 VSS.n8369 VSS.n7405 201.307
R8358 VSS.n8371 VSS.n7397 201.307
R8359 VSS.n8180 VSS.n7536 201.307
R8360 VSS.n8178 VSS.n8021 201.307
R8361 VSS.n8171 VSS.n8170 201.307
R8362 VSS.n8160 VSS.n8159 201.307
R8363 VSS.n8051 VSS.n8042 201.307
R8364 VSS.n8148 VSS.n8147 201.307
R8365 VSS.n8137 VSS.n8136 201.307
R8366 VSS.n8070 VSS.n8061 201.307
R8367 VSS.n8126 VSS.n8125 201.307
R8368 VSS.n8115 VSS.n8114 201.307
R8369 VSS.n8089 VSS.n8080 201.307
R8370 VSS.n8103 VSS.n8102 201.307
R8371 VSS.n7920 VSS.n7919 201.307
R8372 VSS.n7931 VSS.n7930 201.307
R8373 VSS.n7942 VSS.n7587 201.307
R8374 VSS.n7944 VSS.n7579 201.307
R8375 VSS.n7955 VSS.n7954 201.307
R8376 VSS.n7966 VSS.n7965 201.307
R8377 VSS.n7976 VSS.n7566 201.307
R8378 VSS.n7978 VSS.n7558 201.307
R8379 VSS.n7989 VSS.n7988 201.307
R8380 VSS.n8000 VSS.n7999 201.307
R8381 VSS.n8011 VSS.n7545 201.307
R8382 VSS.n8013 VSS.n7537 201.307
R8383 VSS.n7838 VSS.n7673 201.307
R8384 VSS.n7831 VSS.n7830 201.307
R8385 VSS.n7820 VSS.n7819 201.307
R8386 VSS.n7697 VSS.n7688 201.307
R8387 VSS.n7808 VSS.n7807 201.307
R8388 VSS.n7797 VSS.n7796 201.307
R8389 VSS.n7716 VSS.n7707 201.307
R8390 VSS.n7786 VSS.n7785 201.307
R8391 VSS.n7775 VSS.n7774 201.307
R8392 VSS.n7735 VSS.n7726 201.307
R8393 VSS.n7763 VSS.n7762 201.307
R8394 VSS.n7752 VSS.n7751 201.307
R8395 VSS.n5569 VSS.n5416 201.307
R8396 VSS.n5558 VSS.n5557 201.307
R8397 VSS.n5432 VSS.n5423 201.307
R8398 VSS.n5546 VSS.n5545 201.307
R8399 VSS.n5535 VSS.n5534 201.307
R8400 VSS.n5451 VSS.n5442 201.307
R8401 VSS.n5523 VSS.n5522 201.307
R8402 VSS.n5513 VSS.n5512 201.307
R8403 VSS.n5470 VSS.n5461 201.307
R8404 VSS.n5501 VSS.n5500 201.307
R8405 VSS.n5490 VSS.n5489 201.307
R8406 VSS.n5480 VSS.n3641 201.307
R8407 VSS.n5320 VSS.n5319 201.307
R8408 VSS.n5331 VSS.n3745 201.307
R8409 VSS.n5333 VSS.n3737 201.307
R8410 VSS.n5344 VSS.n5343 201.307
R8411 VSS.n5355 VSS.n5354 201.307
R8412 VSS.n5366 VSS.n3724 201.307
R8413 VSS.n5368 VSS.n3716 201.307
R8414 VSS.n5378 VSS.n5377 201.307
R8415 VSS.n5389 VSS.n5388 201.307
R8416 VSS.n5400 VSS.n3703 201.307
R8417 VSS.n5403 VSS.n5402 201.307
R8418 VSS.n5415 VSS.n5414 201.307
R8419 VSS.n5223 VSS.n5059 201.307
R8420 VSS.n5212 VSS.n5211 201.307
R8421 VSS.n5075 VSS.n5066 201.307
R8422 VSS.n5200 VSS.n5199 201.307
R8423 VSS.n5189 VSS.n5188 201.307
R8424 VSS.n5094 VSS.n5085 201.307
R8425 VSS.n5177 VSS.n5176 201.307
R8426 VSS.n5167 VSS.n5166 201.307
R8427 VSS.n5113 VSS.n5104 201.307
R8428 VSS.n5155 VSS.n5154 201.307
R8429 VSS.n5144 VSS.n5143 201.307
R8430 VSS.n5132 VSS.n5123 201.307
R8431 VSS.n4963 VSS.n4962 201.307
R8432 VSS.n4974 VSS.n3886 201.307
R8433 VSS.n4976 VSS.n3878 201.307
R8434 VSS.n4987 VSS.n4986 201.307
R8435 VSS.n4998 VSS.n4997 201.307
R8436 VSS.n5009 VSS.n3865 201.307
R8437 VSS.n5011 VSS.n3857 201.307
R8438 VSS.n5021 VSS.n5020 201.307
R8439 VSS.n5032 VSS.n5031 201.307
R8440 VSS.n5043 VSS.n3844 201.307
R8441 VSS.n5046 VSS.n5045 201.307
R8442 VSS.n5058 VSS.n5057 201.307
R8443 VSS.n4866 VSS.n4702 201.307
R8444 VSS.n4855 VSS.n4854 201.307
R8445 VSS.n4718 VSS.n4709 201.307
R8446 VSS.n4843 VSS.n4842 201.307
R8447 VSS.n4832 VSS.n4831 201.307
R8448 VSS.n4737 VSS.n4728 201.307
R8449 VSS.n4820 VSS.n4819 201.307
R8450 VSS.n4810 VSS.n4809 201.307
R8451 VSS.n4756 VSS.n4747 201.307
R8452 VSS.n4798 VSS.n4797 201.307
R8453 VSS.n4787 VSS.n4786 201.307
R8454 VSS.n4775 VSS.n4766 201.307
R8455 VSS.n4606 VSS.n4605 201.307
R8456 VSS.n4617 VSS.n4027 201.307
R8457 VSS.n4619 VSS.n4019 201.307
R8458 VSS.n4630 VSS.n4629 201.307
R8459 VSS.n4641 VSS.n4640 201.307
R8460 VSS.n4652 VSS.n4006 201.307
R8461 VSS.n4654 VSS.n3998 201.307
R8462 VSS.n4664 VSS.n4663 201.307
R8463 VSS.n4675 VSS.n4674 201.307
R8464 VSS.n4686 VSS.n3985 201.307
R8465 VSS.n4689 VSS.n4688 201.307
R8466 VSS.n4701 VSS.n4700 201.307
R8467 VSS.n4509 VSS.n4345 201.307
R8468 VSS.n4498 VSS.n4497 201.307
R8469 VSS.n4361 VSS.n4352 201.307
R8470 VSS.n4486 VSS.n4485 201.307
R8471 VSS.n4475 VSS.n4474 201.307
R8472 VSS.n4380 VSS.n4371 201.307
R8473 VSS.n4463 VSS.n4462 201.307
R8474 VSS.n4453 VSS.n4452 201.307
R8475 VSS.n4399 VSS.n4390 201.307
R8476 VSS.n4441 VSS.n4440 201.307
R8477 VSS.n4430 VSS.n4429 201.307
R8478 VSS.n4418 VSS.n4409 201.307
R8479 VSS.n4249 VSS.n4248 201.307
R8480 VSS.n4260 VSS.n4168 201.307
R8481 VSS.n4262 VSS.n4160 201.307
R8482 VSS.n4273 VSS.n4272 201.307
R8483 VSS.n4284 VSS.n4283 201.307
R8484 VSS.n4295 VSS.n4147 201.307
R8485 VSS.n4297 VSS.n4139 201.307
R8486 VSS.n4307 VSS.n4306 201.307
R8487 VSS.n4318 VSS.n4317 201.307
R8488 VSS.n4329 VSS.n4126 201.307
R8489 VSS.n4332 VSS.n4331 201.307
R8490 VSS.n4344 VSS.n4343 201.307
R8491 VSS.n2808 VSS.n2807 201.307
R8492 VSS.n2959 VSS.n2958 201.307
R8493 VSS.n2948 VSS.n2947 201.307
R8494 VSS.n2827 VSS.n2818 201.307
R8495 VSS.n2936 VSS.n2935 201.307
R8496 VSS.n2925 VSS.n2924 201.307
R8497 VSS.n2846 VSS.n2837 201.307
R8498 VSS.n2914 VSS.n2913 201.307
R8499 VSS.n2903 VSS.n2902 201.307
R8500 VSS.n2865 VSS.n2856 201.307
R8501 VSS.n2891 VSS.n2890 201.307
R8502 VSS.n2880 VSS.n2879 201.307
R8503 VSS.n2701 VSS.n1373 201.307
R8504 VSS.n2703 VSS.n1365 201.307
R8505 VSS.n2714 VSS.n2713 201.307
R8506 VSS.n2725 VSS.n2724 201.307
R8507 VSS.n2736 VSS.n1352 201.307
R8508 VSS.n2738 VSS.n1344 201.307
R8509 VSS.n2749 VSS.n2748 201.307
R8510 VSS.n2759 VSS.n2758 201.307
R8511 VSS.n2770 VSS.n1331 201.307
R8512 VSS.n2772 VSS.n1323 201.307
R8513 VSS.n2783 VSS.n2782 201.307
R8514 VSS.n2794 VSS.n2793 201.307
R8515 VSS.n2333 VSS.n2332 201.307
R8516 VSS.n2467 VSS.n2466 201.307
R8517 VSS.n2456 VSS.n2455 201.307
R8518 VSS.n2352 VSS.n2343 201.307
R8519 VSS.n2444 VSS.n2443 201.307
R8520 VSS.n2433 VSS.n2432 201.307
R8521 VSS.n2371 VSS.n2362 201.307
R8522 VSS.n2422 VSS.n2421 201.307
R8523 VSS.n2411 VSS.n2410 201.307
R8524 VSS.n2390 VSS.n2381 201.307
R8525 VSS.n2399 VSS.n2398 201.307
R8526 VSS.n2686 VSS.n2685 201.307
R8527 VSS.n2221 VSS.n1479 201.307
R8528 VSS.n2559 VSS.n2558 201.307
R8529 VSS.n2548 VSS.n2547 201.307
R8530 VSS.n2240 VSS.n2231 201.307
R8531 VSS.n2536 VSS.n2535 201.307
R8532 VSS.n2525 VSS.n2524 201.307
R8533 VSS.n2259 VSS.n2250 201.307
R8534 VSS.n2514 VSS.n2513 201.307
R8535 VSS.n2503 VSS.n2502 201.307
R8536 VSS.n2278 VSS.n2269 201.307
R8537 VSS.n2491 VSS.n2490 201.307
R8538 VSS.n2480 VSS.n2479 201.307
R8539 VSS.n2116 VSS.n2115 201.307
R8540 VSS.n2127 VSS.n2126 201.307
R8541 VSS.n2138 VSS.n1529 201.307
R8542 VSS.n2140 VSS.n1521 201.307
R8543 VSS.n2151 VSS.n2150 201.307
R8544 VSS.n2162 VSS.n2161 201.307
R8545 VSS.n2172 VSS.n1508 201.307
R8546 VSS.n2174 VSS.n1500 201.307
R8547 VSS.n2185 VSS.n2184 201.307
R8548 VSS.n2196 VSS.n2195 201.307
R8549 VSS.n2207 VSS.n1487 201.307
R8550 VSS.n2209 VSS.n1480 201.307
R8551 VSS.n1724 VSS.n1723 201.307
R8552 VSS.n1866 VSS.n1865 201.307
R8553 VSS.n1855 VSS.n1854 201.307
R8554 VSS.n1743 VSS.n1734 201.307
R8555 VSS.n1843 VSS.n1842 201.307
R8556 VSS.n1832 VSS.n1831 201.307
R8557 VSS.n1762 VSS.n1753 201.307
R8558 VSS.n1821 VSS.n1820 201.307
R8559 VSS.n1810 VSS.n1809 201.307
R8560 VSS.n1781 VSS.n1772 201.307
R8561 VSS.n1798 VSS.n1797 201.307
R8562 VSS.n1785 VSS.n1543 201.307
R8563 VSS.n1965 VSS.n1606 201.307
R8564 VSS.n1958 VSS.n1957 201.307
R8565 VSS.n1947 VSS.n1946 201.307
R8566 VSS.n1631 VSS.n1622 201.307
R8567 VSS.n1935 VSS.n1934 201.307
R8568 VSS.n1924 VSS.n1923 201.307
R8569 VSS.n1650 VSS.n1641 201.307
R8570 VSS.n1913 VSS.n1912 201.307
R8571 VSS.n1902 VSS.n1901 201.307
R8572 VSS.n1669 VSS.n1660 201.307
R8573 VSS.n1890 VSS.n1889 201.307
R8574 VSS.n1879 VSS.n1878 201.307
R8575 VSS.n10437 VSS.n10433 195.413
R8576 VSS.n10437 VSS.n10436 195.413
R8577 VSS.n6826 VSS.n6757 195.049
R8578 VSS.n10433 sky130_asc_nfet_01v8_lvt_9_0/SOURCE 189.013
R8579 VSS.n6802 VSS.n6770 187.247
R8580 VSS.t30 VSS.n16031 185
R8581 VSS.n17414 VSS.n17413 185
R8582 VSS.n17410 VSS.n17409 185
R8583 VSS.n17406 VSS.n17405 185
R8584 VSS.n17403 VSS.n17402 185
R8585 VSS.n17449 VSS.n17448 185
R8586 VSS.n17458 VSS.n17457 185
R8587 VSS.n17393 VSS.n17392 185
R8588 VSS.n17328 VSS.n17327 185
R8589 VSS.n17417 VSS.n17416 185
R8590 VSS.n17385 VSS.t30 185
R8591 VSS.n17460 VSS.n16034 185
R8592 VSS.t30 VSS.n16034 185
R8593 VSS.t30 VSS.n16037 185
R8594 VSS.n17460 VSS.n16037 185
R8595 VSS.n17460 VSS.n16033 185
R8596 VSS.t30 VSS.n16033 185
R8597 VSS.t30 VSS.n16038 185
R8598 VSS.n17460 VSS.n16038 185
R8599 VSS.n17460 VSS.n16032 185
R8600 VSS.t30 VSS.n16032 185
R8601 VSS.t30 VSS.n16039 185
R8602 VSS.n17460 VSS.n16039 185
R8603 VSS.n17460 VSS.n16031 185
R8604 VSS.t54 VSS.n16075 185
R8605 VSS.n17251 VSS.n17250 185
R8606 VSS.n17248 VSS.n16079 185
R8607 VSS.n17245 VSS.n17244 185
R8608 VSS.n17241 VSS.n17240 185
R8609 VSS.n17237 VSS.n17236 185
R8610 VSS.n17234 VSS.n17233 185
R8611 VSS.n17293 VSS.n17292 185
R8612 VSS.n17302 VSS.n17301 185
R8613 VSS.n17223 VSS.n16082 185
R8614 VSS.n17305 VSS.n16082 185
R8615 VSS.t54 VSS.n16076 185
R8616 VSS.n17305 VSS.n16076 185
R8617 VSS.n17305 VSS.n16073 185
R8618 VSS.t54 VSS.n16073 185
R8619 VSS.t54 VSS.n16077 185
R8620 VSS.n17305 VSS.n16077 185
R8621 VSS.n17305 VSS.n16072 185
R8622 VSS.t54 VSS.n16072 185
R8623 VSS.t54 VSS.n16078 185
R8624 VSS.n17305 VSS.n16078 185
R8625 VSS.n17305 VSS.n16071 185
R8626 VSS.t54 VSS.n16071 185
R8627 VSS.t54 VSS.n17306 185
R8628 VSS.n17306 VSS.n17305 185
R8629 VSS.t50 VSS.n16165 185
R8630 VSS.n17161 VSS.n17160 185
R8631 VSS.n17158 VSS.n16169 185
R8632 VSS.n17155 VSS.n17154 185
R8633 VSS.n17151 VSS.n17150 185
R8634 VSS.n17147 VSS.n17146 185
R8635 VSS.n17144 VSS.n17143 185
R8636 VSS.n17203 VSS.n17202 185
R8637 VSS.n17212 VSS.n17211 185
R8638 VSS.n17133 VSS.n16172 185
R8639 VSS.n17215 VSS.n16172 185
R8640 VSS.t50 VSS.n16166 185
R8641 VSS.n17215 VSS.n16166 185
R8642 VSS.n17215 VSS.n16163 185
R8643 VSS.t50 VSS.n16163 185
R8644 VSS.t50 VSS.n16167 185
R8645 VSS.n17215 VSS.n16167 185
R8646 VSS.n17215 VSS.n16162 185
R8647 VSS.t50 VSS.n16162 185
R8648 VSS.t50 VSS.n16168 185
R8649 VSS.n17215 VSS.n16168 185
R8650 VSS.n17215 VSS.n16161 185
R8651 VSS.t50 VSS.n16161 185
R8652 VSS.t50 VSS.n17216 185
R8653 VSS.n17216 VSS.n17215 185
R8654 VSS.t42 VSS.n16255 185
R8655 VSS.n17071 VSS.n17070 185
R8656 VSS.n17068 VSS.n16259 185
R8657 VSS.n17065 VSS.n17064 185
R8658 VSS.n17061 VSS.n17060 185
R8659 VSS.n17057 VSS.n17056 185
R8660 VSS.n17054 VSS.n17053 185
R8661 VSS.n17113 VSS.n17112 185
R8662 VSS.n17122 VSS.n17121 185
R8663 VSS.n17043 VSS.n16262 185
R8664 VSS.n17125 VSS.n16262 185
R8665 VSS.t42 VSS.n16256 185
R8666 VSS.n17125 VSS.n16256 185
R8667 VSS.n17125 VSS.n16253 185
R8668 VSS.t42 VSS.n16253 185
R8669 VSS.t42 VSS.n16257 185
R8670 VSS.n17125 VSS.n16257 185
R8671 VSS.n17125 VSS.n16252 185
R8672 VSS.t42 VSS.n16252 185
R8673 VSS.t42 VSS.n16258 185
R8674 VSS.n17125 VSS.n16258 185
R8675 VSS.n17125 VSS.n16251 185
R8676 VSS.t42 VSS.n16251 185
R8677 VSS.t42 VSS.n17126 185
R8678 VSS.n17126 VSS.n17125 185
R8679 VSS.t68 VSS.n16345 185
R8680 VSS.n16981 VSS.n16980 185
R8681 VSS.n16978 VSS.n16349 185
R8682 VSS.n16975 VSS.n16974 185
R8683 VSS.n16971 VSS.n16970 185
R8684 VSS.n16967 VSS.n16966 185
R8685 VSS.n16964 VSS.n16963 185
R8686 VSS.n17023 VSS.n17022 185
R8687 VSS.n17032 VSS.n17031 185
R8688 VSS.n16953 VSS.n16352 185
R8689 VSS.n17035 VSS.n16352 185
R8690 VSS.t68 VSS.n16346 185
R8691 VSS.n17035 VSS.n16346 185
R8692 VSS.n17035 VSS.n16343 185
R8693 VSS.t68 VSS.n16343 185
R8694 VSS.t68 VSS.n16347 185
R8695 VSS.n17035 VSS.n16347 185
R8696 VSS.n17035 VSS.n16342 185
R8697 VSS.t68 VSS.n16342 185
R8698 VSS.t68 VSS.n16348 185
R8699 VSS.n17035 VSS.n16348 185
R8700 VSS.n17035 VSS.n16341 185
R8701 VSS.t68 VSS.n16341 185
R8702 VSS.t68 VSS.n17036 185
R8703 VSS.n17036 VSS.n17035 185
R8704 VSS.t74 VSS.n16435 185
R8705 VSS.n16891 VSS.n16890 185
R8706 VSS.n16888 VSS.n16439 185
R8707 VSS.n16885 VSS.n16884 185
R8708 VSS.n16881 VSS.n16880 185
R8709 VSS.n16877 VSS.n16876 185
R8710 VSS.n16874 VSS.n16873 185
R8711 VSS.n16933 VSS.n16932 185
R8712 VSS.n16942 VSS.n16941 185
R8713 VSS.n16863 VSS.n16442 185
R8714 VSS.n16945 VSS.n16442 185
R8715 VSS.t74 VSS.n16436 185
R8716 VSS.n16945 VSS.n16436 185
R8717 VSS.n16945 VSS.n16433 185
R8718 VSS.t74 VSS.n16433 185
R8719 VSS.t74 VSS.n16437 185
R8720 VSS.n16945 VSS.n16437 185
R8721 VSS.n16945 VSS.n16432 185
R8722 VSS.t74 VSS.n16432 185
R8723 VSS.t74 VSS.n16438 185
R8724 VSS.n16945 VSS.n16438 185
R8725 VSS.n16945 VSS.n16431 185
R8726 VSS.t74 VSS.n16431 185
R8727 VSS.t74 VSS.n16946 185
R8728 VSS.n16946 VSS.n16945 185
R8729 VSS.t90 VSS.n16525 185
R8730 VSS.n16801 VSS.n16800 185
R8731 VSS.n16798 VSS.n16529 185
R8732 VSS.n16795 VSS.n16794 185
R8733 VSS.n16791 VSS.n16790 185
R8734 VSS.n16787 VSS.n16786 185
R8735 VSS.n16784 VSS.n16783 185
R8736 VSS.n16843 VSS.n16842 185
R8737 VSS.n16852 VSS.n16851 185
R8738 VSS.n16773 VSS.n16532 185
R8739 VSS.n16855 VSS.n16532 185
R8740 VSS.t90 VSS.n16526 185
R8741 VSS.n16855 VSS.n16526 185
R8742 VSS.n16855 VSS.n16523 185
R8743 VSS.t90 VSS.n16523 185
R8744 VSS.t90 VSS.n16527 185
R8745 VSS.n16855 VSS.n16527 185
R8746 VSS.n16855 VSS.n16522 185
R8747 VSS.t90 VSS.n16522 185
R8748 VSS.t90 VSS.n16528 185
R8749 VSS.n16855 VSS.n16528 185
R8750 VSS.n16855 VSS.n16521 185
R8751 VSS.t90 VSS.n16521 185
R8752 VSS.t90 VSS.n16856 185
R8753 VSS.n16856 VSS.n16855 185
R8754 VSS.t28 VSS.n16615 185
R8755 VSS.n16711 VSS.n16710 185
R8756 VSS.n16708 VSS.n16619 185
R8757 VSS.n16705 VSS.n16704 185
R8758 VSS.n16701 VSS.n16700 185
R8759 VSS.n16697 VSS.n16696 185
R8760 VSS.n16694 VSS.n16693 185
R8761 VSS.n16753 VSS.n16752 185
R8762 VSS.n16762 VSS.n16761 185
R8763 VSS.n16683 VSS.n16622 185
R8764 VSS.n16765 VSS.n16622 185
R8765 VSS.t28 VSS.n16616 185
R8766 VSS.n16765 VSS.n16616 185
R8767 VSS.n16765 VSS.n16613 185
R8768 VSS.t28 VSS.n16613 185
R8769 VSS.t28 VSS.n16617 185
R8770 VSS.n16765 VSS.n16617 185
R8771 VSS.n16765 VSS.n16612 185
R8772 VSS.t28 VSS.n16612 185
R8773 VSS.t28 VSS.n16618 185
R8774 VSS.n16765 VSS.n16618 185
R8775 VSS.n16765 VSS.n16611 185
R8776 VSS.t28 VSS.n16611 185
R8777 VSS.t28 VSS.n16766 185
R8778 VSS.n16766 VSS.n16765 185
R8779 VSS.t58 VSS.n11082 185
R8780 VSS.n11174 VSS.n11173 185
R8781 VSS.n11171 VSS.n11086 185
R8782 VSS.n11179 VSS.n11177 185
R8783 VSS.n11168 VSS.n11167 185
R8784 VSS.n11164 VSS.n11163 185
R8785 VSS.n11161 VSS.n11160 185
R8786 VSS.n11221 VSS.n11220 185
R8787 VSS.n11230 VSS.n11229 185
R8788 VSS.n11151 VSS.n11150 185
R8789 VSS.t58 VSS.n11083 185
R8790 VSS.n11232 VSS.n11080 185
R8791 VSS.t58 VSS.n11080 185
R8792 VSS.t58 VSS.n11084 185
R8793 VSS.n11232 VSS.n11084 185
R8794 VSS.n11232 VSS.n11079 185
R8795 VSS.t58 VSS.n11079 185
R8796 VSS.t58 VSS.n11085 185
R8797 VSS.n11232 VSS.n11085 185
R8798 VSS.n11232 VSS.n11078 185
R8799 VSS.t58 VSS.n11078 185
R8800 VSS.t58 VSS.n11233 185
R8801 VSS.n11233 VSS.n11232 185
R8802 VSS.n11232 VSS.n11082 185
R8803 VSS.t32 VSS.n10992 185
R8804 VSS.n11264 VSS.n11263 185
R8805 VSS.n11261 VSS.n10996 185
R8806 VSS.n11269 VSS.n11267 185
R8807 VSS.n11258 VSS.n11257 185
R8808 VSS.n11254 VSS.n11253 185
R8809 VSS.n11251 VSS.n11250 185
R8810 VSS.n11311 VSS.n11310 185
R8811 VSS.n11320 VSS.n11319 185
R8812 VSS.n11241 VSS.n11240 185
R8813 VSS.t32 VSS.n10993 185
R8814 VSS.n11322 VSS.n10990 185
R8815 VSS.t32 VSS.n10990 185
R8816 VSS.t32 VSS.n10994 185
R8817 VSS.n11322 VSS.n10994 185
R8818 VSS.n11322 VSS.n10989 185
R8819 VSS.t32 VSS.n10989 185
R8820 VSS.t32 VSS.n10995 185
R8821 VSS.n11322 VSS.n10995 185
R8822 VSS.n11322 VSS.n10988 185
R8823 VSS.t32 VSS.n10988 185
R8824 VSS.t32 VSS.n11323 185
R8825 VSS.n11323 VSS.n11322 185
R8826 VSS.n11322 VSS.n10992 185
R8827 VSS.t92 VSS.n10902 185
R8828 VSS.n11354 VSS.n11353 185
R8829 VSS.n11351 VSS.n10906 185
R8830 VSS.n11359 VSS.n11357 185
R8831 VSS.n11348 VSS.n11347 185
R8832 VSS.n11344 VSS.n11343 185
R8833 VSS.n11341 VSS.n11340 185
R8834 VSS.n11401 VSS.n11400 185
R8835 VSS.n11410 VSS.n11409 185
R8836 VSS.n11331 VSS.n11330 185
R8837 VSS.t92 VSS.n10903 185
R8838 VSS.n11412 VSS.n10900 185
R8839 VSS.t92 VSS.n10900 185
R8840 VSS.t92 VSS.n10904 185
R8841 VSS.n11412 VSS.n10904 185
R8842 VSS.n11412 VSS.n10899 185
R8843 VSS.t92 VSS.n10899 185
R8844 VSS.t92 VSS.n10905 185
R8845 VSS.n11412 VSS.n10905 185
R8846 VSS.n11412 VSS.n10898 185
R8847 VSS.t92 VSS.n10898 185
R8848 VSS.t92 VSS.n11413 185
R8849 VSS.n11413 VSS.n11412 185
R8850 VSS.n11412 VSS.n10902 185
R8851 VSS.t88 VSS.n10812 185
R8852 VSS.n13473 VSS.n13472 185
R8853 VSS.n13470 VSS.n10816 185
R8854 VSS.n13478 VSS.n13476 185
R8855 VSS.n13467 VSS.n13466 185
R8856 VSS.n13463 VSS.n13462 185
R8857 VSS.n13460 VSS.n13459 185
R8858 VSS.n13521 VSS.n13520 185
R8859 VSS.n13530 VSS.n13529 185
R8860 VSS.n11421 VSS.n11420 185
R8861 VSS.t88 VSS.n10813 185
R8862 VSS.n13532 VSS.n10810 185
R8863 VSS.t88 VSS.n10810 185
R8864 VSS.t88 VSS.n10814 185
R8865 VSS.n13532 VSS.n10814 185
R8866 VSS.n13532 VSS.n10809 185
R8867 VSS.t88 VSS.n10809 185
R8868 VSS.t88 VSS.n10815 185
R8869 VSS.n13532 VSS.n10815 185
R8870 VSS.n13532 VSS.n10808 185
R8871 VSS.t88 VSS.n10808 185
R8872 VSS.t88 VSS.n13533 185
R8873 VSS.n13533 VSS.n13532 185
R8874 VSS.n13532 VSS.n10812 185
R8875 VSS.t72 VSS.n10722 185
R8876 VSS.n13564 VSS.n13563 185
R8877 VSS.n13561 VSS.n10726 185
R8878 VSS.n13569 VSS.n13567 185
R8879 VSS.n13558 VSS.n13557 185
R8880 VSS.n13554 VSS.n13553 185
R8881 VSS.n13551 VSS.n13550 185
R8882 VSS.n13611 VSS.n13610 185
R8883 VSS.n13620 VSS.n13619 185
R8884 VSS.n13541 VSS.n13540 185
R8885 VSS.t72 VSS.n10723 185
R8886 VSS.n13622 VSS.n10720 185
R8887 VSS.t72 VSS.n10720 185
R8888 VSS.t72 VSS.n10724 185
R8889 VSS.n13622 VSS.n10724 185
R8890 VSS.n13622 VSS.n10719 185
R8891 VSS.t72 VSS.n10719 185
R8892 VSS.t72 VSS.n10725 185
R8893 VSS.n13622 VSS.n10725 185
R8894 VSS.n13622 VSS.n10718 185
R8895 VSS.t72 VSS.n10718 185
R8896 VSS.t72 VSS.n13623 185
R8897 VSS.n13623 VSS.n13622 185
R8898 VSS.n13622 VSS.n10722 185
R8899 VSS.t78 VSS.n10632 185
R8900 VSS.n13654 VSS.n13653 185
R8901 VSS.n13651 VSS.n10636 185
R8902 VSS.n13659 VSS.n13657 185
R8903 VSS.n13648 VSS.n13647 185
R8904 VSS.n13644 VSS.n13643 185
R8905 VSS.n13641 VSS.n13640 185
R8906 VSS.n13701 VSS.n13700 185
R8907 VSS.n13710 VSS.n13709 185
R8908 VSS.n13631 VSS.n13630 185
R8909 VSS.t78 VSS.n10633 185
R8910 VSS.n13712 VSS.n10630 185
R8911 VSS.t78 VSS.n10630 185
R8912 VSS.t78 VSS.n10634 185
R8913 VSS.n13712 VSS.n10634 185
R8914 VSS.n13712 VSS.n10629 185
R8915 VSS.t78 VSS.n10629 185
R8916 VSS.t78 VSS.n10635 185
R8917 VSS.n13712 VSS.n10635 185
R8918 VSS.n13712 VSS.n10628 185
R8919 VSS.t78 VSS.n10628 185
R8920 VSS.t78 VSS.n13713 185
R8921 VSS.n13713 VSS.n13712 185
R8922 VSS.n13712 VSS.n10632 185
R8923 VSS.t82 VSS.n10542 185
R8924 VSS.n13744 VSS.n13743 185
R8925 VSS.n13741 VSS.n10546 185
R8926 VSS.n13749 VSS.n13747 185
R8927 VSS.n13738 VSS.n13737 185
R8928 VSS.n13734 VSS.n13733 185
R8929 VSS.n13731 VSS.n13730 185
R8930 VSS.n13791 VSS.n13790 185
R8931 VSS.n13800 VSS.n13799 185
R8932 VSS.n13721 VSS.n13720 185
R8933 VSS.t82 VSS.n10543 185
R8934 VSS.n13802 VSS.n10540 185
R8935 VSS.t82 VSS.n10540 185
R8936 VSS.t82 VSS.n10544 185
R8937 VSS.n13802 VSS.n10544 185
R8938 VSS.n13802 VSS.n10539 185
R8939 VSS.t82 VSS.n10539 185
R8940 VSS.t82 VSS.n10545 185
R8941 VSS.n13802 VSS.n10545 185
R8942 VSS.n13802 VSS.n10538 185
R8943 VSS.t82 VSS.n10538 185
R8944 VSS.t82 VSS.n13803 185
R8945 VSS.n13803 VSS.n13802 185
R8946 VSS.n13802 VSS.n10542 185
R8947 VSS.t62 VSS.n10500 185
R8948 VSS.n13915 VSS.n13914 185
R8949 VSS.n13910 VSS.n13909 185
R8950 VSS.n13906 VSS.n13905 185
R8951 VSS.n13903 VSS.n13902 185
R8952 VSS.n13941 VSS.n13940 185
R8953 VSS.n13950 VSS.n13949 185
R8954 VSS.n13893 VSS.n13892 185
R8955 VSS.n13825 VSS.n13824 185
R8956 VSS.n13956 VSS.n13955 185
R8957 VSS.n13885 VSS.t62 185
R8958 VSS.n13952 VSS.n10503 185
R8959 VSS.t62 VSS.n10503 185
R8960 VSS.t62 VSS.n10505 185
R8961 VSS.n13952 VSS.n10505 185
R8962 VSS.n13952 VSS.n10502 185
R8963 VSS.t62 VSS.n10502 185
R8964 VSS.t62 VSS.n10506 185
R8965 VSS.n13952 VSS.n10506 185
R8966 VSS.n13952 VSS.n10501 185
R8967 VSS.t62 VSS.n10501 185
R8968 VSS.t62 VSS.n10507 185
R8969 VSS.n13952 VSS.n10507 185
R8970 VSS.n13952 VSS.n10500 185
R8971 VSS.n9094 VSS.n9093 185
R8972 VSS.n9078 VSS.n9077 185
R8973 VSS.n9062 VSS.n9061 185
R8974 VSS.n9046 VSS.n9045 185
R8975 VSS.n9158 VSS.n9157 185
R8976 VSS.n9038 VSS.n9037 185
R8977 VSS.n9054 VSS.n9053 185
R8978 VSS.n9070 VSS.n9069 185
R8979 VSS.n9086 VSS.n9085 185
R8980 VSS.t34 VSS.n9210 185
R8981 VSS.n10206 VSS.n10205 185
R8982 VSS.n10203 VSS.n9214 185
R8983 VSS.n10200 VSS.n10199 185
R8984 VSS.n10196 VSS.n10195 185
R8985 VSS.n10192 VSS.n10191 185
R8986 VSS.n10189 VSS.n10188 185
R8987 VSS.n10248 VSS.n10247 185
R8988 VSS.n10257 VSS.n10256 185
R8989 VSS.n10178 VSS.n9217 185
R8990 VSS.n10260 VSS.n9217 185
R8991 VSS.t34 VSS.n9211 185
R8992 VSS.n10260 VSS.n9211 185
R8993 VSS.n10260 VSS.n9208 185
R8994 VSS.t34 VSS.n9208 185
R8995 VSS.t34 VSS.n9212 185
R8996 VSS.n10260 VSS.n9212 185
R8997 VSS.n10260 VSS.n9207 185
R8998 VSS.t34 VSS.n9207 185
R8999 VSS.t34 VSS.n9213 185
R9000 VSS.n10260 VSS.n9213 185
R9001 VSS.n10260 VSS.n9206 185
R9002 VSS.t34 VSS.n9206 185
R9003 VSS.t34 VSS.n10261 185
R9004 VSS.n10261 VSS.n10260 185
R9005 VSS.t26 VSS.n9300 185
R9006 VSS.n10116 VSS.n10115 185
R9007 VSS.n10113 VSS.n9304 185
R9008 VSS.n10110 VSS.n10109 185
R9009 VSS.n10106 VSS.n10105 185
R9010 VSS.n10102 VSS.n10101 185
R9011 VSS.n10099 VSS.n10098 185
R9012 VSS.n10158 VSS.n10157 185
R9013 VSS.n10167 VSS.n10166 185
R9014 VSS.n10088 VSS.n9307 185
R9015 VSS.n10170 VSS.n9307 185
R9016 VSS.t26 VSS.n9301 185
R9017 VSS.n10170 VSS.n9301 185
R9018 VSS.n10170 VSS.n9298 185
R9019 VSS.t26 VSS.n9298 185
R9020 VSS.t26 VSS.n9302 185
R9021 VSS.n10170 VSS.n9302 185
R9022 VSS.n10170 VSS.n9297 185
R9023 VSS.t26 VSS.n9297 185
R9024 VSS.t26 VSS.n9303 185
R9025 VSS.n10170 VSS.n9303 185
R9026 VSS.n10170 VSS.n9296 185
R9027 VSS.t26 VSS.n9296 185
R9028 VSS.t26 VSS.n10171 185
R9029 VSS.n10171 VSS.n10170 185
R9030 VSS.t52 VSS.n9390 185
R9031 VSS.n10026 VSS.n10025 185
R9032 VSS.n10023 VSS.n9394 185
R9033 VSS.n10020 VSS.n10019 185
R9034 VSS.n10016 VSS.n10015 185
R9035 VSS.n10012 VSS.n10011 185
R9036 VSS.n10009 VSS.n10008 185
R9037 VSS.n10068 VSS.n10067 185
R9038 VSS.n10077 VSS.n10076 185
R9039 VSS.n9998 VSS.n9397 185
R9040 VSS.n10080 VSS.n9397 185
R9041 VSS.t52 VSS.n9391 185
R9042 VSS.n10080 VSS.n9391 185
R9043 VSS.n10080 VSS.n9388 185
R9044 VSS.t52 VSS.n9388 185
R9045 VSS.t52 VSS.n9392 185
R9046 VSS.n10080 VSS.n9392 185
R9047 VSS.n10080 VSS.n9387 185
R9048 VSS.t52 VSS.n9387 185
R9049 VSS.t52 VSS.n9393 185
R9050 VSS.n10080 VSS.n9393 185
R9051 VSS.n10080 VSS.n9386 185
R9052 VSS.t52 VSS.n9386 185
R9053 VSS.t52 VSS.n10081 185
R9054 VSS.n10081 VSS.n10080 185
R9055 VSS.t56 VSS.n9480 185
R9056 VSS.n9936 VSS.n9935 185
R9057 VSS.n9933 VSS.n9484 185
R9058 VSS.n9930 VSS.n9929 185
R9059 VSS.n9926 VSS.n9925 185
R9060 VSS.n9922 VSS.n9921 185
R9061 VSS.n9919 VSS.n9918 185
R9062 VSS.n9978 VSS.n9977 185
R9063 VSS.n9987 VSS.n9986 185
R9064 VSS.n9908 VSS.n9487 185
R9065 VSS.n9990 VSS.n9487 185
R9066 VSS.t56 VSS.n9481 185
R9067 VSS.n9990 VSS.n9481 185
R9068 VSS.n9990 VSS.n9478 185
R9069 VSS.t56 VSS.n9478 185
R9070 VSS.t56 VSS.n9482 185
R9071 VSS.n9990 VSS.n9482 185
R9072 VSS.n9990 VSS.n9477 185
R9073 VSS.t56 VSS.n9477 185
R9074 VSS.t56 VSS.n9483 185
R9075 VSS.n9990 VSS.n9483 185
R9076 VSS.n9990 VSS.n9476 185
R9077 VSS.t56 VSS.n9476 185
R9078 VSS.t56 VSS.n9991 185
R9079 VSS.n9991 VSS.n9990 185
R9080 VSS.t80 VSS.n9570 185
R9081 VSS.n9846 VSS.n9845 185
R9082 VSS.n9843 VSS.n9574 185
R9083 VSS.n9840 VSS.n9839 185
R9084 VSS.n9836 VSS.n9835 185
R9085 VSS.n9832 VSS.n9831 185
R9086 VSS.n9829 VSS.n9828 185
R9087 VSS.n9888 VSS.n9887 185
R9088 VSS.n9897 VSS.n9896 185
R9089 VSS.n9818 VSS.n9577 185
R9090 VSS.n9900 VSS.n9577 185
R9091 VSS.t80 VSS.n9571 185
R9092 VSS.n9900 VSS.n9571 185
R9093 VSS.n9900 VSS.n9568 185
R9094 VSS.t80 VSS.n9568 185
R9095 VSS.t80 VSS.n9572 185
R9096 VSS.n9900 VSS.n9572 185
R9097 VSS.n9900 VSS.n9567 185
R9098 VSS.t80 VSS.n9567 185
R9099 VSS.t80 VSS.n9573 185
R9100 VSS.n9900 VSS.n9573 185
R9101 VSS.n9900 VSS.n9566 185
R9102 VSS.t80 VSS.n9566 185
R9103 VSS.t80 VSS.n9901 185
R9104 VSS.n9901 VSS.n9900 185
R9105 VSS.t18 VSS.n9660 185
R9106 VSS.n9756 VSS.n9755 185
R9107 VSS.n9753 VSS.n9664 185
R9108 VSS.n9750 VSS.n9749 185
R9109 VSS.n9746 VSS.n9745 185
R9110 VSS.n9742 VSS.n9741 185
R9111 VSS.n9739 VSS.n9738 185
R9112 VSS.n9798 VSS.n9797 185
R9113 VSS.n9807 VSS.n9806 185
R9114 VSS.n9728 VSS.n9667 185
R9115 VSS.n9810 VSS.n9667 185
R9116 VSS.t18 VSS.n9661 185
R9117 VSS.n9810 VSS.n9661 185
R9118 VSS.n9810 VSS.n9658 185
R9119 VSS.t18 VSS.n9658 185
R9120 VSS.t18 VSS.n9662 185
R9121 VSS.n9810 VSS.n9662 185
R9122 VSS.n9810 VSS.n9657 185
R9123 VSS.t18 VSS.n9657 185
R9124 VSS.t18 VSS.n9663 185
R9125 VSS.n9810 VSS.n9663 185
R9126 VSS.n9810 VSS.n9656 185
R9127 VSS.t18 VSS.n9656 185
R9128 VSS.t18 VSS.n9811 185
R9129 VSS.n9811 VSS.n9810 185
R9130 VSS.t38 VSS.n10323 185
R9131 VSS.n10314 VSS.n9181 185
R9132 VSS.n8936 VSS.n8935 185
R9133 VSS.n8941 VSS.n8935 185
R9134 VSS.n8947 VSS.n8935 185
R9135 VSS.n8953 VSS.n8935 185
R9136 VSS.n8958 VSS.n8935 185
R9137 VSS.n8965 VSS.n8935 185
R9138 VSS.t38 VSS.n8936 185
R9139 VSS.t38 VSS.n8941 185
R9140 VSS.t38 VSS.n8947 185
R9141 VSS.t38 VSS.n8953 185
R9142 VSS.t38 VSS.n8958 185
R9143 VSS.t38 VSS.n8965 185
R9144 VSS.t38 VSS.n8971 185
R9145 VSS.n10330 VSS.n10329 185
R9146 VSS.n10336 VSS.n10335 185
R9147 VSS.n10342 VSS.n10341 185
R9148 VSS.n10348 VSS.n10347 185
R9149 VSS.n10354 VSS.n10353 185
R9150 VSS.n10360 VSS.n10359 185
R9151 VSS.n10366 VSS.n10365 185
R9152 VSS.n9184 VSS.n9183 185
R9153 VSS.t46 VSS.n3624 185
R9154 VSS.n5739 VSS.n5738 185
R9155 VSS.n5745 VSS.n5744 185
R9156 VSS.n5751 VSS.n5750 185
R9157 VSS.n5757 VSS.n5756 185
R9158 VSS.n5763 VSS.n5762 185
R9159 VSS.n5769 VSS.n5768 185
R9160 VSS.n5775 VSS.n5774 185
R9161 VSS.n5781 VSS.n5780 185
R9162 VSS.n5669 VSS.n5668 185
R9163 VSS.n5669 VSS.n3582 185
R9164 VSS.t46 VSS.n3583 185
R9165 VSS.n3583 VSS.n3582 185
R9166 VSS.n3588 VSS.n3582 185
R9167 VSS.t46 VSS.n3588 185
R9168 VSS.t46 VSS.n3594 185
R9169 VSS.n3594 VSS.n3582 185
R9170 VSS.n3600 VSS.n3582 185
R9171 VSS.t46 VSS.n3600 185
R9172 VSS.t46 VSS.n3606 185
R9173 VSS.n3606 VSS.n3582 185
R9174 VSS.n3611 VSS.n3582 185
R9175 VSS.t46 VSS.n3611 185
R9176 VSS.t46 VSS.n3618 185
R9177 VSS.n3618 VSS.n3582 185
R9178 VSS.t70 VSS.n3566 185
R9179 VSS.n5861 VSS.n5860 185
R9180 VSS.n5867 VSS.n5866 185
R9181 VSS.n5873 VSS.n5872 185
R9182 VSS.n5879 VSS.n5878 185
R9183 VSS.n5885 VSS.n5884 185
R9184 VSS.n5891 VSS.n5890 185
R9185 VSS.n5897 VSS.n5896 185
R9186 VSS.n5903 VSS.n5902 185
R9187 VSS.n5791 VSS.n5790 185
R9188 VSS.n5791 VSS.n3524 185
R9189 VSS.t70 VSS.n3525 185
R9190 VSS.n3525 VSS.n3524 185
R9191 VSS.n3530 VSS.n3524 185
R9192 VSS.t70 VSS.n3530 185
R9193 VSS.t70 VSS.n3536 185
R9194 VSS.n3536 VSS.n3524 185
R9195 VSS.n3542 VSS.n3524 185
R9196 VSS.t70 VSS.n3542 185
R9197 VSS.t70 VSS.n3548 185
R9198 VSS.n3548 VSS.n3524 185
R9199 VSS.n3553 VSS.n3524 185
R9200 VSS.t70 VSS.n3553 185
R9201 VSS.t70 VSS.n3560 185
R9202 VSS.n3560 VSS.n3524 185
R9203 VSS.t66 VSS.n3508 185
R9204 VSS.n5983 VSS.n5982 185
R9205 VSS.n5989 VSS.n5988 185
R9206 VSS.n5995 VSS.n5994 185
R9207 VSS.n6001 VSS.n6000 185
R9208 VSS.n6007 VSS.n6006 185
R9209 VSS.n6013 VSS.n6012 185
R9210 VSS.n6019 VSS.n6018 185
R9211 VSS.n6025 VSS.n6024 185
R9212 VSS.n5913 VSS.n5912 185
R9213 VSS.n5913 VSS.n3466 185
R9214 VSS.t66 VSS.n3467 185
R9215 VSS.n3467 VSS.n3466 185
R9216 VSS.n3472 VSS.n3466 185
R9217 VSS.t66 VSS.n3472 185
R9218 VSS.t66 VSS.n3478 185
R9219 VSS.n3478 VSS.n3466 185
R9220 VSS.n3484 VSS.n3466 185
R9221 VSS.t66 VSS.n3484 185
R9222 VSS.t66 VSS.n3490 185
R9223 VSS.n3490 VSS.n3466 185
R9224 VSS.n3495 VSS.n3466 185
R9225 VSS.t66 VSS.n3495 185
R9226 VSS.t66 VSS.n3502 185
R9227 VSS.n3502 VSS.n3466 185
R9228 VSS.t64 VSS.n3450 185
R9229 VSS.n6105 VSS.n6104 185
R9230 VSS.n6111 VSS.n6110 185
R9231 VSS.n6117 VSS.n6116 185
R9232 VSS.n6123 VSS.n6122 185
R9233 VSS.n6129 VSS.n6128 185
R9234 VSS.n6135 VSS.n6134 185
R9235 VSS.n6141 VSS.n6140 185
R9236 VSS.n6147 VSS.n6146 185
R9237 VSS.n6035 VSS.n6034 185
R9238 VSS.n6035 VSS.n3408 185
R9239 VSS.t64 VSS.n3409 185
R9240 VSS.n3409 VSS.n3408 185
R9241 VSS.n3414 VSS.n3408 185
R9242 VSS.t64 VSS.n3414 185
R9243 VSS.t64 VSS.n3420 185
R9244 VSS.n3420 VSS.n3408 185
R9245 VSS.n3426 VSS.n3408 185
R9246 VSS.t64 VSS.n3426 185
R9247 VSS.t64 VSS.n3432 185
R9248 VSS.n3432 VSS.n3408 185
R9249 VSS.n3437 VSS.n3408 185
R9250 VSS.t64 VSS.n3437 185
R9251 VSS.t64 VSS.n3444 185
R9252 VSS.n3444 VSS.n3408 185
R9253 VSS.t84 VSS.n3392 185
R9254 VSS.n6227 VSS.n6226 185
R9255 VSS.n6233 VSS.n6232 185
R9256 VSS.n6239 VSS.n6238 185
R9257 VSS.n6245 VSS.n6244 185
R9258 VSS.n6251 VSS.n6250 185
R9259 VSS.n6257 VSS.n6256 185
R9260 VSS.n6263 VSS.n6262 185
R9261 VSS.n6269 VSS.n6268 185
R9262 VSS.n6157 VSS.n6156 185
R9263 VSS.n6157 VSS.n3350 185
R9264 VSS.t84 VSS.n3351 185
R9265 VSS.n3351 VSS.n3350 185
R9266 VSS.n3356 VSS.n3350 185
R9267 VSS.t84 VSS.n3356 185
R9268 VSS.t84 VSS.n3362 185
R9269 VSS.n3362 VSS.n3350 185
R9270 VSS.n3368 VSS.n3350 185
R9271 VSS.t84 VSS.n3368 185
R9272 VSS.t84 VSS.n3374 185
R9273 VSS.n3374 VSS.n3350 185
R9274 VSS.n3379 VSS.n3350 185
R9275 VSS.t84 VSS.n3379 185
R9276 VSS.t84 VSS.n3386 185
R9277 VSS.n3386 VSS.n3350 185
R9278 VSS.t86 VSS.n3334 185
R9279 VSS.n6349 VSS.n6348 185
R9280 VSS.n6355 VSS.n6354 185
R9281 VSS.n6361 VSS.n6360 185
R9282 VSS.n6367 VSS.n6366 185
R9283 VSS.n6373 VSS.n6372 185
R9284 VSS.n6379 VSS.n6378 185
R9285 VSS.n6385 VSS.n6384 185
R9286 VSS.n6391 VSS.n6390 185
R9287 VSS.n6279 VSS.n6278 185
R9288 VSS.n6279 VSS.n3292 185
R9289 VSS.t86 VSS.n3293 185
R9290 VSS.n3293 VSS.n3292 185
R9291 VSS.n3298 VSS.n3292 185
R9292 VSS.t86 VSS.n3298 185
R9293 VSS.t86 VSS.n3304 185
R9294 VSS.n3304 VSS.n3292 185
R9295 VSS.n3310 VSS.n3292 185
R9296 VSS.t86 VSS.n3310 185
R9297 VSS.t86 VSS.n3316 185
R9298 VSS.n3316 VSS.n3292 185
R9299 VSS.n3321 VSS.n3292 185
R9300 VSS.t86 VSS.n3321 185
R9301 VSS.t86 VSS.n3328 185
R9302 VSS.n3328 VSS.n3292 185
R9303 VSS.t24 VSS.n3276 185
R9304 VSS.n6471 VSS.n6470 185
R9305 VSS.n6477 VSS.n6476 185
R9306 VSS.n6483 VSS.n6482 185
R9307 VSS.n6489 VSS.n6488 185
R9308 VSS.n6495 VSS.n6494 185
R9309 VSS.n6501 VSS.n6500 185
R9310 VSS.n6507 VSS.n6506 185
R9311 VSS.n6513 VSS.n6512 185
R9312 VSS.n6401 VSS.n6400 185
R9313 VSS.n6401 VSS.n3234 185
R9314 VSS.t24 VSS.n3235 185
R9315 VSS.n3235 VSS.n3234 185
R9316 VSS.n3240 VSS.n3234 185
R9317 VSS.t24 VSS.n3240 185
R9318 VSS.t24 VSS.n3246 185
R9319 VSS.n3246 VSS.n3234 185
R9320 VSS.n3252 VSS.n3234 185
R9321 VSS.t24 VSS.n3252 185
R9322 VSS.t24 VSS.n3258 185
R9323 VSS.n3258 VSS.n3234 185
R9324 VSS.n3263 VSS.n3234 185
R9325 VSS.t24 VSS.n3263 185
R9326 VSS.t24 VSS.n3270 185
R9327 VSS.n3270 VSS.n3234 185
R9328 VSS.n3157 VSS.t44 185
R9329 VSS.n3226 VSS.n3225 185
R9330 VSS.n3218 VSS.n3217 185
R9331 VSS.n3210 VSS.n3209 185
R9332 VSS.n3202 VSS.n3201 185
R9333 VSS.n3194 VSS.n3193 185
R9334 VSS.n3186 VSS.n3185 185
R9335 VSS.n3178 VSS.n3177 185
R9336 VSS.n6601 VSS.n6600 185
R9337 VSS.n6537 VSS.n3149 185
R9338 VSS.n6598 VSS.n3149 185
R9339 VSS.n6599 VSS.t44 185
R9340 VSS.n6599 VSS.n6598 185
R9341 VSS.n6598 VSS.n3144 185
R9342 VSS.n3144 VSS.t44 185
R9343 VSS.n3146 VSS.t44 185
R9344 VSS.n6598 VSS.n3146 185
R9345 VSS.n6598 VSS.n3143 185
R9346 VSS.n3143 VSS.t44 185
R9347 VSS.n3147 VSS.t44 185
R9348 VSS.n6598 VSS.n3147 185
R9349 VSS.n6598 VSS.n3142 185
R9350 VSS.n3142 VSS.t44 185
R9351 VSS.n3148 VSS.t44 185
R9352 VSS.n6598 VSS.n3148 185
R9353 VSS.t60 VSS.n27 185
R9354 VSS.n1204 VSS.n1203 185
R9355 VSS.n1201 VSS.n31 185
R9356 VSS.n1198 VSS.n1197 185
R9357 VSS.n1194 VSS.n1193 185
R9358 VSS.n1190 VSS.n1189 185
R9359 VSS.n1187 VSS.n1186 185
R9360 VSS.n1241 VSS.n1240 185
R9361 VSS.n1250 VSS.n1249 185
R9362 VSS.n1176 VSS.n34 185
R9363 VSS.n1252 VSS.n34 185
R9364 VSS.t60 VSS.n28 185
R9365 VSS.n1252 VSS.n28 185
R9366 VSS.n1252 VSS.n25 185
R9367 VSS.t60 VSS.n25 185
R9368 VSS.t60 VSS.n29 185
R9369 VSS.n1252 VSS.n29 185
R9370 VSS.n1252 VSS.n24 185
R9371 VSS.t60 VSS.n24 185
R9372 VSS.t60 VSS.n30 185
R9373 VSS.n1252 VSS.n30 185
R9374 VSS.n1252 VSS.n23 185
R9375 VSS.t60 VSS.n23 185
R9376 VSS.t60 VSS.n1253 185
R9377 VSS.n1253 VSS.n1252 185
R9378 VSS.t48 VSS.n118 185
R9379 VSS.n1114 VSS.n1113 185
R9380 VSS.n1111 VSS.n122 185
R9381 VSS.n1108 VSS.n1107 185
R9382 VSS.n1104 VSS.n1103 185
R9383 VSS.n1100 VSS.n1099 185
R9384 VSS.n1097 VSS.n1096 185
R9385 VSS.n1156 VSS.n1155 185
R9386 VSS.n1165 VSS.n1164 185
R9387 VSS.n1086 VSS.n125 185
R9388 VSS.n1168 VSS.n125 185
R9389 VSS.t48 VSS.n119 185
R9390 VSS.n1168 VSS.n119 185
R9391 VSS.n1168 VSS.n116 185
R9392 VSS.t48 VSS.n116 185
R9393 VSS.t48 VSS.n120 185
R9394 VSS.n1168 VSS.n120 185
R9395 VSS.n1168 VSS.n115 185
R9396 VSS.t48 VSS.n115 185
R9397 VSS.t48 VSS.n121 185
R9398 VSS.n1168 VSS.n121 185
R9399 VSS.n1168 VSS.n114 185
R9400 VSS.t48 VSS.n114 185
R9401 VSS.t48 VSS.n1169 185
R9402 VSS.n1169 VSS.n1168 185
R9403 VSS.t76 VSS.n208 185
R9404 VSS.n1024 VSS.n1023 185
R9405 VSS.n1021 VSS.n212 185
R9406 VSS.n1018 VSS.n1017 185
R9407 VSS.n1014 VSS.n1013 185
R9408 VSS.n1010 VSS.n1009 185
R9409 VSS.n1007 VSS.n1006 185
R9410 VSS.n1066 VSS.n1065 185
R9411 VSS.n1075 VSS.n1074 185
R9412 VSS.n996 VSS.n215 185
R9413 VSS.n1078 VSS.n215 185
R9414 VSS.t76 VSS.n209 185
R9415 VSS.n1078 VSS.n209 185
R9416 VSS.n1078 VSS.n206 185
R9417 VSS.t76 VSS.n206 185
R9418 VSS.t76 VSS.n210 185
R9419 VSS.n1078 VSS.n210 185
R9420 VSS.n1078 VSS.n205 185
R9421 VSS.t76 VSS.n205 185
R9422 VSS.t76 VSS.n211 185
R9423 VSS.n1078 VSS.n211 185
R9424 VSS.n1078 VSS.n204 185
R9425 VSS.t76 VSS.n204 185
R9426 VSS.t76 VSS.n1079 185
R9427 VSS.n1079 VSS.n1078 185
R9428 VSS.t22 VSS.n298 185
R9429 VSS.n934 VSS.n933 185
R9430 VSS.n931 VSS.n302 185
R9431 VSS.n928 VSS.n927 185
R9432 VSS.n924 VSS.n923 185
R9433 VSS.n920 VSS.n919 185
R9434 VSS.n917 VSS.n916 185
R9435 VSS.n976 VSS.n975 185
R9436 VSS.n985 VSS.n984 185
R9437 VSS.n906 VSS.n305 185
R9438 VSS.n988 VSS.n305 185
R9439 VSS.t22 VSS.n299 185
R9440 VSS.n988 VSS.n299 185
R9441 VSS.n988 VSS.n296 185
R9442 VSS.t22 VSS.n296 185
R9443 VSS.t22 VSS.n300 185
R9444 VSS.n988 VSS.n300 185
R9445 VSS.n988 VSS.n295 185
R9446 VSS.t22 VSS.n295 185
R9447 VSS.t22 VSS.n301 185
R9448 VSS.n988 VSS.n301 185
R9449 VSS.n988 VSS.n294 185
R9450 VSS.t22 VSS.n294 185
R9451 VSS.t22 VSS.n989 185
R9452 VSS.n989 VSS.n988 185
R9453 VSS.t16 VSS.n388 185
R9454 VSS.n844 VSS.n843 185
R9455 VSS.n841 VSS.n392 185
R9456 VSS.n838 VSS.n837 185
R9457 VSS.n834 VSS.n833 185
R9458 VSS.n830 VSS.n829 185
R9459 VSS.n827 VSS.n826 185
R9460 VSS.n886 VSS.n885 185
R9461 VSS.n895 VSS.n894 185
R9462 VSS.n816 VSS.n395 185
R9463 VSS.n898 VSS.n395 185
R9464 VSS.t16 VSS.n389 185
R9465 VSS.n898 VSS.n389 185
R9466 VSS.n898 VSS.n386 185
R9467 VSS.t16 VSS.n386 185
R9468 VSS.t16 VSS.n390 185
R9469 VSS.n898 VSS.n390 185
R9470 VSS.n898 VSS.n385 185
R9471 VSS.t16 VSS.n385 185
R9472 VSS.t16 VSS.n391 185
R9473 VSS.n898 VSS.n391 185
R9474 VSS.n898 VSS.n384 185
R9475 VSS.t16 VSS.n384 185
R9476 VSS.t16 VSS.n899 185
R9477 VSS.n899 VSS.n898 185
R9478 VSS.t36 VSS.n478 185
R9479 VSS.n754 VSS.n753 185
R9480 VSS.n751 VSS.n482 185
R9481 VSS.n748 VSS.n747 185
R9482 VSS.n744 VSS.n743 185
R9483 VSS.n740 VSS.n739 185
R9484 VSS.n737 VSS.n736 185
R9485 VSS.n796 VSS.n795 185
R9486 VSS.n805 VSS.n804 185
R9487 VSS.n726 VSS.n485 185
R9488 VSS.n808 VSS.n485 185
R9489 VSS.t36 VSS.n479 185
R9490 VSS.n808 VSS.n479 185
R9491 VSS.n808 VSS.n476 185
R9492 VSS.t36 VSS.n476 185
R9493 VSS.t36 VSS.n480 185
R9494 VSS.n808 VSS.n480 185
R9495 VSS.n808 VSS.n475 185
R9496 VSS.t36 VSS.n475 185
R9497 VSS.t36 VSS.n481 185
R9498 VSS.n808 VSS.n481 185
R9499 VSS.n808 VSS.n474 185
R9500 VSS.t36 VSS.n474 185
R9501 VSS.t36 VSS.n809 185
R9502 VSS.n809 VSS.n808 185
R9503 VSS.t40 VSS.n568 185
R9504 VSS.n664 VSS.n663 185
R9505 VSS.n661 VSS.n572 185
R9506 VSS.n658 VSS.n657 185
R9507 VSS.n654 VSS.n653 185
R9508 VSS.n650 VSS.n649 185
R9509 VSS.n647 VSS.n646 185
R9510 VSS.n706 VSS.n705 185
R9511 VSS.n715 VSS.n714 185
R9512 VSS.n636 VSS.n575 185
R9513 VSS.n718 VSS.n575 185
R9514 VSS.t40 VSS.n569 185
R9515 VSS.n718 VSS.n569 185
R9516 VSS.n718 VSS.n566 185
R9517 VSS.t40 VSS.n566 185
R9518 VSS.t40 VSS.n570 185
R9519 VSS.n718 VSS.n570 185
R9520 VSS.n718 VSS.n565 185
R9521 VSS.t40 VSS.n565 185
R9522 VSS.t40 VSS.n571 185
R9523 VSS.n718 VSS.n571 185
R9524 VSS.n718 VSS.n564 185
R9525 VSS.t40 VSS.n564 185
R9526 VSS.t40 VSS.n719 185
R9527 VSS.n719 VSS.n718 185
R9528 VSS.n14723 VSS.n14363 181.396
R9529 VSS.n12794 VSS.n12723 181.396
R9530 VSS.n7837 VSS.n7672 181.396
R9531 VSS.n4247 VSS.n4176 181.396
R9532 VSS.n1964 VSS.n1604 181.396
R9533 VSS.n14727 VSS.n14361 175.544
R9534 VSS.n14731 VSS.n14361 175.544
R9535 VSS.n14731 VSS.n14359 175.544
R9536 VSS.n14735 VSS.n14359 175.544
R9537 VSS.n14735 VSS.n14357 175.544
R9538 VSS.n14739 VSS.n14357 175.544
R9539 VSS.n14739 VSS.n14355 175.544
R9540 VSS.n14743 VSS.n14355 175.544
R9541 VSS.n14743 VSS.n14353 175.544
R9542 VSS.n14747 VSS.n14353 175.544
R9543 VSS.n14747 VSS.n14351 175.544
R9544 VSS.n14782 VSS.n14334 175.544
R9545 VSS.n14782 VSS.n14332 175.544
R9546 VSS.n14786 VSS.n14332 175.544
R9547 VSS.n14786 VSS.n14330 175.544
R9548 VSS.n14790 VSS.n14330 175.544
R9549 VSS.n14790 VSS.n14328 175.544
R9550 VSS.n14794 VSS.n14328 175.544
R9551 VSS.n14794 VSS.n14326 175.544
R9552 VSS.n14798 VSS.n14326 175.544
R9553 VSS.n14798 VSS.n14323 175.544
R9554 VSS.n14837 VSS.n14323 175.544
R9555 VSS.n14751 VSS.n14349 175.544
R9556 VSS.n14755 VSS.n14349 175.544
R9557 VSS.n14755 VSS.n14347 175.544
R9558 VSS.n14759 VSS.n14347 175.544
R9559 VSS.n14759 VSS.n14345 175.544
R9560 VSS.n14763 VSS.n14345 175.544
R9561 VSS.n14763 VSS.n14343 175.544
R9562 VSS.n14768 VSS.n14343 175.544
R9563 VSS.n14768 VSS.n14341 175.544
R9564 VSS.n14772 VSS.n14341 175.544
R9565 VSS.n14773 VSS.n14772 175.544
R9566 VSS.n15361 VSS.n14220 175.544
R9567 VSS.n15365 VSS.n14220 175.544
R9568 VSS.n15365 VSS.n14218 175.544
R9569 VSS.n15369 VSS.n14218 175.544
R9570 VSS.n15369 VSS.n14216 175.544
R9571 VSS.n15373 VSS.n14216 175.544
R9572 VSS.n15373 VSS.n14214 175.544
R9573 VSS.n15378 VSS.n14214 175.544
R9574 VSS.n15378 VSS.n14212 175.544
R9575 VSS.n15382 VSS.n14212 175.544
R9576 VSS.n15383 VSS.n15382 175.544
R9577 VSS.n14833 VSS.n14832 175.544
R9578 VSS.n14832 VSS.n14802 175.544
R9579 VSS.n14828 VSS.n14802 175.544
R9580 VSS.n14828 VSS.n14804 175.544
R9581 VSS.n14824 VSS.n14804 175.544
R9582 VSS.n14824 VSS.n14807 175.544
R9583 VSS.n14820 VSS.n14807 175.544
R9584 VSS.n14820 VSS.n14809 175.544
R9585 VSS.n14816 VSS.n14809 175.544
R9586 VSS.n14816 VSS.n14813 175.544
R9587 VSS.n14813 VSS.n14812 175.544
R9588 VSS.n14192 VSS.n14160 175.544
R9589 VSS.n14188 VSS.n14160 175.544
R9590 VSS.n14188 VSS.n14162 175.544
R9591 VSS.n14184 VSS.n14162 175.544
R9592 VSS.n14184 VSS.n14164 175.544
R9593 VSS.n14180 VSS.n14164 175.544
R9594 VSS.n14180 VSS.n14166 175.544
R9595 VSS.n14176 VSS.n14166 175.544
R9596 VSS.n14176 VSS.n14168 175.544
R9597 VSS.n14172 VSS.n14168 175.544
R9598 VSS.n14172 VSS.n14170 175.544
R9599 VSS.n15392 VSS.n14205 175.544
R9600 VSS.n15392 VSS.n14203 175.544
R9601 VSS.n15396 VSS.n14203 175.544
R9602 VSS.n15396 VSS.n14201 175.544
R9603 VSS.n15400 VSS.n14201 175.544
R9604 VSS.n15400 VSS.n14199 175.544
R9605 VSS.n15404 VSS.n14199 175.544
R9606 VSS.n15404 VSS.n14197 175.544
R9607 VSS.n15408 VSS.n14197 175.544
R9608 VSS.n15408 VSS.n14195 175.544
R9609 VSS.n15412 VSS.n14195 175.544
R9610 VSS.n15921 VSS.n14053 175.544
R9611 VSS.n15925 VSS.n14053 175.544
R9612 VSS.n15925 VSS.n14051 175.544
R9613 VSS.n15929 VSS.n14051 175.544
R9614 VSS.n15929 VSS.n14049 175.544
R9615 VSS.n15933 VSS.n14049 175.544
R9616 VSS.n15933 VSS.n14047 175.544
R9617 VSS.n15938 VSS.n14047 175.544
R9618 VSS.n15938 VSS.n14045 175.544
R9619 VSS.n15942 VSS.n14045 175.544
R9620 VSS.n15943 VSS.n15942 175.544
R9621 VSS.n15952 VSS.n14038 175.544
R9622 VSS.n15952 VSS.n14036 175.544
R9623 VSS.n15956 VSS.n14036 175.544
R9624 VSS.n15956 VSS.n14034 175.544
R9625 VSS.n15960 VSS.n14034 175.544
R9626 VSS.n15960 VSS.n14032 175.544
R9627 VSS.n15964 VSS.n14032 175.544
R9628 VSS.n15964 VSS.n14030 175.544
R9629 VSS.n15968 VSS.n14030 175.544
R9630 VSS.n15968 VSS.n14028 175.544
R9631 VSS.n15972 VSS.n14028 175.544
R9632 VSS.n15996 VSS.n14016 175.544
R9633 VSS.n15992 VSS.n14016 175.544
R9634 VSS.n15992 VSS.n14018 175.544
R9635 VSS.n15988 VSS.n14018 175.544
R9636 VSS.n15988 VSS.n14020 175.544
R9637 VSS.n15984 VSS.n14020 175.544
R9638 VSS.n15984 VSS.n14022 175.544
R9639 VSS.n15980 VSS.n14022 175.544
R9640 VSS.n15980 VSS.n14024 175.544
R9641 VSS.n15976 VSS.n14024 175.544
R9642 VSS.n15976 VSS.n14026 175.544
R9643 VSS.n12788 VSS.n12787 175.544
R9644 VSS.n12787 VSS.n12726 175.544
R9645 VSS.n12783 VSS.n12726 175.544
R9646 VSS.n12783 VSS.n12728 175.544
R9647 VSS.n12779 VSS.n12728 175.544
R9648 VSS.n12779 VSS.n12731 175.544
R9649 VSS.n12775 VSS.n12731 175.544
R9650 VSS.n12775 VSS.n12733 175.544
R9651 VSS.n12771 VSS.n12733 175.544
R9652 VSS.n12771 VSS.n12735 175.544
R9653 VSS.n12767 VSS.n12735 175.544
R9654 VSS.n13099 VSS.n12640 175.544
R9655 VSS.n13099 VSS.n12638 175.544
R9656 VSS.n13103 VSS.n12638 175.544
R9657 VSS.n13103 VSS.n12636 175.544
R9658 VSS.n13107 VSS.n12636 175.544
R9659 VSS.n13107 VSS.n12634 175.544
R9660 VSS.n13111 VSS.n12634 175.544
R9661 VSS.n13111 VSS.n12632 175.544
R9662 VSS.n13115 VSS.n12632 175.544
R9663 VSS.n13115 VSS.n12630 175.544
R9664 VSS.n13119 VSS.n12630 175.544
R9665 VSS.n12763 VSS.n12737 175.544
R9666 VSS.n12763 VSS.n12739 175.544
R9667 VSS.n12759 VSS.n12739 175.544
R9668 VSS.n12759 VSS.n12741 175.544
R9669 VSS.n12755 VSS.n12741 175.544
R9670 VSS.n12755 VSS.n12743 175.544
R9671 VSS.n12751 VSS.n12743 175.544
R9672 VSS.n12751 VSS.n12745 175.544
R9673 VSS.n12747 VSS.n12745 175.544
R9674 VSS.n12747 VSS.n12643 175.544
R9675 VSS.n13094 VSS.n12643 175.544
R9676 VSS.n13348 VSS.n12499 175.544
R9677 VSS.n13348 VSS.n12497 175.544
R9678 VSS.n13352 VSS.n12497 175.544
R9679 VSS.n13352 VSS.n12495 175.544
R9680 VSS.n13356 VSS.n12495 175.544
R9681 VSS.n13356 VSS.n12493 175.544
R9682 VSS.n13360 VSS.n12493 175.544
R9683 VSS.n13360 VSS.n12491 175.544
R9684 VSS.n13364 VSS.n12491 175.544
R9685 VSS.n13364 VSS.n12489 175.544
R9686 VSS.n13368 VSS.n12489 175.544
R9687 VSS.n12627 VSS.n12600 175.544
R9688 VSS.n12623 VSS.n12600 175.544
R9689 VSS.n12623 VSS.n12602 175.544
R9690 VSS.n12619 VSS.n12602 175.544
R9691 VSS.n12619 VSS.n12604 175.544
R9692 VSS.n12615 VSS.n12604 175.544
R9693 VSS.n12615 VSS.n12606 175.544
R9694 VSS.n12611 VSS.n12606 175.544
R9695 VSS.n12611 VSS.n12608 175.544
R9696 VSS.n12608 VSS.n12502 175.544
R9697 VSS.n13343 VSS.n12502 175.544
R9698 VSS.n12457 VSS.n12456 175.544
R9699 VSS.n12456 VSS.n11516 175.544
R9700 VSS.n12452 VSS.n11516 175.544
R9701 VSS.n12452 VSS.n11518 175.544
R9702 VSS.n12448 VSS.n11518 175.544
R9703 VSS.n12448 VSS.n11521 175.544
R9704 VSS.n12444 VSS.n11521 175.544
R9705 VSS.n12444 VSS.n11523 175.544
R9706 VSS.n12440 VSS.n11523 175.544
R9707 VSS.n12440 VSS.n11525 175.544
R9708 VSS.n12436 VSS.n11525 175.544
R9709 VSS.n12486 VSS.n11499 175.544
R9710 VSS.n12482 VSS.n11499 175.544
R9711 VSS.n12482 VSS.n11501 175.544
R9712 VSS.n12478 VSS.n11501 175.544
R9713 VSS.n12478 VSS.n11503 175.544
R9714 VSS.n12474 VSS.n11503 175.544
R9715 VSS.n12474 VSS.n11505 175.544
R9716 VSS.n12470 VSS.n11505 175.544
R9717 VSS.n12470 VSS.n11507 175.544
R9718 VSS.n12466 VSS.n11507 175.544
R9719 VSS.n12466 VSS.n11509 175.544
R9720 VSS.n12137 VSS.n12136 175.544
R9721 VSS.n12140 VSS.n12137 175.544
R9722 VSS.n12140 VSS.n12133 175.544
R9723 VSS.n12144 VSS.n12133 175.544
R9724 VSS.n12144 VSS.n12131 175.544
R9725 VSS.n12148 VSS.n12131 175.544
R9726 VSS.n12148 VSS.n12129 175.544
R9727 VSS.n12153 VSS.n12129 175.544
R9728 VSS.n12153 VSS.n12127 175.544
R9729 VSS.n12157 VSS.n12127 175.544
R9730 VSS.n12158 VSS.n12157 175.544
R9731 VSS.n12167 VSS.n12087 175.544
R9732 VSS.n12167 VSS.n12085 175.544
R9733 VSS.n12171 VSS.n12085 175.544
R9734 VSS.n12171 VSS.n12083 175.544
R9735 VSS.n12175 VSS.n12083 175.544
R9736 VSS.n12175 VSS.n12081 175.544
R9737 VSS.n12179 VSS.n12081 175.544
R9738 VSS.n12179 VSS.n12079 175.544
R9739 VSS.n12183 VSS.n12079 175.544
R9740 VSS.n12183 VSS.n12077 175.544
R9741 VSS.n12187 VSS.n12077 175.544
R9742 VSS.n12211 VSS.n12065 175.544
R9743 VSS.n12207 VSS.n12065 175.544
R9744 VSS.n12207 VSS.n12067 175.544
R9745 VSS.n12203 VSS.n12067 175.544
R9746 VSS.n12203 VSS.n12069 175.544
R9747 VSS.n12199 VSS.n12069 175.544
R9748 VSS.n12199 VSS.n12071 175.544
R9749 VSS.n12195 VSS.n12071 175.544
R9750 VSS.n12195 VSS.n12073 175.544
R9751 VSS.n12191 VSS.n12073 175.544
R9752 VSS.n12191 VSS.n12075 175.544
R9753 VSS.n7844 VSS.n7670 175.544
R9754 VSS.n7844 VSS.n7668 175.544
R9755 VSS.n7848 VSS.n7668 175.544
R9756 VSS.n7848 VSS.n7666 175.544
R9757 VSS.n7852 VSS.n7666 175.544
R9758 VSS.n7852 VSS.n7664 175.544
R9759 VSS.n7856 VSS.n7664 175.544
R9760 VSS.n7856 VSS.n7662 175.544
R9761 VSS.n7860 VSS.n7662 175.544
R9762 VSS.n7860 VSS.n7660 175.544
R9763 VSS.n7864 VSS.n7660 175.544
R9764 VSS.n7645 VSS.n7618 175.544
R9765 VSS.n7641 VSS.n7618 175.544
R9766 VSS.n7641 VSS.n7620 175.544
R9767 VSS.n7637 VSS.n7620 175.544
R9768 VSS.n7637 VSS.n7622 175.544
R9769 VSS.n7633 VSS.n7622 175.544
R9770 VSS.n7633 VSS.n7624 175.544
R9771 VSS.n7629 VSS.n7624 175.544
R9772 VSS.n7629 VSS.n7626 175.544
R9773 VSS.n7626 VSS.n7521 175.544
R9774 VSS.n8221 VSS.n7521 175.544
R9775 VSS.n7868 VSS.n7658 175.544
R9776 VSS.n7868 VSS.n7656 175.544
R9777 VSS.n7872 VSS.n7656 175.544
R9778 VSS.n7872 VSS.n7654 175.544
R9779 VSS.n7876 VSS.n7654 175.544
R9780 VSS.n7876 VSS.n7652 175.544
R9781 VSS.n7880 VSS.n7652 175.544
R9782 VSS.n7880 VSS.n7650 175.544
R9783 VSS.n7884 VSS.n7650 175.544
R9784 VSS.n7884 VSS.n7648 175.544
R9785 VSS.n7888 VSS.n7648 175.544
R9786 VSS.n7505 VSS.n7478 175.544
R9787 VSS.n7501 VSS.n7478 175.544
R9788 VSS.n7501 VSS.n7480 175.544
R9789 VSS.n7497 VSS.n7480 175.544
R9790 VSS.n7497 VSS.n7482 175.544
R9791 VSS.n7493 VSS.n7482 175.544
R9792 VSS.n7493 VSS.n7484 175.544
R9793 VSS.n7489 VSS.n7484 175.544
R9794 VSS.n7489 VSS.n7486 175.544
R9795 VSS.n7486 VSS.n7381 175.544
R9796 VSS.n8579 VSS.n7381 175.544
R9797 VSS.n8226 VSS.n7518 175.544
R9798 VSS.n8226 VSS.n7516 175.544
R9799 VSS.n8230 VSS.n7516 175.544
R9800 VSS.n8230 VSS.n7514 175.544
R9801 VSS.n8234 VSS.n7514 175.544
R9802 VSS.n8234 VSS.n7512 175.544
R9803 VSS.n8238 VSS.n7512 175.544
R9804 VSS.n8238 VSS.n7510 175.544
R9805 VSS.n8242 VSS.n7510 175.544
R9806 VSS.n8242 VSS.n7508 175.544
R9807 VSS.n8246 VSS.n7508 175.544
R9808 VSS.n7365 VSS.n7338 175.544
R9809 VSS.n7361 VSS.n7338 175.544
R9810 VSS.n7361 VSS.n7340 175.544
R9811 VSS.n7357 VSS.n7340 175.544
R9812 VSS.n7357 VSS.n7342 175.544
R9813 VSS.n7353 VSS.n7342 175.544
R9814 VSS.n7353 VSS.n7344 175.544
R9815 VSS.n7349 VSS.n7344 175.544
R9816 VSS.n7349 VSS.n7346 175.544
R9817 VSS.n7346 VSS.n7241 175.544
R9818 VSS.n8801 VSS.n7241 175.544
R9819 VSS.n8584 VSS.n7378 175.544
R9820 VSS.n8584 VSS.n7376 175.544
R9821 VSS.n8588 VSS.n7376 175.544
R9822 VSS.n8588 VSS.n7374 175.544
R9823 VSS.n8592 VSS.n7374 175.544
R9824 VSS.n8592 VSS.n7372 175.544
R9825 VSS.n8596 VSS.n7372 175.544
R9826 VSS.n8596 VSS.n7370 175.544
R9827 VSS.n8600 VSS.n7370 175.544
R9828 VSS.n8600 VSS.n7368 175.544
R9829 VSS.n8604 VSS.n7368 175.544
R9830 VSS.n8806 VSS.n7238 175.544
R9831 VSS.n8806 VSS.n7236 175.544
R9832 VSS.n8810 VSS.n7236 175.544
R9833 VSS.n8810 VSS.n7234 175.544
R9834 VSS.n8814 VSS.n7234 175.544
R9835 VSS.n8814 VSS.n7232 175.544
R9836 VSS.n8818 VSS.n7232 175.544
R9837 VSS.n8818 VSS.n7230 175.544
R9838 VSS.n8822 VSS.n7230 175.544
R9839 VSS.n8822 VSS.n7228 175.544
R9840 VSS.n8826 VSS.n7228 175.544
R9841 VSS.n7225 VSS.n6982 175.544
R9842 VSS.n7221 VSS.n6982 175.544
R9843 VSS.n7221 VSS.n6984 175.544
R9844 VSS.n7217 VSS.n6984 175.544
R9845 VSS.n7217 VSS.n6986 175.544
R9846 VSS.n7213 VSS.n6986 175.544
R9847 VSS.n7213 VSS.n6988 175.544
R9848 VSS.n7209 VSS.n6988 175.544
R9849 VSS.n7209 VSS.n6990 175.544
R9850 VSS.n7205 VSS.n6990 175.544
R9851 VSS.n7205 VSS.n6992 175.544
R9852 VSS.n7181 VSS.n7004 175.544
R9853 VSS.n7181 VSS.n7002 175.544
R9854 VSS.n7185 VSS.n7002 175.544
R9855 VSS.n7185 VSS.n7000 175.544
R9856 VSS.n7189 VSS.n7000 175.544
R9857 VSS.n7189 VSS.n6998 175.544
R9858 VSS.n7193 VSS.n6998 175.544
R9859 VSS.n7193 VSS.n6996 175.544
R9860 VSS.n7197 VSS.n6996 175.544
R9861 VSS.n7197 VSS.n6994 175.544
R9862 VSS.n7201 VSS.n6994 175.544
R9863 VSS.n6798 VSS.n6772 175.544
R9864 VSS.n6798 VSS.n6774 175.544
R9865 VSS.n6794 VSS.n6774 175.544
R9866 VSS.n6794 VSS.n6776 175.544
R9867 VSS.n6790 VSS.n6776 175.544
R9868 VSS.n6790 VSS.n6778 175.544
R9869 VSS.n6786 VSS.n6778 175.544
R9870 VSS.n6786 VSS.n6780 175.544
R9871 VSS.n6782 VSS.n6780 175.544
R9872 VSS.n6782 VSS.n6731 175.544
R9873 VSS.n6878 VSS.n6731 175.544
R9874 VSS.n6854 VSS.n6743 175.544
R9875 VSS.n6858 VSS.n6743 175.544
R9876 VSS.n6858 VSS.n6741 175.544
R9877 VSS.n6862 VSS.n6741 175.544
R9878 VSS.n6862 VSS.n6739 175.544
R9879 VSS.n6866 VSS.n6739 175.544
R9880 VSS.n6866 VSS.n6737 175.544
R9881 VSS.n6870 VSS.n6737 175.544
R9882 VSS.n6870 VSS.n6735 175.544
R9883 VSS.n6874 VSS.n6735 175.544
R9884 VSS.n6874 VSS.n6732 175.544
R9885 VSS.n6830 VSS.n6755 175.544
R9886 VSS.n6834 VSS.n6755 175.544
R9887 VSS.n6834 VSS.n6753 175.544
R9888 VSS.n6838 VSS.n6753 175.544
R9889 VSS.n6838 VSS.n6751 175.544
R9890 VSS.n6842 VSS.n6751 175.544
R9891 VSS.n6842 VSS.n6749 175.544
R9892 VSS.n6846 VSS.n6749 175.544
R9893 VSS.n6846 VSS.n6747 175.544
R9894 VSS.n6850 VSS.n6747 175.544
R9895 VSS.n6850 VSS.n6745 175.544
R9896 VSS.n6826 VSS.n6760 175.544
R9897 VSS.n6822 VSS.n6760 175.544
R9898 VSS.n6822 VSS.n6762 175.544
R9899 VSS.n6818 VSS.n6762 175.544
R9900 VSS.n6818 VSS.n6764 175.544
R9901 VSS.n6814 VSS.n6764 175.544
R9902 VSS.n6814 VSS.n6765 175.544
R9903 VSS.n6810 VSS.n6765 175.544
R9904 VSS.n6810 VSS.n6767 175.544
R9905 VSS.n6806 VSS.n6767 175.544
R9906 VSS.n6806 VSS.n6770 175.544
R9907 VSS.n4241 VSS.n4240 175.544
R9908 VSS.n4240 VSS.n4179 175.544
R9909 VSS.n4236 VSS.n4179 175.544
R9910 VSS.n4236 VSS.n4181 175.544
R9911 VSS.n4232 VSS.n4181 175.544
R9912 VSS.n4232 VSS.n4184 175.544
R9913 VSS.n4228 VSS.n4184 175.544
R9914 VSS.n4228 VSS.n4186 175.544
R9915 VSS.n4224 VSS.n4186 175.544
R9916 VSS.n4224 VSS.n4188 175.544
R9917 VSS.n4220 VSS.n4188 175.544
R9918 VSS.n4552 VSS.n4093 175.544
R9919 VSS.n4552 VSS.n4091 175.544
R9920 VSS.n4556 VSS.n4091 175.544
R9921 VSS.n4556 VSS.n4089 175.544
R9922 VSS.n4560 VSS.n4089 175.544
R9923 VSS.n4560 VSS.n4087 175.544
R9924 VSS.n4564 VSS.n4087 175.544
R9925 VSS.n4564 VSS.n4085 175.544
R9926 VSS.n4568 VSS.n4085 175.544
R9927 VSS.n4568 VSS.n4083 175.544
R9928 VSS.n4572 VSS.n4083 175.544
R9929 VSS.n4216 VSS.n4190 175.544
R9930 VSS.n4216 VSS.n4192 175.544
R9931 VSS.n4212 VSS.n4192 175.544
R9932 VSS.n4212 VSS.n4194 175.544
R9933 VSS.n4208 VSS.n4194 175.544
R9934 VSS.n4208 VSS.n4196 175.544
R9935 VSS.n4204 VSS.n4196 175.544
R9936 VSS.n4204 VSS.n4198 175.544
R9937 VSS.n4200 VSS.n4198 175.544
R9938 VSS.n4200 VSS.n4096 175.544
R9939 VSS.n4547 VSS.n4096 175.544
R9940 VSS.n4909 VSS.n3952 175.544
R9941 VSS.n4909 VSS.n3950 175.544
R9942 VSS.n4913 VSS.n3950 175.544
R9943 VSS.n4913 VSS.n3948 175.544
R9944 VSS.n4917 VSS.n3948 175.544
R9945 VSS.n4917 VSS.n3946 175.544
R9946 VSS.n4921 VSS.n3946 175.544
R9947 VSS.n4921 VSS.n3944 175.544
R9948 VSS.n4925 VSS.n3944 175.544
R9949 VSS.n4925 VSS.n3942 175.544
R9950 VSS.n4929 VSS.n3942 175.544
R9951 VSS.n4080 VSS.n4053 175.544
R9952 VSS.n4076 VSS.n4053 175.544
R9953 VSS.n4076 VSS.n4055 175.544
R9954 VSS.n4072 VSS.n4055 175.544
R9955 VSS.n4072 VSS.n4057 175.544
R9956 VSS.n4068 VSS.n4057 175.544
R9957 VSS.n4068 VSS.n4059 175.544
R9958 VSS.n4064 VSS.n4059 175.544
R9959 VSS.n4064 VSS.n4061 175.544
R9960 VSS.n4061 VSS.n3955 175.544
R9961 VSS.n4904 VSS.n3955 175.544
R9962 VSS.n5266 VSS.n3811 175.544
R9963 VSS.n5266 VSS.n3809 175.544
R9964 VSS.n5270 VSS.n3809 175.544
R9965 VSS.n5270 VSS.n3807 175.544
R9966 VSS.n5274 VSS.n3807 175.544
R9967 VSS.n5274 VSS.n3805 175.544
R9968 VSS.n5278 VSS.n3805 175.544
R9969 VSS.n5278 VSS.n3803 175.544
R9970 VSS.n5282 VSS.n3803 175.544
R9971 VSS.n5282 VSS.n3801 175.544
R9972 VSS.n5286 VSS.n3801 175.544
R9973 VSS.n3939 VSS.n3912 175.544
R9974 VSS.n3935 VSS.n3912 175.544
R9975 VSS.n3935 VSS.n3914 175.544
R9976 VSS.n3931 VSS.n3914 175.544
R9977 VSS.n3931 VSS.n3916 175.544
R9978 VSS.n3927 VSS.n3916 175.544
R9979 VSS.n3927 VSS.n3918 175.544
R9980 VSS.n3923 VSS.n3918 175.544
R9981 VSS.n3923 VSS.n3920 175.544
R9982 VSS.n3920 VSS.n3814 175.544
R9983 VSS.n5261 VSS.n3814 175.544
R9984 VSS.n3798 VSS.n3771 175.544
R9985 VSS.n3794 VSS.n3771 175.544
R9986 VSS.n3794 VSS.n3773 175.544
R9987 VSS.n3790 VSS.n3773 175.544
R9988 VSS.n3790 VSS.n3775 175.544
R9989 VSS.n3786 VSS.n3775 175.544
R9990 VSS.n3786 VSS.n3777 175.544
R9991 VSS.n3782 VSS.n3777 175.544
R9992 VSS.n3782 VSS.n3779 175.544
R9993 VSS.n3779 VSS.n3673 175.544
R9994 VSS.n5607 VSS.n3673 175.544
R9995 VSS.n5612 VSS.n3670 175.544
R9996 VSS.n5612 VSS.n3668 175.544
R9997 VSS.n5616 VSS.n3668 175.544
R9998 VSS.n5616 VSS.n3666 175.544
R9999 VSS.n5620 VSS.n3666 175.544
R10000 VSS.n5620 VSS.n3664 175.544
R10001 VSS.n5624 VSS.n3664 175.544
R10002 VSS.n5624 VSS.n3662 175.544
R10003 VSS.n5628 VSS.n3662 175.544
R10004 VSS.n5628 VSS.n3660 175.544
R10005 VSS.n5632 VSS.n3660 175.544
R10006 VSS.n5656 VSS.n3643 175.544
R10007 VSS.n5652 VSS.n3643 175.544
R10008 VSS.n5652 VSS.n3650 175.544
R10009 VSS.n5648 VSS.n3650 175.544
R10010 VSS.n5648 VSS.n3652 175.544
R10011 VSS.n5644 VSS.n3652 175.544
R10012 VSS.n5644 VSS.n3654 175.544
R10013 VSS.n5640 VSS.n3654 175.544
R10014 VSS.n5640 VSS.n3656 175.544
R10015 VSS.n5636 VSS.n3656 175.544
R10016 VSS.n5636 VSS.n3658 175.544
R10017 VSS.n1968 VSS.n1602 175.544
R10018 VSS.n1972 VSS.n1602 175.544
R10019 VSS.n1972 VSS.n1600 175.544
R10020 VSS.n1976 VSS.n1600 175.544
R10021 VSS.n1976 VSS.n1598 175.544
R10022 VSS.n1980 VSS.n1598 175.544
R10023 VSS.n1980 VSS.n1596 175.544
R10024 VSS.n1984 VSS.n1596 175.544
R10025 VSS.n1984 VSS.n1594 175.544
R10026 VSS.n1988 VSS.n1594 175.544
R10027 VSS.n1988 VSS.n1592 175.544
R10028 VSS.n2023 VSS.n1575 175.544
R10029 VSS.n2023 VSS.n1573 175.544
R10030 VSS.n2027 VSS.n1573 175.544
R10031 VSS.n2027 VSS.n1571 175.544
R10032 VSS.n2031 VSS.n1571 175.544
R10033 VSS.n2031 VSS.n1569 175.544
R10034 VSS.n2035 VSS.n1569 175.544
R10035 VSS.n2035 VSS.n1567 175.544
R10036 VSS.n2039 VSS.n1567 175.544
R10037 VSS.n2039 VSS.n1564 175.544
R10038 VSS.n2078 VSS.n1564 175.544
R10039 VSS.n1992 VSS.n1590 175.544
R10040 VSS.n1996 VSS.n1590 175.544
R10041 VSS.n1996 VSS.n1588 175.544
R10042 VSS.n2000 VSS.n1588 175.544
R10043 VSS.n2000 VSS.n1586 175.544
R10044 VSS.n2004 VSS.n1586 175.544
R10045 VSS.n2004 VSS.n1584 175.544
R10046 VSS.n2009 VSS.n1584 175.544
R10047 VSS.n2009 VSS.n1582 175.544
R10048 VSS.n2013 VSS.n1582 175.544
R10049 VSS.n2014 VSS.n2013 175.544
R10050 VSS.n2602 VSS.n1461 175.544
R10051 VSS.n2606 VSS.n1461 175.544
R10052 VSS.n2606 VSS.n1459 175.544
R10053 VSS.n2610 VSS.n1459 175.544
R10054 VSS.n2610 VSS.n1457 175.544
R10055 VSS.n2614 VSS.n1457 175.544
R10056 VSS.n2614 VSS.n1455 175.544
R10057 VSS.n2619 VSS.n1455 175.544
R10058 VSS.n2619 VSS.n1453 175.544
R10059 VSS.n2623 VSS.n1453 175.544
R10060 VSS.n2624 VSS.n2623 175.544
R10061 VSS.n2074 VSS.n2073 175.544
R10062 VSS.n2073 VSS.n2043 175.544
R10063 VSS.n2069 VSS.n2043 175.544
R10064 VSS.n2069 VSS.n2045 175.544
R10065 VSS.n2065 VSS.n2045 175.544
R10066 VSS.n2065 VSS.n2048 175.544
R10067 VSS.n2061 VSS.n2048 175.544
R10068 VSS.n2061 VSS.n2050 175.544
R10069 VSS.n2057 VSS.n2050 175.544
R10070 VSS.n2057 VSS.n2054 175.544
R10071 VSS.n2054 VSS.n2053 175.544
R10072 VSS.n1433 VSS.n1401 175.544
R10073 VSS.n1429 VSS.n1401 175.544
R10074 VSS.n1429 VSS.n1403 175.544
R10075 VSS.n1425 VSS.n1403 175.544
R10076 VSS.n1425 VSS.n1405 175.544
R10077 VSS.n1421 VSS.n1405 175.544
R10078 VSS.n1421 VSS.n1407 175.544
R10079 VSS.n1417 VSS.n1407 175.544
R10080 VSS.n1417 VSS.n1409 175.544
R10081 VSS.n1413 VSS.n1409 175.544
R10082 VSS.n1413 VSS.n1411 175.544
R10083 VSS.n2633 VSS.n1446 175.544
R10084 VSS.n2633 VSS.n1444 175.544
R10085 VSS.n2637 VSS.n1444 175.544
R10086 VSS.n2637 VSS.n1442 175.544
R10087 VSS.n2641 VSS.n1442 175.544
R10088 VSS.n2641 VSS.n1440 175.544
R10089 VSS.n2645 VSS.n1440 175.544
R10090 VSS.n2645 VSS.n1438 175.544
R10091 VSS.n2649 VSS.n1438 175.544
R10092 VSS.n2649 VSS.n1436 175.544
R10093 VSS.n2653 VSS.n1436 175.544
R10094 VSS.n3039 VSS.n1271 175.544
R10095 VSS.n3039 VSS.n1274 175.544
R10096 VSS.n3035 VSS.n1274 175.544
R10097 VSS.n3035 VSS.n1276 175.544
R10098 VSS.n3031 VSS.n1276 175.544
R10099 VSS.n3031 VSS.n1278 175.544
R10100 VSS.n3027 VSS.n1278 175.544
R10101 VSS.n3027 VSS.n1280 175.544
R10102 VSS.n3023 VSS.n1280 175.544
R10103 VSS.n3023 VSS.n1282 175.544
R10104 VSS.n3019 VSS.n1282 175.544
R10105 VSS.n2995 VSS.n1294 175.544
R10106 VSS.n2999 VSS.n1294 175.544
R10107 VSS.n2999 VSS.n1292 175.544
R10108 VSS.n3003 VSS.n1292 175.544
R10109 VSS.n3003 VSS.n1290 175.544
R10110 VSS.n3007 VSS.n1290 175.544
R10111 VSS.n3007 VSS.n1288 175.544
R10112 VSS.n3011 VSS.n1288 175.544
R10113 VSS.n3011 VSS.n1286 175.544
R10114 VSS.n3015 VSS.n1286 175.544
R10115 VSS.n3015 VSS.n1284 175.544
R10116 VSS.n16004 VSS.n14012 167.742
R10117 VSS.n12219 VSS.n12061 167.742
R10118 VSS.n7172 VSS.n7010 167.742
R10119 VSS.n5660 VSS.n3640 167.742
R10120 VSS.n3043 VSS.n1270 167.742
R10121 VSS.n17327 VSS.n17313 151.666
R10122 VSS.n16082 VSS.n16057 151.666
R10123 VSS.n16172 VSS.n16147 151.666
R10124 VSS.n16262 VSS.n16237 151.666
R10125 VSS.n16352 VSS.n16327 151.666
R10126 VSS.n16442 VSS.n16417 151.666
R10127 VSS.n16532 VSS.n16507 151.666
R10128 VSS.n16622 VSS.n16597 151.666
R10129 VSS.n11150 VSS.n11064 151.666
R10130 VSS.n11240 VSS.n10974 151.666
R10131 VSS.n11330 VSS.n10884 151.666
R10132 VSS.n11420 VSS.n10794 151.666
R10133 VSS.n13540 VSS.n10704 151.666
R10134 VSS.n13630 VSS.n10614 151.666
R10135 VSS.n13720 VSS.n10524 151.666
R10136 VSS.n13824 VSS.n13810 151.666
R10137 VSS.n9157 VSS.n8984 151.666
R10138 VSS.n9217 VSS.n9192 151.666
R10139 VSS.n9307 VSS.n9282 151.666
R10140 VSS.n9397 VSS.n9372 151.666
R10141 VSS.n9487 VSS.n9462 151.666
R10142 VSS.n9577 VSS.n9552 151.666
R10143 VSS.n9667 VSS.n9642 151.666
R10144 VSS.n10315 VSS.n10314 151.666
R10145 VSS.n5670 VSS.n5669 151.666
R10146 VSS.n5792 VSS.n5791 151.666
R10147 VSS.n5914 VSS.n5913 151.666
R10148 VSS.n6036 VSS.n6035 151.666
R10149 VSS.n6158 VSS.n6157 151.666
R10150 VSS.n6280 VSS.n6279 151.666
R10151 VSS.n6402 VSS.n6401 151.666
R10152 VSS.n6540 VSS.n3149 151.666
R10153 VSS.n34 VSS.n9 151.666
R10154 VSS.n125 VSS.n100 151.666
R10155 VSS.n215 VSS.n190 151.666
R10156 VSS.n305 VSS.n280 151.666
R10157 VSS.n395 VSS.n370 151.666
R10158 VSS.n485 VSS.n460 151.666
R10159 VSS.n575 VSS.n550 151.666
R10160 VSS.n17383 VSS.n17313 150
R10161 VSS.n17379 VSS.n17326 150
R10162 VSS.n17377 VSS.n17376 150
R10163 VSS.n17373 VSS.n17372 150
R10164 VSS.n17365 VSS.n17364 150
R10165 VSS.n17361 VSS.n17360 150
R10166 VSS.n17357 VSS.n17356 150
R10167 VSS.n17353 VSS.n17321 150
R10168 VSS.n17336 VSS.n16030 150
R10169 VSS.n17340 VSS.n17339 150
R10170 VSS.n17344 VSS.n17343 150
R10171 VSS.n17348 VSS.n17347 150
R10172 VSS.n16139 VSS.n16057 150
R10173 VSS.n16137 VSS.n16136 150
R10174 VSS.n16133 VSS.n16132 150
R10175 VSS.n16129 VSS.n16128 150
R10176 VSS.n16121 VSS.n16120 150
R10177 VSS.n16117 VSS.n16116 150
R10178 VSS.n16113 VSS.n16112 150
R10179 VSS.n16109 VSS.n16065 150
R10180 VSS.n17307 VSS.n16056 150
R10181 VSS.n16096 VSS.n16095 150
R10182 VSS.n16100 VSS.n16099 150
R10183 VSS.n16104 VSS.n16103 150
R10184 VSS.n16229 VSS.n16147 150
R10185 VSS.n16227 VSS.n16226 150
R10186 VSS.n16223 VSS.n16222 150
R10187 VSS.n16219 VSS.n16218 150
R10188 VSS.n16211 VSS.n16210 150
R10189 VSS.n16207 VSS.n16206 150
R10190 VSS.n16203 VSS.n16202 150
R10191 VSS.n16199 VSS.n16155 150
R10192 VSS.n17217 VSS.n16146 150
R10193 VSS.n16186 VSS.n16185 150
R10194 VSS.n16190 VSS.n16189 150
R10195 VSS.n16194 VSS.n16193 150
R10196 VSS.n16319 VSS.n16237 150
R10197 VSS.n16317 VSS.n16316 150
R10198 VSS.n16313 VSS.n16312 150
R10199 VSS.n16309 VSS.n16308 150
R10200 VSS.n16301 VSS.n16300 150
R10201 VSS.n16297 VSS.n16296 150
R10202 VSS.n16293 VSS.n16292 150
R10203 VSS.n16289 VSS.n16245 150
R10204 VSS.n17127 VSS.n16236 150
R10205 VSS.n16276 VSS.n16275 150
R10206 VSS.n16280 VSS.n16279 150
R10207 VSS.n16284 VSS.n16283 150
R10208 VSS.n16409 VSS.n16327 150
R10209 VSS.n16407 VSS.n16406 150
R10210 VSS.n16403 VSS.n16402 150
R10211 VSS.n16399 VSS.n16398 150
R10212 VSS.n16391 VSS.n16390 150
R10213 VSS.n16387 VSS.n16386 150
R10214 VSS.n16383 VSS.n16382 150
R10215 VSS.n16379 VSS.n16335 150
R10216 VSS.n17037 VSS.n16326 150
R10217 VSS.n16366 VSS.n16365 150
R10218 VSS.n16370 VSS.n16369 150
R10219 VSS.n16374 VSS.n16373 150
R10220 VSS.n16499 VSS.n16417 150
R10221 VSS.n16497 VSS.n16496 150
R10222 VSS.n16493 VSS.n16492 150
R10223 VSS.n16489 VSS.n16488 150
R10224 VSS.n16481 VSS.n16480 150
R10225 VSS.n16477 VSS.n16476 150
R10226 VSS.n16473 VSS.n16472 150
R10227 VSS.n16469 VSS.n16425 150
R10228 VSS.n16947 VSS.n16416 150
R10229 VSS.n16456 VSS.n16455 150
R10230 VSS.n16460 VSS.n16459 150
R10231 VSS.n16464 VSS.n16463 150
R10232 VSS.n16589 VSS.n16507 150
R10233 VSS.n16587 VSS.n16586 150
R10234 VSS.n16583 VSS.n16582 150
R10235 VSS.n16579 VSS.n16578 150
R10236 VSS.n16571 VSS.n16570 150
R10237 VSS.n16567 VSS.n16566 150
R10238 VSS.n16563 VSS.n16562 150
R10239 VSS.n16559 VSS.n16515 150
R10240 VSS.n16857 VSS.n16506 150
R10241 VSS.n16546 VSS.n16545 150
R10242 VSS.n16550 VSS.n16549 150
R10243 VSS.n16554 VSS.n16553 150
R10244 VSS.n16679 VSS.n16597 150
R10245 VSS.n16677 VSS.n16676 150
R10246 VSS.n16673 VSS.n16672 150
R10247 VSS.n16669 VSS.n16668 150
R10248 VSS.n16661 VSS.n16660 150
R10249 VSS.n16657 VSS.n16656 150
R10250 VSS.n16653 VSS.n16652 150
R10251 VSS.n16649 VSS.n16605 150
R10252 VSS.n16767 VSS.n16596 150
R10253 VSS.n16636 VSS.n16635 150
R10254 VSS.n16640 VSS.n16639 150
R10255 VSS.n16644 VSS.n16643 150
R10256 VSS.n11146 VSS.n11064 150
R10257 VSS.n11144 VSS.n11143 150
R10258 VSS.n11140 VSS.n11139 150
R10259 VSS.n11136 VSS.n11135 150
R10260 VSS.n11128 VSS.n11127 150
R10261 VSS.n11124 VSS.n11123 150
R10262 VSS.n11120 VSS.n11119 150
R10263 VSS.n11116 VSS.n11072 150
R10264 VSS.n11234 VSS.n11063 150
R10265 VSS.n11103 VSS.n11102 150
R10266 VSS.n11107 VSS.n11106 150
R10267 VSS.n11111 VSS.n11110 150
R10268 VSS.n11056 VSS.n10974 150
R10269 VSS.n11054 VSS.n11053 150
R10270 VSS.n11050 VSS.n11049 150
R10271 VSS.n11046 VSS.n11045 150
R10272 VSS.n11038 VSS.n11037 150
R10273 VSS.n11034 VSS.n11033 150
R10274 VSS.n11030 VSS.n11029 150
R10275 VSS.n11026 VSS.n10982 150
R10276 VSS.n11324 VSS.n10973 150
R10277 VSS.n11013 VSS.n11012 150
R10278 VSS.n11017 VSS.n11016 150
R10279 VSS.n11021 VSS.n11020 150
R10280 VSS.n10966 VSS.n10884 150
R10281 VSS.n10964 VSS.n10963 150
R10282 VSS.n10960 VSS.n10959 150
R10283 VSS.n10956 VSS.n10955 150
R10284 VSS.n10948 VSS.n10947 150
R10285 VSS.n10944 VSS.n10943 150
R10286 VSS.n10940 VSS.n10939 150
R10287 VSS.n10936 VSS.n10892 150
R10288 VSS.n11414 VSS.n10883 150
R10289 VSS.n10923 VSS.n10922 150
R10290 VSS.n10927 VSS.n10926 150
R10291 VSS.n10931 VSS.n10930 150
R10292 VSS.n10876 VSS.n10794 150
R10293 VSS.n10874 VSS.n10873 150
R10294 VSS.n10870 VSS.n10869 150
R10295 VSS.n10866 VSS.n10865 150
R10296 VSS.n10858 VSS.n10857 150
R10297 VSS.n10854 VSS.n10853 150
R10298 VSS.n10850 VSS.n10849 150
R10299 VSS.n10846 VSS.n10802 150
R10300 VSS.n13534 VSS.n10793 150
R10301 VSS.n10833 VSS.n10832 150
R10302 VSS.n10837 VSS.n10836 150
R10303 VSS.n10841 VSS.n10840 150
R10304 VSS.n10786 VSS.n10704 150
R10305 VSS.n10784 VSS.n10783 150
R10306 VSS.n10780 VSS.n10779 150
R10307 VSS.n10776 VSS.n10775 150
R10308 VSS.n10768 VSS.n10767 150
R10309 VSS.n10764 VSS.n10763 150
R10310 VSS.n10760 VSS.n10759 150
R10311 VSS.n10756 VSS.n10712 150
R10312 VSS.n13624 VSS.n10703 150
R10313 VSS.n10743 VSS.n10742 150
R10314 VSS.n10747 VSS.n10746 150
R10315 VSS.n10751 VSS.n10750 150
R10316 VSS.n10696 VSS.n10614 150
R10317 VSS.n10694 VSS.n10693 150
R10318 VSS.n10690 VSS.n10689 150
R10319 VSS.n10686 VSS.n10685 150
R10320 VSS.n10678 VSS.n10677 150
R10321 VSS.n10674 VSS.n10673 150
R10322 VSS.n10670 VSS.n10669 150
R10323 VSS.n10666 VSS.n10622 150
R10324 VSS.n13714 VSS.n10613 150
R10325 VSS.n10653 VSS.n10652 150
R10326 VSS.n10657 VSS.n10656 150
R10327 VSS.n10661 VSS.n10660 150
R10328 VSS.n10606 VSS.n10524 150
R10329 VSS.n10604 VSS.n10603 150
R10330 VSS.n10600 VSS.n10599 150
R10331 VSS.n10596 VSS.n10595 150
R10332 VSS.n10588 VSS.n10587 150
R10333 VSS.n10584 VSS.n10583 150
R10334 VSS.n10580 VSS.n10579 150
R10335 VSS.n10576 VSS.n10532 150
R10336 VSS.n13804 VSS.n10523 150
R10337 VSS.n10563 VSS.n10562 150
R10338 VSS.n10567 VSS.n10566 150
R10339 VSS.n10571 VSS.n10570 150
R10340 VSS.n13883 VSS.n13810 150
R10341 VSS.n13879 VSS.n13823 150
R10342 VSS.n13877 VSS.n13876 150
R10343 VSS.n13873 VSS.n13872 150
R10344 VSS.n13865 VSS.n13864 150
R10345 VSS.n13861 VSS.n13860 150
R10346 VSS.n13857 VSS.n13856 150
R10347 VSS.n13853 VSS.n13818 150
R10348 VSS.n13836 VSS.n10497 150
R10349 VSS.n13840 VSS.n13839 150
R10350 VSS.n13844 VSS.n13843 150
R10351 VSS.n13848 VSS.n13847 150
R10352 VSS.n9100 VSS.n9099 150
R10353 VSS.n9104 VSS.n9103 150
R10354 VSS.n9108 VSS.n9107 150
R10355 VSS.n9110 VSS.n8993 150
R10356 VSS.n9117 VSS.n9116 150
R10357 VSS.n9121 VSS.n9120 150
R10358 VSS.n9125 VSS.n9124 150
R10359 VSS.n9129 VSS.n9128 150
R10360 VSS.n9145 VSS.n9144 150
R10361 VSS.n9141 VSS.n9140 150
R10362 VSS.n9137 VSS.n9136 150
R10363 VSS.n9133 VSS.n9132 150
R10364 VSS.n9274 VSS.n9192 150
R10365 VSS.n9272 VSS.n9271 150
R10366 VSS.n9268 VSS.n9267 150
R10367 VSS.n9264 VSS.n9263 150
R10368 VSS.n9256 VSS.n9255 150
R10369 VSS.n9252 VSS.n9251 150
R10370 VSS.n9248 VSS.n9247 150
R10371 VSS.n9244 VSS.n9200 150
R10372 VSS.n10262 VSS.n9191 150
R10373 VSS.n9231 VSS.n9230 150
R10374 VSS.n9235 VSS.n9234 150
R10375 VSS.n9239 VSS.n9238 150
R10376 VSS.n9364 VSS.n9282 150
R10377 VSS.n9362 VSS.n9361 150
R10378 VSS.n9358 VSS.n9357 150
R10379 VSS.n9354 VSS.n9353 150
R10380 VSS.n9346 VSS.n9345 150
R10381 VSS.n9342 VSS.n9341 150
R10382 VSS.n9338 VSS.n9337 150
R10383 VSS.n9334 VSS.n9290 150
R10384 VSS.n10172 VSS.n9281 150
R10385 VSS.n9321 VSS.n9320 150
R10386 VSS.n9325 VSS.n9324 150
R10387 VSS.n9329 VSS.n9328 150
R10388 VSS.n9454 VSS.n9372 150
R10389 VSS.n9452 VSS.n9451 150
R10390 VSS.n9448 VSS.n9447 150
R10391 VSS.n9444 VSS.n9443 150
R10392 VSS.n9436 VSS.n9435 150
R10393 VSS.n9432 VSS.n9431 150
R10394 VSS.n9428 VSS.n9427 150
R10395 VSS.n9424 VSS.n9380 150
R10396 VSS.n10082 VSS.n9371 150
R10397 VSS.n9411 VSS.n9410 150
R10398 VSS.n9415 VSS.n9414 150
R10399 VSS.n9419 VSS.n9418 150
R10400 VSS.n9544 VSS.n9462 150
R10401 VSS.n9542 VSS.n9541 150
R10402 VSS.n9538 VSS.n9537 150
R10403 VSS.n9534 VSS.n9533 150
R10404 VSS.n9526 VSS.n9525 150
R10405 VSS.n9522 VSS.n9521 150
R10406 VSS.n9518 VSS.n9517 150
R10407 VSS.n9514 VSS.n9470 150
R10408 VSS.n9992 VSS.n9461 150
R10409 VSS.n9501 VSS.n9500 150
R10410 VSS.n9505 VSS.n9504 150
R10411 VSS.n9509 VSS.n9508 150
R10412 VSS.n9634 VSS.n9552 150
R10413 VSS.n9632 VSS.n9631 150
R10414 VSS.n9628 VSS.n9627 150
R10415 VSS.n9624 VSS.n9623 150
R10416 VSS.n9616 VSS.n9615 150
R10417 VSS.n9612 VSS.n9611 150
R10418 VSS.n9608 VSS.n9607 150
R10419 VSS.n9604 VSS.n9560 150
R10420 VSS.n9902 VSS.n9551 150
R10421 VSS.n9591 VSS.n9590 150
R10422 VSS.n9595 VSS.n9594 150
R10423 VSS.n9599 VSS.n9598 150
R10424 VSS.n9724 VSS.n9642 150
R10425 VSS.n9722 VSS.n9721 150
R10426 VSS.n9718 VSS.n9717 150
R10427 VSS.n9714 VSS.n9713 150
R10428 VSS.n9706 VSS.n9705 150
R10429 VSS.n9702 VSS.n9701 150
R10430 VSS.n9698 VSS.n9697 150
R10431 VSS.n9694 VSS.n9650 150
R10432 VSS.n9812 VSS.n9641 150
R10433 VSS.n9681 VSS.n9680 150
R10434 VSS.n9685 VSS.n9684 150
R10435 VSS.n9689 VSS.n9688 150
R10436 VSS.n10312 VSS.n10311 150
R10437 VSS.n10308 VSS.n10307 150
R10438 VSS.n10304 VSS.n10303 150
R10439 VSS.n10300 VSS.n9165 150
R10440 VSS.n10295 VSS.n10294 150
R10441 VSS.n10291 VSS.n10290 150
R10442 VSS.n10287 VSS.n10286 150
R10443 VSS.n10283 VSS.n10282 150
R10444 VSS.n10267 VSS.n9164 150
R10445 VSS.n10271 VSS.n10270 150
R10446 VSS.n10275 VSS.n10274 150
R10447 VSS.n10279 VSS.n10278 150
R10448 VSS.n6694 VSS.n6693 150
R10449 VSS.n6698 VSS.n6697 150
R10450 VSS.n6702 VSS.n6701 150
R10451 VSS.n6706 VSS.n6705 150
R10452 VSS.n6714 VSS.n6713 150
R10453 VSS.n6718 VSS.n6717 150
R10454 VSS.n6723 VSS.n6658 150
R10455 VSS.n6725 VSS.n6638 150
R10456 VSS.n6673 VSS.n6672 150
R10457 VSS.n6669 VSS.n6668 150
R10458 VSS.n6665 VSS.n6664 150
R10459 VSS.n6661 VSS.n6660 150
R10460 VSS.n6677 VSS.n6676 150
R10461 VSS.n5731 VSS.n5670 150
R10462 VSS.n5727 VSS.n5683 150
R10463 VSS.n5725 VSS.n5724 150
R10464 VSS.n5721 VSS.n5720 150
R10465 VSS.n5713 VSS.n5712 150
R10466 VSS.n5709 VSS.n5708 150
R10467 VSS.n5705 VSS.n5704 150
R10468 VSS.n5701 VSS.n5678 150
R10469 VSS.n5734 VSS.n3631 150
R10470 VSS.n5688 VSS.n5687 150
R10471 VSS.n5692 VSS.n5691 150
R10472 VSS.n5696 VSS.n5695 150
R10473 VSS.n5853 VSS.n5792 150
R10474 VSS.n5849 VSS.n5805 150
R10475 VSS.n5847 VSS.n5846 150
R10476 VSS.n5843 VSS.n5842 150
R10477 VSS.n5835 VSS.n5834 150
R10478 VSS.n5831 VSS.n5830 150
R10479 VSS.n5827 VSS.n5826 150
R10480 VSS.n5823 VSS.n5800 150
R10481 VSS.n5856 VSS.n3573 150
R10482 VSS.n5810 VSS.n5809 150
R10483 VSS.n5814 VSS.n5813 150
R10484 VSS.n5818 VSS.n5817 150
R10485 VSS.n5975 VSS.n5914 150
R10486 VSS.n5971 VSS.n5927 150
R10487 VSS.n5969 VSS.n5968 150
R10488 VSS.n5965 VSS.n5964 150
R10489 VSS.n5957 VSS.n5956 150
R10490 VSS.n5953 VSS.n5952 150
R10491 VSS.n5949 VSS.n5948 150
R10492 VSS.n5945 VSS.n5922 150
R10493 VSS.n5978 VSS.n3515 150
R10494 VSS.n5932 VSS.n5931 150
R10495 VSS.n5936 VSS.n5935 150
R10496 VSS.n5940 VSS.n5939 150
R10497 VSS.n6097 VSS.n6036 150
R10498 VSS.n6093 VSS.n6049 150
R10499 VSS.n6091 VSS.n6090 150
R10500 VSS.n6087 VSS.n6086 150
R10501 VSS.n6079 VSS.n6078 150
R10502 VSS.n6075 VSS.n6074 150
R10503 VSS.n6071 VSS.n6070 150
R10504 VSS.n6067 VSS.n6044 150
R10505 VSS.n6100 VSS.n3457 150
R10506 VSS.n6054 VSS.n6053 150
R10507 VSS.n6058 VSS.n6057 150
R10508 VSS.n6062 VSS.n6061 150
R10509 VSS.n6219 VSS.n6158 150
R10510 VSS.n6215 VSS.n6171 150
R10511 VSS.n6213 VSS.n6212 150
R10512 VSS.n6209 VSS.n6208 150
R10513 VSS.n6201 VSS.n6200 150
R10514 VSS.n6197 VSS.n6196 150
R10515 VSS.n6193 VSS.n6192 150
R10516 VSS.n6189 VSS.n6166 150
R10517 VSS.n6222 VSS.n3399 150
R10518 VSS.n6176 VSS.n6175 150
R10519 VSS.n6180 VSS.n6179 150
R10520 VSS.n6184 VSS.n6183 150
R10521 VSS.n6341 VSS.n6280 150
R10522 VSS.n6337 VSS.n6293 150
R10523 VSS.n6335 VSS.n6334 150
R10524 VSS.n6331 VSS.n6330 150
R10525 VSS.n6323 VSS.n6322 150
R10526 VSS.n6319 VSS.n6318 150
R10527 VSS.n6315 VSS.n6314 150
R10528 VSS.n6311 VSS.n6288 150
R10529 VSS.n6344 VSS.n3341 150
R10530 VSS.n6298 VSS.n6297 150
R10531 VSS.n6302 VSS.n6301 150
R10532 VSS.n6306 VSS.n6305 150
R10533 VSS.n6463 VSS.n6402 150
R10534 VSS.n6459 VSS.n6415 150
R10535 VSS.n6457 VSS.n6456 150
R10536 VSS.n6453 VSS.n6452 150
R10537 VSS.n6445 VSS.n6444 150
R10538 VSS.n6441 VSS.n6440 150
R10539 VSS.n6437 VSS.n6436 150
R10540 VSS.n6433 VSS.n6410 150
R10541 VSS.n6466 VSS.n3283 150
R10542 VSS.n6420 VSS.n6419 150
R10543 VSS.n6424 VSS.n6423 150
R10544 VSS.n6428 VSS.n6427 150
R10545 VSS.n6542 VSS.n6540 150
R10546 VSS.n6546 VSS.n6533 150
R10547 VSS.n6550 VSS.n6548 150
R10548 VSS.n6554 VSS.n6531 150
R10549 VSS.n6562 VSS.n6529 150
R10550 VSS.n6566 VSS.n6564 150
R10551 VSS.n6570 VSS.n6527 150
R10552 VSS.n6573 VSS.n6572 150
R10553 VSS.n6587 VSS.n3158 150
R10554 VSS.n6585 VSS.n6584 150
R10555 VSS.n6581 VSS.n6580 150
R10556 VSS.n6578 VSS.n6523 150
R10557 VSS.n92 VSS.n9 150
R10558 VSS.n90 VSS.n89 150
R10559 VSS.n86 VSS.n85 150
R10560 VSS.n82 VSS.n81 150
R10561 VSS.n74 VSS.n73 150
R10562 VSS.n70 VSS.n69 150
R10563 VSS.n66 VSS.n65 150
R10564 VSS.n62 VSS.n17 150
R10565 VSS.n1254 VSS.n8 150
R10566 VSS.n49 VSS.n48 150
R10567 VSS.n53 VSS.n52 150
R10568 VSS.n57 VSS.n56 150
R10569 VSS.n182 VSS.n100 150
R10570 VSS.n180 VSS.n179 150
R10571 VSS.n176 VSS.n175 150
R10572 VSS.n172 VSS.n171 150
R10573 VSS.n164 VSS.n163 150
R10574 VSS.n160 VSS.n159 150
R10575 VSS.n156 VSS.n155 150
R10576 VSS.n152 VSS.n108 150
R10577 VSS.n1170 VSS.n99 150
R10578 VSS.n139 VSS.n138 150
R10579 VSS.n143 VSS.n142 150
R10580 VSS.n147 VSS.n146 150
R10581 VSS.n272 VSS.n190 150
R10582 VSS.n270 VSS.n269 150
R10583 VSS.n266 VSS.n265 150
R10584 VSS.n262 VSS.n261 150
R10585 VSS.n254 VSS.n253 150
R10586 VSS.n250 VSS.n249 150
R10587 VSS.n246 VSS.n245 150
R10588 VSS.n242 VSS.n198 150
R10589 VSS.n1080 VSS.n189 150
R10590 VSS.n229 VSS.n228 150
R10591 VSS.n233 VSS.n232 150
R10592 VSS.n237 VSS.n236 150
R10593 VSS.n362 VSS.n280 150
R10594 VSS.n360 VSS.n359 150
R10595 VSS.n356 VSS.n355 150
R10596 VSS.n352 VSS.n351 150
R10597 VSS.n344 VSS.n343 150
R10598 VSS.n340 VSS.n339 150
R10599 VSS.n336 VSS.n335 150
R10600 VSS.n332 VSS.n288 150
R10601 VSS.n990 VSS.n279 150
R10602 VSS.n319 VSS.n318 150
R10603 VSS.n323 VSS.n322 150
R10604 VSS.n327 VSS.n326 150
R10605 VSS.n452 VSS.n370 150
R10606 VSS.n450 VSS.n449 150
R10607 VSS.n446 VSS.n445 150
R10608 VSS.n442 VSS.n441 150
R10609 VSS.n434 VSS.n433 150
R10610 VSS.n430 VSS.n429 150
R10611 VSS.n426 VSS.n425 150
R10612 VSS.n422 VSS.n378 150
R10613 VSS.n900 VSS.n369 150
R10614 VSS.n409 VSS.n408 150
R10615 VSS.n413 VSS.n412 150
R10616 VSS.n417 VSS.n416 150
R10617 VSS.n542 VSS.n460 150
R10618 VSS.n540 VSS.n539 150
R10619 VSS.n536 VSS.n535 150
R10620 VSS.n532 VSS.n531 150
R10621 VSS.n524 VSS.n523 150
R10622 VSS.n520 VSS.n519 150
R10623 VSS.n516 VSS.n515 150
R10624 VSS.n512 VSS.n468 150
R10625 VSS.n810 VSS.n459 150
R10626 VSS.n499 VSS.n498 150
R10627 VSS.n503 VSS.n502 150
R10628 VSS.n507 VSS.n506 150
R10629 VSS.n632 VSS.n550 150
R10630 VSS.n630 VSS.n629 150
R10631 VSS.n626 VSS.n625 150
R10632 VSS.n622 VSS.n621 150
R10633 VSS.n614 VSS.n613 150
R10634 VSS.n610 VSS.n609 150
R10635 VSS.n606 VSS.n605 150
R10636 VSS.n602 VSS.n558 150
R10637 VSS.n720 VSS.n549 150
R10638 VSS.n589 VSS.n588 150
R10639 VSS.n593 VSS.n592 150
R10640 VSS.n597 VSS.n596 150
R10641 VSS.n15664 VSS.n15663 146.25
R10642 VSS.n15665 VSS.n15664 146.25
R10643 VSS.n15662 VSS.n15640 146.25
R10644 VSS.n15640 VSS.n15639 146.25
R10645 VSS.n15661 VSS.n15660 146.25
R10646 VSS.n15660 VSS.n15659 146.25
R10647 VSS.n15642 VSS.n15641 146.25
R10648 VSS.n15658 VSS.n15642 146.25
R10649 VSS.n15656 VSS.n15655 146.25
R10650 VSS.n15657 VSS.n15656 146.25
R10651 VSS.n15654 VSS.n15644 146.25
R10652 VSS.n15644 VSS.n15643 146.25
R10653 VSS.n15653 VSS.n15652 146.25
R10654 VSS.n15652 VSS.n15651 146.25
R10655 VSS.n15646 VSS.n15645 146.25
R10656 VSS.n15650 VSS.n15646 146.25
R10657 VSS.n15648 VSS.n15647 146.25
R10658 VSS.n15649 VSS.n15648 146.25
R10659 VSS.n14041 VSS.n14040 146.25
R10660 VSS.n14043 VSS.n14041 146.25
R10661 VSS.n15948 VSS.n15947 146.25
R10662 VSS.n15947 VSS.n15946 146.25
R10663 VSS.n15638 VSS.n15637 146.25
R10664 VSS.n15666 VSS.n15638 146.25
R10665 VSS.n15669 VSS.n15668 146.25
R10666 VSS.n15668 VSS.n15667 146.25
R10667 VSS.n15898 VSS.n15897 146.25
R10668 VSS.n15897 VSS.n15896 146.25
R10669 VSS.n15899 VSS.n14066 146.25
R10670 VSS.n14066 VSS.n14065 146.25
R10671 VSS.n15901 VSS.n15900 146.25
R10672 VSS.n15902 VSS.n15901 146.25
R10673 VSS.n14064 VSS.n14063 146.25
R10674 VSS.n15903 VSS.n14064 146.25
R10675 VSS.n15906 VSS.n15905 146.25
R10676 VSS.n15905 VSS.n15904 146.25
R10677 VSS.n15907 VSS.n14062 146.25
R10678 VSS.n14062 VSS.n14061 146.25
R10679 VSS.n15909 VSS.n15908 146.25
R10680 VSS.n15910 VSS.n15909 146.25
R10681 VSS.n14060 VSS.n14059 146.25
R10682 VSS.n15911 VSS.n14060 146.25
R10683 VSS.n15914 VSS.n15913 146.25
R10684 VSS.n15913 VSS.n15912 146.25
R10685 VSS.n15915 VSS.n14058 146.25
R10686 VSS.n14058 VSS.n14057 146.25
R10687 VSS.n15917 VSS.n15916 146.25
R10688 VSS.n15918 VSS.n15917 146.25
R10689 VSS.n14068 VSS.n14067 146.25
R10690 VSS.n15895 VSS.n14068 146.25
R10691 VSS.n15893 VSS.n15892 146.25
R10692 VSS.n15894 VSS.n15893 146.25
R10693 VSS.n15436 VSS.n15435 146.25
R10694 VSS.n15437 VSS.n15436 146.25
R10695 VSS.n15434 VSS.n14147 146.25
R10696 VSS.n14147 VSS.n14146 146.25
R10697 VSS.n15433 VSS.n15432 146.25
R10698 VSS.n15432 VSS.n15431 146.25
R10699 VSS.n14150 VSS.n14149 146.25
R10700 VSS.n15430 VSS.n14150 146.25
R10701 VSS.n15428 VSS.n15427 146.25
R10702 VSS.n15429 VSS.n15428 146.25
R10703 VSS.n15426 VSS.n14152 146.25
R10704 VSS.n14152 VSS.n14151 146.25
R10705 VSS.n15425 VSS.n15424 146.25
R10706 VSS.n15424 VSS.n15423 146.25
R10707 VSS.n14154 VSS.n14153 146.25
R10708 VSS.n15422 VSS.n14154 146.25
R10709 VSS.n15420 VSS.n15419 146.25
R10710 VSS.n15421 VSS.n15420 146.25
R10711 VSS.n15418 VSS.n14156 146.25
R10712 VSS.n14156 VSS.n14155 146.25
R10713 VSS.n15417 VSS.n15416 146.25
R10714 VSS.n15416 VSS.n15415 146.25
R10715 VSS.n14148 VSS.n14145 146.25
R10716 VSS.n15438 VSS.n14145 146.25
R10717 VSS.n15440 VSS.n14136 146.25
R10718 VSS.n15440 VSS.n15439 146.25
R10719 VSS.n15077 VSS.n15076 146.25
R10720 VSS.n15078 VSS.n15077 146.25
R10721 VSS.n15075 VSS.n15053 146.25
R10722 VSS.n15053 VSS.n15052 146.25
R10723 VSS.n15074 VSS.n15073 146.25
R10724 VSS.n15073 VSS.n15072 146.25
R10725 VSS.n15055 VSS.n15054 146.25
R10726 VSS.n15071 VSS.n15055 146.25
R10727 VSS.n15069 VSS.n15068 146.25
R10728 VSS.n15070 VSS.n15069 146.25
R10729 VSS.n15067 VSS.n15057 146.25
R10730 VSS.n15057 VSS.n15056 146.25
R10731 VSS.n15066 VSS.n15065 146.25
R10732 VSS.n15065 VSS.n15064 146.25
R10733 VSS.n15059 VSS.n15058 146.25
R10734 VSS.n15063 VSS.n15059 146.25
R10735 VSS.n15061 VSS.n15060 146.25
R10736 VSS.n15062 VSS.n15061 146.25
R10737 VSS.n14210 VSS.n14208 146.25
R10738 VSS.n14208 VSS.n14207 146.25
R10739 VSS.n15387 VSS.n15386 146.25
R10740 VSS.n15388 VSS.n15387 146.25
R10741 VSS.n15051 VSS.n15050 146.25
R10742 VSS.n15079 VSS.n15051 146.25
R10743 VSS.n15082 VSS.n15081 146.25
R10744 VSS.n15081 VSS.n15080 146.25
R10745 VSS.n15337 VSS.n15336 146.25
R10746 VSS.n15338 VSS.n15337 146.25
R10747 VSS.n14233 VSS.n14232 146.25
R10748 VSS.n15339 VSS.n14233 146.25
R10749 VSS.n15342 VSS.n15341 146.25
R10750 VSS.n15341 VSS.n15340 146.25
R10751 VSS.n15343 VSS.n14231 146.25
R10752 VSS.n14231 VSS.n14230 146.25
R10753 VSS.n15345 VSS.n15344 146.25
R10754 VSS.n15346 VSS.n15345 146.25
R10755 VSS.n14229 VSS.n14228 146.25
R10756 VSS.n15347 VSS.n14229 146.25
R10757 VSS.n15350 VSS.n15349 146.25
R10758 VSS.n15349 VSS.n15348 146.25
R10759 VSS.n15351 VSS.n14227 146.25
R10760 VSS.n14227 VSS.n14226 146.25
R10761 VSS.n15353 VSS.n15352 146.25
R10762 VSS.n15354 VSS.n15353 146.25
R10763 VSS.n14225 VSS.n14224 146.25
R10764 VSS.n15355 VSS.n14225 146.25
R10765 VSS.n15358 VSS.n15357 146.25
R10766 VSS.n15357 VSS.n15356 146.25
R10767 VSS.n15335 VSS.n14235 146.25
R10768 VSS.n14235 VSS.n14234 146.25
R10769 VSS.n15334 VSS.n15333 146.25
R10770 VSS.n15333 VSS.n15332 146.25
R10771 VSS.n14312 VSS.n14309 146.25
R10772 VSS.n14860 VSS.n14309 146.25
R10773 VSS.n14858 VSS.n14857 146.25
R10774 VSS.n14859 VSS.n14858 146.25
R10775 VSS.n14856 VSS.n14311 146.25
R10776 VSS.n14311 VSS.n14310 146.25
R10777 VSS.n14855 VSS.n14854 146.25
R10778 VSS.n14854 VSS.n14853 146.25
R10779 VSS.n14314 VSS.n14313 146.25
R10780 VSS.n14852 VSS.n14314 146.25
R10781 VSS.n14850 VSS.n14849 146.25
R10782 VSS.n14851 VSS.n14850 146.25
R10783 VSS.n14848 VSS.n14316 146.25
R10784 VSS.n14316 VSS.n14315 146.25
R10785 VSS.n14847 VSS.n14846 146.25
R10786 VSS.n14846 VSS.n14845 146.25
R10787 VSS.n14318 VSS.n14317 146.25
R10788 VSS.n14844 VSS.n14318 146.25
R10789 VSS.n14842 VSS.n14841 146.25
R10790 VSS.n14843 VSS.n14842 146.25
R10791 VSS.n14840 VSS.n14320 146.25
R10792 VSS.n14320 VSS.n14319 146.25
R10793 VSS.n14862 VSS.n14308 146.25
R10794 VSS.n14862 VSS.n14861 146.25
R10795 VSS.n14864 VSS.n14863 146.25
R10796 VSS.n14863 VSS.n14301 146.25
R10797 VSS.n14468 VSS.n14467 146.25
R10798 VSS.n14469 VSS.n14468 146.25
R10799 VSS.n14466 VSS.n14444 146.25
R10800 VSS.n14444 VSS.n14443 146.25
R10801 VSS.n14465 VSS.n14464 146.25
R10802 VSS.n14464 VSS.n14463 146.25
R10803 VSS.n14446 VSS.n14445 146.25
R10804 VSS.n14462 VSS.n14446 146.25
R10805 VSS.n14460 VSS.n14459 146.25
R10806 VSS.n14461 VSS.n14460 146.25
R10807 VSS.n14458 VSS.n14448 146.25
R10808 VSS.n14448 VSS.n14447 146.25
R10809 VSS.n14457 VSS.n14456 146.25
R10810 VSS.n14456 VSS.n14455 146.25
R10811 VSS.n14450 VSS.n14449 146.25
R10812 VSS.n14454 VSS.n14450 146.25
R10813 VSS.n14452 VSS.n14451 146.25
R10814 VSS.n14453 VSS.n14452 146.25
R10815 VSS.n14337 VSS.n14336 146.25
R10816 VSS.n14339 VSS.n14337 146.25
R10817 VSS.n14778 VSS.n14777 146.25
R10818 VSS.n14777 VSS.n14776 146.25
R10819 VSS.n14442 VSS.n14441 146.25
R10820 VSS.n14470 VSS.n14442 146.25
R10821 VSS.n14473 VSS.n14472 146.25
R10822 VSS.n14472 VSS.n14471 146.25
R10823 VSS.n12107 VSS.n12106 146.25
R10824 VSS.n12108 VSS.n12107 146.25
R10825 VSS.n12099 VSS.n12098 146.25
R10826 VSS.n12109 VSS.n12099 146.25
R10827 VSS.n12112 VSS.n12111 146.25
R10828 VSS.n12111 VSS.n12110 146.25
R10829 VSS.n12113 VSS.n12097 146.25
R10830 VSS.n12097 VSS.n12096 146.25
R10831 VSS.n12115 VSS.n12114 146.25
R10832 VSS.n12116 VSS.n12115 146.25
R10833 VSS.n12095 VSS.n12094 146.25
R10834 VSS.n12117 VSS.n12095 146.25
R10835 VSS.n12120 VSS.n12119 146.25
R10836 VSS.n12119 VSS.n12118 146.25
R10837 VSS.n12121 VSS.n12093 146.25
R10838 VSS.n12093 VSS.n12092 146.25
R10839 VSS.n12123 VSS.n12122 146.25
R10840 VSS.n12124 VSS.n12123 146.25
R10841 VSS.n12090 VSS.n12089 146.25
R10842 VSS.n12125 VSS.n12090 146.25
R10843 VSS.n12163 VSS.n12162 146.25
R10844 VSS.n12162 VSS.n12161 146.25
R10845 VSS.n12105 VSS.n12101 146.25
R10846 VSS.n12101 VSS.n12100 146.25
R10847 VSS.n12104 VSS.n12103 146.25
R10848 VSS.n12103 VSS.n12102 146.25
R10849 VSS.n12412 VSS.n12411 146.25
R10850 VSS.n12413 VSS.n12412 146.25
R10851 VSS.n11538 VSS.n11537 146.25
R10852 VSS.n12414 VSS.n11538 146.25
R10853 VSS.n12417 VSS.n12416 146.25
R10854 VSS.n12416 VSS.n12415 146.25
R10855 VSS.n12418 VSS.n11536 146.25
R10856 VSS.n11536 VSS.n11535 146.25
R10857 VSS.n12420 VSS.n12419 146.25
R10858 VSS.n12421 VSS.n12420 146.25
R10859 VSS.n11534 VSS.n11533 146.25
R10860 VSS.n12422 VSS.n11534 146.25
R10861 VSS.n12425 VSS.n12424 146.25
R10862 VSS.n12424 VSS.n12423 146.25
R10863 VSS.n12426 VSS.n11532 146.25
R10864 VSS.n11532 VSS.n11531 146.25
R10865 VSS.n12428 VSS.n12427 146.25
R10866 VSS.n12429 VSS.n12428 146.25
R10867 VSS.n11530 VSS.n11529 146.25
R10868 VSS.n12430 VSS.n11530 146.25
R10869 VSS.n12433 VSS.n12432 146.25
R10870 VSS.n12432 VSS.n12431 146.25
R10871 VSS.n12410 VSS.n11540 146.25
R10872 VSS.n11540 VSS.n11539 146.25
R10873 VSS.n12409 VSS.n12408 146.25
R10874 VSS.n12408 VSS.n12407 146.25
R10875 VSS.n11802 VSS.n11801 146.25
R10876 VSS.n11801 VSS.n11800 146.25
R10877 VSS.n11777 VSS.n11776 146.25
R10878 VSS.n11799 VSS.n11777 146.25
R10879 VSS.n11797 VSS.n11796 146.25
R10880 VSS.n11798 VSS.n11797 146.25
R10881 VSS.n11795 VSS.n11779 146.25
R10882 VSS.n11779 VSS.n11778 146.25
R10883 VSS.n11794 VSS.n11793 146.25
R10884 VSS.n11793 VSS.n11792 146.25
R10885 VSS.n11781 VSS.n11780 146.25
R10886 VSS.n11791 VSS.n11781 146.25
R10887 VSS.n11789 VSS.n11788 146.25
R10888 VSS.n11790 VSS.n11789 146.25
R10889 VSS.n11787 VSS.n11783 146.25
R10890 VSS.n11783 VSS.n11782 146.25
R10891 VSS.n11786 VSS.n11785 146.25
R10892 VSS.n11785 VSS.n11784 146.25
R10893 VSS.n11514 VSS.n11512 146.25
R10894 VSS.n11512 VSS.n11511 146.25
R10895 VSS.n12461 VSS.n12460 146.25
R10896 VSS.n12462 VSS.n12461 146.25
R10897 VSS.n11803 VSS.n11609 146.25
R10898 VSS.n11609 VSS.n11607 146.25
R10899 VSS.n11805 VSS.n11804 146.25
R10900 VSS.n11806 VSS.n11805 146.25
R10901 VSS.n13392 VSS.n13391 146.25
R10902 VSS.n13393 VSS.n13392 146.25
R10903 VSS.n13390 VSS.n11487 146.25
R10904 VSS.n11487 VSS.n11486 146.25
R10905 VSS.n13389 VSS.n13388 146.25
R10906 VSS.n13388 VSS.n13387 146.25
R10907 VSS.n11489 VSS.n11488 146.25
R10908 VSS.n13386 VSS.n11489 146.25
R10909 VSS.n13384 VSS.n13383 146.25
R10910 VSS.n13385 VSS.n13384 146.25
R10911 VSS.n13382 VSS.n11491 146.25
R10912 VSS.n11491 VSS.n11490 146.25
R10913 VSS.n13381 VSS.n13380 146.25
R10914 VSS.n13380 VSS.n13379 146.25
R10915 VSS.n11493 VSS.n11492 146.25
R10916 VSS.n13378 VSS.n11493 146.25
R10917 VSS.n13376 VSS.n13375 146.25
R10918 VSS.n13377 VSS.n13376 146.25
R10919 VSS.n13374 VSS.n11495 146.25
R10920 VSS.n11495 VSS.n11494 146.25
R10921 VSS.n13373 VSS.n13372 146.25
R10922 VSS.n13372 VSS.n13371 146.25
R10923 VSS.n11484 VSS.n11482 146.25
R10924 VSS.n13394 VSS.n11484 146.25
R10925 VSS.n13397 VSS.n13396 146.25
R10926 VSS.n13396 VSS.n13395 146.25
R10927 VSS.n12514 VSS.n12513 146.25
R10928 VSS.n13319 VSS.n12514 146.25
R10929 VSS.n13322 VSS.n13321 146.25
R10930 VSS.n13321 VSS.n13320 146.25
R10931 VSS.n13323 VSS.n12512 146.25
R10932 VSS.n12512 VSS.n12511 146.25
R10933 VSS.n13325 VSS.n13324 146.25
R10934 VSS.n13326 VSS.n13325 146.25
R10935 VSS.n12510 VSS.n12509 146.25
R10936 VSS.n13327 VSS.n12510 146.25
R10937 VSS.n13330 VSS.n13329 146.25
R10938 VSS.n13329 VSS.n13328 146.25
R10939 VSS.n13331 VSS.n12508 146.25
R10940 VSS.n12508 VSS.n12507 146.25
R10941 VSS.n13334 VSS.n13333 146.25
R10942 VSS.n13335 VSS.n13334 146.25
R10943 VSS.n13332 VSS.n12506 146.25
R10944 VSS.n13336 VSS.n12506 146.25
R10945 VSS.n13338 VSS.n12505 146.25
R10946 VSS.n13338 VSS.n13337 146.25
R10947 VSS.n13340 VSS.n13339 146.25
R10948 VSS.n13339 VSS.n12500 146.25
R10949 VSS.n13317 VSS.n13316 146.25
R10950 VSS.n13318 VSS.n13317 146.25
R10951 VSS.n13315 VSS.n12516 146.25
R10952 VSS.n12516 VSS.n12515 146.25
R10953 VSS.n13143 VSS.n13142 146.25
R10954 VSS.n13144 VSS.n13143 146.25
R10955 VSS.n13141 VSS.n12588 146.25
R10956 VSS.n12588 VSS.n12587 146.25
R10957 VSS.n13140 VSS.n13139 146.25
R10958 VSS.n13139 VSS.n13138 146.25
R10959 VSS.n12590 VSS.n12589 146.25
R10960 VSS.n13137 VSS.n12590 146.25
R10961 VSS.n13135 VSS.n13134 146.25
R10962 VSS.n13136 VSS.n13135 146.25
R10963 VSS.n13133 VSS.n12592 146.25
R10964 VSS.n12592 VSS.n12591 146.25
R10965 VSS.n13132 VSS.n13131 146.25
R10966 VSS.n13131 VSS.n13130 146.25
R10967 VSS.n12594 VSS.n12593 146.25
R10968 VSS.n13129 VSS.n12594 146.25
R10969 VSS.n13127 VSS.n13126 146.25
R10970 VSS.n13128 VSS.n13127 146.25
R10971 VSS.n13125 VSS.n12596 146.25
R10972 VSS.n12596 VSS.n12595 146.25
R10973 VSS.n13124 VSS.n13123 146.25
R10974 VSS.n13123 VSS.n13122 146.25
R10975 VSS.n12586 VSS.n12585 146.25
R10976 VSS.n13145 VSS.n12586 146.25
R10977 VSS.n13148 VSS.n13147 146.25
R10978 VSS.n13147 VSS.n13146 146.25
R10979 VSS.n12655 VSS.n12654 146.25
R10980 VSS.n13070 VSS.n12655 146.25
R10981 VSS.n13073 VSS.n13072 146.25
R10982 VSS.n13072 VSS.n13071 146.25
R10983 VSS.n13074 VSS.n12653 146.25
R10984 VSS.n12653 VSS.n12652 146.25
R10985 VSS.n13076 VSS.n13075 146.25
R10986 VSS.n13077 VSS.n13076 146.25
R10987 VSS.n12651 VSS.n12650 146.25
R10988 VSS.n13078 VSS.n12651 146.25
R10989 VSS.n13081 VSS.n13080 146.25
R10990 VSS.n13080 VSS.n13079 146.25
R10991 VSS.n13082 VSS.n12649 146.25
R10992 VSS.n12649 VSS.n12648 146.25
R10993 VSS.n13085 VSS.n13084 146.25
R10994 VSS.n13086 VSS.n13085 146.25
R10995 VSS.n13083 VSS.n12647 146.25
R10996 VSS.n13087 VSS.n12647 146.25
R10997 VSS.n13089 VSS.n12646 146.25
R10998 VSS.n13089 VSS.n13088 146.25
R10999 VSS.n13091 VSS.n13090 146.25
R11000 VSS.n13090 VSS.n12641 146.25
R11001 VSS.n13068 VSS.n13067 146.25
R11002 VSS.n13069 VSS.n13068 146.25
R11003 VSS.n13066 VSS.n12657 146.25
R11004 VSS.n12657 VSS.n12656 146.25
R11005 VSS.n8851 VSS.n8850 146.25
R11006 VSS.n8850 VSS.n8849 146.25
R11007 VSS.n6970 VSS.n6969 146.25
R11008 VSS.n8848 VSS.n6970 146.25
R11009 VSS.n8846 VSS.n8845 146.25
R11010 VSS.n8847 VSS.n8846 146.25
R11011 VSS.n8844 VSS.n6972 146.25
R11012 VSS.n6972 VSS.n6971 146.25
R11013 VSS.n8843 VSS.n8842 146.25
R11014 VSS.n8842 VSS.n8841 146.25
R11015 VSS.n6974 VSS.n6973 146.25
R11016 VSS.n8840 VSS.n6974 146.25
R11017 VSS.n8838 VSS.n8837 146.25
R11018 VSS.n8839 VSS.n8838 146.25
R11019 VSS.n8836 VSS.n6976 146.25
R11020 VSS.n6976 VSS.n6975 146.25
R11021 VSS.n8835 VSS.n8834 146.25
R11022 VSS.n8834 VSS.n8833 146.25
R11023 VSS.n6978 VSS.n6977 146.25
R11024 VSS.n8832 VSS.n6978 146.25
R11025 VSS.n8830 VSS.n8829 146.25
R11026 VSS.n8831 VSS.n8830 146.25
R11027 VSS.n8852 VSS.n6967 146.25
R11028 VSS.n6967 VSS.n6966 146.25
R11029 VSS.n8854 VSS.n8853 146.25
R11030 VSS.n8855 VSS.n8854 146.25
R11031 VSS.n8777 VSS.n7253 146.25
R11032 VSS.n7253 VSS.n7252 146.25
R11033 VSS.n8779 VSS.n8778 146.25
R11034 VSS.n8780 VSS.n8779 146.25
R11035 VSS.n7251 VSS.n7250 146.25
R11036 VSS.n8781 VSS.n7251 146.25
R11037 VSS.n8784 VSS.n8783 146.25
R11038 VSS.n8783 VSS.n8782 146.25
R11039 VSS.n8785 VSS.n7249 146.25
R11040 VSS.n7249 VSS.n7248 146.25
R11041 VSS.n8787 VSS.n8786 146.25
R11042 VSS.n8788 VSS.n8787 146.25
R11043 VSS.n7247 VSS.n7246 146.25
R11044 VSS.n8789 VSS.n7247 146.25
R11045 VSS.n8793 VSS.n8792 146.25
R11046 VSS.n8792 VSS.n8791 146.25
R11047 VSS.n8794 VSS.n7245 146.25
R11048 VSS.n8790 VSS.n7245 146.25
R11049 VSS.n8796 VSS.n8795 146.25
R11050 VSS.n8796 VSS.n7244 146.25
R11051 VSS.n8797 VSS.n7239 146.25
R11052 VSS.n8798 VSS.n8797 146.25
R11053 VSS.n8776 VSS.n8775 146.25
R11054 VSS.n8775 VSS.n8774 146.25
R11055 VSS.n7255 VSS.n7254 146.25
R11056 VSS.n8773 VSS.n7255 146.25
R11057 VSS.n8629 VSS.n8628 146.25
R11058 VSS.n8628 VSS.n8627 146.25
R11059 VSS.n7326 VSS.n7325 146.25
R11060 VSS.n8626 VSS.n7326 146.25
R11061 VSS.n8624 VSS.n8623 146.25
R11062 VSS.n8625 VSS.n8624 146.25
R11063 VSS.n8622 VSS.n7328 146.25
R11064 VSS.n7328 VSS.n7327 146.25
R11065 VSS.n8621 VSS.n8620 146.25
R11066 VSS.n8620 VSS.n8619 146.25
R11067 VSS.n7330 VSS.n7329 146.25
R11068 VSS.n8618 VSS.n7330 146.25
R11069 VSS.n8616 VSS.n8615 146.25
R11070 VSS.n8617 VSS.n8616 146.25
R11071 VSS.n8614 VSS.n7332 146.25
R11072 VSS.n7332 VSS.n7331 146.25
R11073 VSS.n8613 VSS.n8612 146.25
R11074 VSS.n8612 VSS.n8611 146.25
R11075 VSS.n7334 VSS.n7333 146.25
R11076 VSS.n8610 VSS.n7334 146.25
R11077 VSS.n8608 VSS.n8607 146.25
R11078 VSS.n8609 VSS.n8608 146.25
R11079 VSS.n8630 VSS.n7323 146.25
R11080 VSS.n7323 VSS.n7321 146.25
R11081 VSS.n8632 VSS.n8631 146.25
R11082 VSS.n8633 VSS.n8632 146.25
R11083 VSS.n8555 VSS.n7393 146.25
R11084 VSS.n7393 VSS.n7392 146.25
R11085 VSS.n8557 VSS.n8556 146.25
R11086 VSS.n8558 VSS.n8557 146.25
R11087 VSS.n7391 VSS.n7390 146.25
R11088 VSS.n8559 VSS.n7391 146.25
R11089 VSS.n8562 VSS.n8561 146.25
R11090 VSS.n8561 VSS.n8560 146.25
R11091 VSS.n8563 VSS.n7389 146.25
R11092 VSS.n7389 VSS.n7388 146.25
R11093 VSS.n8565 VSS.n8564 146.25
R11094 VSS.n8566 VSS.n8565 146.25
R11095 VSS.n7387 VSS.n7386 146.25
R11096 VSS.n8567 VSS.n7387 146.25
R11097 VSS.n8571 VSS.n8570 146.25
R11098 VSS.n8570 VSS.n8569 146.25
R11099 VSS.n8572 VSS.n7385 146.25
R11100 VSS.n8568 VSS.n7385 146.25
R11101 VSS.n8574 VSS.n8573 146.25
R11102 VSS.n8574 VSS.n7384 146.25
R11103 VSS.n8575 VSS.n7379 146.25
R11104 VSS.n8576 VSS.n8575 146.25
R11105 VSS.n8554 VSS.n8553 146.25
R11106 VSS.n8553 VSS.n8552 146.25
R11107 VSS.n7395 VSS.n7394 146.25
R11108 VSS.n8551 VSS.n7395 146.25
R11109 VSS.n8271 VSS.n8270 146.25
R11110 VSS.n8270 VSS.n8269 146.25
R11111 VSS.n7466 VSS.n7465 146.25
R11112 VSS.n8268 VSS.n7466 146.25
R11113 VSS.n8266 VSS.n8265 146.25
R11114 VSS.n8267 VSS.n8266 146.25
R11115 VSS.n8264 VSS.n7468 146.25
R11116 VSS.n7468 VSS.n7467 146.25
R11117 VSS.n8263 VSS.n8262 146.25
R11118 VSS.n8262 VSS.n8261 146.25
R11119 VSS.n7470 VSS.n7469 146.25
R11120 VSS.n8260 VSS.n7470 146.25
R11121 VSS.n8258 VSS.n8257 146.25
R11122 VSS.n8259 VSS.n8258 146.25
R11123 VSS.n8256 VSS.n7472 146.25
R11124 VSS.n7472 VSS.n7471 146.25
R11125 VSS.n8255 VSS.n8254 146.25
R11126 VSS.n8254 VSS.n8253 146.25
R11127 VSS.n7474 VSS.n7473 146.25
R11128 VSS.n8252 VSS.n7474 146.25
R11129 VSS.n8250 VSS.n8249 146.25
R11130 VSS.n8251 VSS.n8250 146.25
R11131 VSS.n8272 VSS.n7463 146.25
R11132 VSS.n7463 VSS.n7461 146.25
R11133 VSS.n8274 VSS.n8273 146.25
R11134 VSS.n8275 VSS.n8274 146.25
R11135 VSS.n8197 VSS.n7533 146.25
R11136 VSS.n7533 VSS.n7532 146.25
R11137 VSS.n8199 VSS.n8198 146.25
R11138 VSS.n8200 VSS.n8199 146.25
R11139 VSS.n7531 VSS.n7530 146.25
R11140 VSS.n8201 VSS.n7531 146.25
R11141 VSS.n8204 VSS.n8203 146.25
R11142 VSS.n8203 VSS.n8202 146.25
R11143 VSS.n8205 VSS.n7529 146.25
R11144 VSS.n7529 VSS.n7528 146.25
R11145 VSS.n8207 VSS.n8206 146.25
R11146 VSS.n8208 VSS.n8207 146.25
R11147 VSS.n7527 VSS.n7526 146.25
R11148 VSS.n8209 VSS.n7527 146.25
R11149 VSS.n8213 VSS.n8212 146.25
R11150 VSS.n8212 VSS.n8211 146.25
R11151 VSS.n8214 VSS.n7525 146.25
R11152 VSS.n8210 VSS.n7525 146.25
R11153 VSS.n8216 VSS.n8215 146.25
R11154 VSS.n8216 VSS.n7524 146.25
R11155 VSS.n8217 VSS.n7519 146.25
R11156 VSS.n8218 VSS.n8217 146.25
R11157 VSS.n8196 VSS.n8195 146.25
R11158 VSS.n8195 VSS.n8194 146.25
R11159 VSS.n7535 VSS.n7534 146.25
R11160 VSS.n8193 VSS.n7535 146.25
R11161 VSS.n7913 VSS.n7912 146.25
R11162 VSS.n7912 VSS.n7911 146.25
R11163 VSS.n7606 VSS.n7605 146.25
R11164 VSS.n7910 VSS.n7606 146.25
R11165 VSS.n7908 VSS.n7907 146.25
R11166 VSS.n7909 VSS.n7908 146.25
R11167 VSS.n7906 VSS.n7608 146.25
R11168 VSS.n7608 VSS.n7607 146.25
R11169 VSS.n7905 VSS.n7904 146.25
R11170 VSS.n7904 VSS.n7903 146.25
R11171 VSS.n7610 VSS.n7609 146.25
R11172 VSS.n7902 VSS.n7610 146.25
R11173 VSS.n7900 VSS.n7899 146.25
R11174 VSS.n7901 VSS.n7900 146.25
R11175 VSS.n7898 VSS.n7612 146.25
R11176 VSS.n7612 VSS.n7611 146.25
R11177 VSS.n7897 VSS.n7896 146.25
R11178 VSS.n7896 VSS.n7895 146.25
R11179 VSS.n7614 VSS.n7613 146.25
R11180 VSS.n7894 VSS.n7614 146.25
R11181 VSS.n7892 VSS.n7891 146.25
R11182 VSS.n7893 VSS.n7892 146.25
R11183 VSS.n7914 VSS.n7603 146.25
R11184 VSS.n7603 VSS.n7601 146.25
R11185 VSS.n7916 VSS.n7915 146.25
R11186 VSS.n7917 VSS.n7916 146.25
R11187 VSS.n3685 VSS.n3684 146.25
R11188 VSS.n5583 VSS.n3685 146.25
R11189 VSS.n5586 VSS.n5585 146.25
R11190 VSS.n5585 VSS.n5584 146.25
R11191 VSS.n5587 VSS.n3683 146.25
R11192 VSS.n3683 VSS.n3682 146.25
R11193 VSS.n5589 VSS.n5588 146.25
R11194 VSS.n5590 VSS.n5589 146.25
R11195 VSS.n3681 VSS.n3680 146.25
R11196 VSS.n5591 VSS.n3681 146.25
R11197 VSS.n5594 VSS.n5593 146.25
R11198 VSS.n5593 VSS.n5592 146.25
R11199 VSS.n5595 VSS.n3679 146.25
R11200 VSS.n3679 VSS.n3678 146.25
R11201 VSS.n5598 VSS.n5597 146.25
R11202 VSS.n5599 VSS.n5598 146.25
R11203 VSS.n5596 VSS.n3677 146.25
R11204 VSS.n5600 VSS.n3677 146.25
R11205 VSS.n5602 VSS.n3676 146.25
R11206 VSS.n5602 VSS.n5601 146.25
R11207 VSS.n5604 VSS.n5603 146.25
R11208 VSS.n5603 VSS.n3671 146.25
R11209 VSS.n5581 VSS.n5580 146.25
R11210 VSS.n5582 VSS.n5581 146.25
R11211 VSS.n5579 VSS.n3687 146.25
R11212 VSS.n3687 VSS.n3686 146.25
R11213 VSS.n5310 VSS.n5309 146.25
R11214 VSS.n5311 VSS.n5310 146.25
R11215 VSS.n5308 VSS.n3759 146.25
R11216 VSS.n3759 VSS.n3758 146.25
R11217 VSS.n5307 VSS.n5306 146.25
R11218 VSS.n5306 VSS.n5305 146.25
R11219 VSS.n3761 VSS.n3760 146.25
R11220 VSS.n5304 VSS.n3761 146.25
R11221 VSS.n5302 VSS.n5301 146.25
R11222 VSS.n5303 VSS.n5302 146.25
R11223 VSS.n5300 VSS.n3763 146.25
R11224 VSS.n3763 VSS.n3762 146.25
R11225 VSS.n5299 VSS.n5298 146.25
R11226 VSS.n5298 VSS.n5297 146.25
R11227 VSS.n3765 VSS.n3764 146.25
R11228 VSS.n5296 VSS.n3765 146.25
R11229 VSS.n5294 VSS.n5293 146.25
R11230 VSS.n5295 VSS.n5294 146.25
R11231 VSS.n5292 VSS.n3767 146.25
R11232 VSS.n3767 VSS.n3766 146.25
R11233 VSS.n5291 VSS.n5290 146.25
R11234 VSS.n5290 VSS.n5289 146.25
R11235 VSS.n3757 VSS.n3756 146.25
R11236 VSS.n5312 VSS.n3757 146.25
R11237 VSS.n5315 VSS.n5314 146.25
R11238 VSS.n5314 VSS.n5313 146.25
R11239 VSS.n3826 VSS.n3825 146.25
R11240 VSS.n5237 VSS.n3826 146.25
R11241 VSS.n5240 VSS.n5239 146.25
R11242 VSS.n5239 VSS.n5238 146.25
R11243 VSS.n5241 VSS.n3824 146.25
R11244 VSS.n3824 VSS.n3823 146.25
R11245 VSS.n5243 VSS.n5242 146.25
R11246 VSS.n5244 VSS.n5243 146.25
R11247 VSS.n3822 VSS.n3821 146.25
R11248 VSS.n5245 VSS.n3822 146.25
R11249 VSS.n5248 VSS.n5247 146.25
R11250 VSS.n5247 VSS.n5246 146.25
R11251 VSS.n5249 VSS.n3820 146.25
R11252 VSS.n3820 VSS.n3819 146.25
R11253 VSS.n5252 VSS.n5251 146.25
R11254 VSS.n5253 VSS.n5252 146.25
R11255 VSS.n5250 VSS.n3818 146.25
R11256 VSS.n5254 VSS.n3818 146.25
R11257 VSS.n5256 VSS.n3817 146.25
R11258 VSS.n5256 VSS.n5255 146.25
R11259 VSS.n5258 VSS.n5257 146.25
R11260 VSS.n5257 VSS.n3812 146.25
R11261 VSS.n5235 VSS.n5234 146.25
R11262 VSS.n5236 VSS.n5235 146.25
R11263 VSS.n5233 VSS.n3828 146.25
R11264 VSS.n3828 VSS.n3827 146.25
R11265 VSS.n4953 VSS.n4952 146.25
R11266 VSS.n4954 VSS.n4953 146.25
R11267 VSS.n4951 VSS.n3900 146.25
R11268 VSS.n3900 VSS.n3899 146.25
R11269 VSS.n4950 VSS.n4949 146.25
R11270 VSS.n4949 VSS.n4948 146.25
R11271 VSS.n3902 VSS.n3901 146.25
R11272 VSS.n4947 VSS.n3902 146.25
R11273 VSS.n4945 VSS.n4944 146.25
R11274 VSS.n4946 VSS.n4945 146.25
R11275 VSS.n4943 VSS.n3904 146.25
R11276 VSS.n3904 VSS.n3903 146.25
R11277 VSS.n4942 VSS.n4941 146.25
R11278 VSS.n4941 VSS.n4940 146.25
R11279 VSS.n3906 VSS.n3905 146.25
R11280 VSS.n4939 VSS.n3906 146.25
R11281 VSS.n4937 VSS.n4936 146.25
R11282 VSS.n4938 VSS.n4937 146.25
R11283 VSS.n4935 VSS.n3908 146.25
R11284 VSS.n3908 VSS.n3907 146.25
R11285 VSS.n4934 VSS.n4933 146.25
R11286 VSS.n4933 VSS.n4932 146.25
R11287 VSS.n3898 VSS.n3897 146.25
R11288 VSS.n4955 VSS.n3898 146.25
R11289 VSS.n4958 VSS.n4957 146.25
R11290 VSS.n4957 VSS.n4956 146.25
R11291 VSS.n3967 VSS.n3966 146.25
R11292 VSS.n4880 VSS.n3967 146.25
R11293 VSS.n4883 VSS.n4882 146.25
R11294 VSS.n4882 VSS.n4881 146.25
R11295 VSS.n4884 VSS.n3965 146.25
R11296 VSS.n3965 VSS.n3964 146.25
R11297 VSS.n4886 VSS.n4885 146.25
R11298 VSS.n4887 VSS.n4886 146.25
R11299 VSS.n3963 VSS.n3962 146.25
R11300 VSS.n4888 VSS.n3963 146.25
R11301 VSS.n4891 VSS.n4890 146.25
R11302 VSS.n4890 VSS.n4889 146.25
R11303 VSS.n4892 VSS.n3961 146.25
R11304 VSS.n3961 VSS.n3960 146.25
R11305 VSS.n4895 VSS.n4894 146.25
R11306 VSS.n4896 VSS.n4895 146.25
R11307 VSS.n4893 VSS.n3959 146.25
R11308 VSS.n4897 VSS.n3959 146.25
R11309 VSS.n4899 VSS.n3958 146.25
R11310 VSS.n4899 VSS.n4898 146.25
R11311 VSS.n4901 VSS.n4900 146.25
R11312 VSS.n4900 VSS.n3953 146.25
R11313 VSS.n4878 VSS.n4877 146.25
R11314 VSS.n4879 VSS.n4878 146.25
R11315 VSS.n4876 VSS.n3969 146.25
R11316 VSS.n3969 VSS.n3968 146.25
R11317 VSS.n4596 VSS.n4595 146.25
R11318 VSS.n4597 VSS.n4596 146.25
R11319 VSS.n4594 VSS.n4041 146.25
R11320 VSS.n4041 VSS.n4040 146.25
R11321 VSS.n4593 VSS.n4592 146.25
R11322 VSS.n4592 VSS.n4591 146.25
R11323 VSS.n4043 VSS.n4042 146.25
R11324 VSS.n4590 VSS.n4043 146.25
R11325 VSS.n4588 VSS.n4587 146.25
R11326 VSS.n4589 VSS.n4588 146.25
R11327 VSS.n4586 VSS.n4045 146.25
R11328 VSS.n4045 VSS.n4044 146.25
R11329 VSS.n4585 VSS.n4584 146.25
R11330 VSS.n4584 VSS.n4583 146.25
R11331 VSS.n4047 VSS.n4046 146.25
R11332 VSS.n4582 VSS.n4047 146.25
R11333 VSS.n4580 VSS.n4579 146.25
R11334 VSS.n4581 VSS.n4580 146.25
R11335 VSS.n4578 VSS.n4049 146.25
R11336 VSS.n4049 VSS.n4048 146.25
R11337 VSS.n4577 VSS.n4576 146.25
R11338 VSS.n4576 VSS.n4575 146.25
R11339 VSS.n4039 VSS.n4038 146.25
R11340 VSS.n4598 VSS.n4039 146.25
R11341 VSS.n4601 VSS.n4600 146.25
R11342 VSS.n4600 VSS.n4599 146.25
R11343 VSS.n4108 VSS.n4107 146.25
R11344 VSS.n4523 VSS.n4108 146.25
R11345 VSS.n4526 VSS.n4525 146.25
R11346 VSS.n4525 VSS.n4524 146.25
R11347 VSS.n4527 VSS.n4106 146.25
R11348 VSS.n4106 VSS.n4105 146.25
R11349 VSS.n4529 VSS.n4528 146.25
R11350 VSS.n4530 VSS.n4529 146.25
R11351 VSS.n4104 VSS.n4103 146.25
R11352 VSS.n4531 VSS.n4104 146.25
R11353 VSS.n4534 VSS.n4533 146.25
R11354 VSS.n4533 VSS.n4532 146.25
R11355 VSS.n4535 VSS.n4102 146.25
R11356 VSS.n4102 VSS.n4101 146.25
R11357 VSS.n4538 VSS.n4537 146.25
R11358 VSS.n4539 VSS.n4538 146.25
R11359 VSS.n4536 VSS.n4100 146.25
R11360 VSS.n4540 VSS.n4100 146.25
R11361 VSS.n4542 VSS.n4099 146.25
R11362 VSS.n4542 VSS.n4541 146.25
R11363 VSS.n4544 VSS.n4543 146.25
R11364 VSS.n4543 VSS.n4094 146.25
R11365 VSS.n4521 VSS.n4520 146.25
R11366 VSS.n4522 VSS.n4521 146.25
R11367 VSS.n4519 VSS.n4110 146.25
R11368 VSS.n4110 VSS.n4109 146.25
R11369 VSS.n2972 VSS.n2971 146.25
R11370 VSS.n2971 VSS.n2970 146.25
R11371 VSS.n2973 VSS.n1307 146.25
R11372 VSS.n1307 VSS.n1306 146.25
R11373 VSS.n2975 VSS.n2974 146.25
R11374 VSS.n2976 VSS.n2975 146.25
R11375 VSS.n1305 VSS.n1304 146.25
R11376 VSS.n2977 VSS.n1305 146.25
R11377 VSS.n2980 VSS.n2979 146.25
R11378 VSS.n2979 VSS.n2978 146.25
R11379 VSS.n2981 VSS.n1303 146.25
R11380 VSS.n1303 VSS.n1302 146.25
R11381 VSS.n2983 VSS.n2982 146.25
R11382 VSS.n2984 VSS.n2983 146.25
R11383 VSS.n1301 VSS.n1300 146.25
R11384 VSS.n2985 VSS.n1301 146.25
R11385 VSS.n2988 VSS.n2987 146.25
R11386 VSS.n2987 VSS.n2986 146.25
R11387 VSS.n2989 VSS.n1299 146.25
R11388 VSS.n1299 VSS.n1298 146.25
R11389 VSS.n2991 VSS.n2990 146.25
R11390 VSS.n2992 VSS.n2991 146.25
R11391 VSS.n1309 VSS.n1308 146.25
R11392 VSS.n2969 VSS.n1309 146.25
R11393 VSS.n2967 VSS.n2966 146.25
R11394 VSS.n2968 VSS.n2967 146.25
R11395 VSS.n2677 VSS.n2676 146.25
R11396 VSS.n2678 VSS.n2677 146.25
R11397 VSS.n2675 VSS.n1388 146.25
R11398 VSS.n1388 VSS.n1387 146.25
R11399 VSS.n2674 VSS.n2673 146.25
R11400 VSS.n2673 VSS.n2672 146.25
R11401 VSS.n1391 VSS.n1390 146.25
R11402 VSS.n2671 VSS.n1391 146.25
R11403 VSS.n2669 VSS.n2668 146.25
R11404 VSS.n2670 VSS.n2669 146.25
R11405 VSS.n2667 VSS.n1393 146.25
R11406 VSS.n1393 VSS.n1392 146.25
R11407 VSS.n2666 VSS.n2665 146.25
R11408 VSS.n2665 VSS.n2664 146.25
R11409 VSS.n1395 VSS.n1394 146.25
R11410 VSS.n2663 VSS.n1395 146.25
R11411 VSS.n2661 VSS.n2660 146.25
R11412 VSS.n2662 VSS.n2661 146.25
R11413 VSS.n2659 VSS.n1397 146.25
R11414 VSS.n1397 VSS.n1396 146.25
R11415 VSS.n2658 VSS.n2657 146.25
R11416 VSS.n2657 VSS.n2656 146.25
R11417 VSS.n1389 VSS.n1386 146.25
R11418 VSS.n2679 VSS.n1386 146.25
R11419 VSS.n2681 VSS.n1377 146.25
R11420 VSS.n2681 VSS.n2680 146.25
R11421 VSS.n2318 VSS.n2317 146.25
R11422 VSS.n2319 VSS.n2318 146.25
R11423 VSS.n2316 VSS.n2294 146.25
R11424 VSS.n2294 VSS.n2293 146.25
R11425 VSS.n2315 VSS.n2314 146.25
R11426 VSS.n2314 VSS.n2313 146.25
R11427 VSS.n2296 VSS.n2295 146.25
R11428 VSS.n2312 VSS.n2296 146.25
R11429 VSS.n2310 VSS.n2309 146.25
R11430 VSS.n2311 VSS.n2310 146.25
R11431 VSS.n2308 VSS.n2298 146.25
R11432 VSS.n2298 VSS.n2297 146.25
R11433 VSS.n2307 VSS.n2306 146.25
R11434 VSS.n2306 VSS.n2305 146.25
R11435 VSS.n2300 VSS.n2299 146.25
R11436 VSS.n2304 VSS.n2300 146.25
R11437 VSS.n2302 VSS.n2301 146.25
R11438 VSS.n2303 VSS.n2302 146.25
R11439 VSS.n1451 VSS.n1449 146.25
R11440 VSS.n1449 VSS.n1448 146.25
R11441 VSS.n2628 VSS.n2627 146.25
R11442 VSS.n2629 VSS.n2628 146.25
R11443 VSS.n2292 VSS.n2291 146.25
R11444 VSS.n2320 VSS.n2292 146.25
R11445 VSS.n2323 VSS.n2322 146.25
R11446 VSS.n2322 VSS.n2321 146.25
R11447 VSS.n2578 VSS.n2577 146.25
R11448 VSS.n2579 VSS.n2578 146.25
R11449 VSS.n1474 VSS.n1473 146.25
R11450 VSS.n2580 VSS.n1474 146.25
R11451 VSS.n2583 VSS.n2582 146.25
R11452 VSS.n2582 VSS.n2581 146.25
R11453 VSS.n2584 VSS.n1472 146.25
R11454 VSS.n1472 VSS.n1471 146.25
R11455 VSS.n2586 VSS.n2585 146.25
R11456 VSS.n2587 VSS.n2586 146.25
R11457 VSS.n1470 VSS.n1469 146.25
R11458 VSS.n2588 VSS.n1470 146.25
R11459 VSS.n2591 VSS.n2590 146.25
R11460 VSS.n2590 VSS.n2589 146.25
R11461 VSS.n2592 VSS.n1468 146.25
R11462 VSS.n1468 VSS.n1467 146.25
R11463 VSS.n2594 VSS.n2593 146.25
R11464 VSS.n2595 VSS.n2594 146.25
R11465 VSS.n1466 VSS.n1465 146.25
R11466 VSS.n2596 VSS.n1466 146.25
R11467 VSS.n2599 VSS.n2598 146.25
R11468 VSS.n2598 VSS.n2597 146.25
R11469 VSS.n2576 VSS.n1476 146.25
R11470 VSS.n1476 VSS.n1475 146.25
R11471 VSS.n2575 VSS.n2574 146.25
R11472 VSS.n2574 VSS.n2573 146.25
R11473 VSS.n1553 VSS.n1550 146.25
R11474 VSS.n2101 VSS.n1550 146.25
R11475 VSS.n2099 VSS.n2098 146.25
R11476 VSS.n2100 VSS.n2099 146.25
R11477 VSS.n2097 VSS.n1552 146.25
R11478 VSS.n1552 VSS.n1551 146.25
R11479 VSS.n2096 VSS.n2095 146.25
R11480 VSS.n2095 VSS.n2094 146.25
R11481 VSS.n1555 VSS.n1554 146.25
R11482 VSS.n2093 VSS.n1555 146.25
R11483 VSS.n2091 VSS.n2090 146.25
R11484 VSS.n2092 VSS.n2091 146.25
R11485 VSS.n2089 VSS.n1557 146.25
R11486 VSS.n1557 VSS.n1556 146.25
R11487 VSS.n2088 VSS.n2087 146.25
R11488 VSS.n2087 VSS.n2086 146.25
R11489 VSS.n1559 VSS.n1558 146.25
R11490 VSS.n2085 VSS.n1559 146.25
R11491 VSS.n2083 VSS.n2082 146.25
R11492 VSS.n2084 VSS.n2083 146.25
R11493 VSS.n2081 VSS.n1561 146.25
R11494 VSS.n1561 VSS.n1560 146.25
R11495 VSS.n2103 VSS.n1549 146.25
R11496 VSS.n2103 VSS.n2102 146.25
R11497 VSS.n2105 VSS.n2104 146.25
R11498 VSS.n2104 VSS.n1542 146.25
R11499 VSS.n1709 VSS.n1708 146.25
R11500 VSS.n1710 VSS.n1709 146.25
R11501 VSS.n1707 VSS.n1685 146.25
R11502 VSS.n1685 VSS.n1684 146.25
R11503 VSS.n1706 VSS.n1705 146.25
R11504 VSS.n1705 VSS.n1704 146.25
R11505 VSS.n1687 VSS.n1686 146.25
R11506 VSS.n1703 VSS.n1687 146.25
R11507 VSS.n1701 VSS.n1700 146.25
R11508 VSS.n1702 VSS.n1701 146.25
R11509 VSS.n1699 VSS.n1689 146.25
R11510 VSS.n1689 VSS.n1688 146.25
R11511 VSS.n1698 VSS.n1697 146.25
R11512 VSS.n1697 VSS.n1696 146.25
R11513 VSS.n1691 VSS.n1690 146.25
R11514 VSS.n1695 VSS.n1691 146.25
R11515 VSS.n1693 VSS.n1692 146.25
R11516 VSS.n1694 VSS.n1693 146.25
R11517 VSS.n1578 VSS.n1577 146.25
R11518 VSS.n1580 VSS.n1578 146.25
R11519 VSS.n2019 VSS.n2018 146.25
R11520 VSS.n2018 VSS.n2017 146.25
R11521 VSS.n1683 VSS.n1682 146.25
R11522 VSS.n1711 VSS.n1683 146.25
R11523 VSS.n1714 VSS.n1713 146.25
R11524 VSS.n1713 VSS.n1712 146.25
R11525 VSS.n14719 VSS.n14370 142.386
R11526 VSS.n14707 VSS.n14372 142.386
R11527 VSS.n14703 VSS.n14382 142.386
R11528 VSS.n14696 VSS.n14389 142.386
R11529 VSS.n14684 VSS.n14392 142.386
R11530 VSS.n14680 VSS.n14401 142.386
R11531 VSS.n14674 VSS.n14408 142.386
R11532 VSS.n14662 VSS.n14411 142.386
R11533 VSS.n14658 VSS.n14420 142.386
R11534 VSS.n14651 VSS.n14427 142.386
R11535 VSS.n14639 VSS.n14430 142.386
R11536 VSS.n14884 VSS.n14296 142.386
R11537 VSS.n14888 VSS.n14289 142.386
R11538 VSS.n14900 VSS.n14287 142.386
R11539 VSS.n14907 VSS.n14279 142.386
R11540 VSS.n14919 VSS.n14275 142.386
R11541 VSS.n14923 VSS.n14268 142.386
R11542 VSS.n14934 VSS.n14266 142.386
R11543 VSS.n14941 VSS.n14258 142.386
R11544 VSS.n14953 VSS.n14254 142.386
R11545 VSS.n14957 VSS.n14247 142.386
R11546 VSS.n14969 VSS.n14245 142.386
R11547 VSS.n14627 VSS.n14479 142.386
R11548 VSS.n14615 VSS.n14485 142.386
R11549 VSS.n14611 VSS.n14494 142.386
R11550 VSS.n14604 VSS.n14501 142.386
R11551 VSS.n14592 VSS.n14504 142.386
R11552 VSS.n14588 VSS.n14513 142.386
R11553 VSS.n14582 VSS.n14520 142.386
R11554 VSS.n14570 VSS.n14523 142.386
R11555 VSS.n14566 VSS.n14532 142.386
R11556 VSS.n14559 VSS.n14539 142.386
R11557 VSS.n14545 VSS.n14542 142.386
R11558 VSS.n15228 VSS.n15088 142.386
R11559 VSS.n15216 VSS.n15094 142.386
R11560 VSS.n15212 VSS.n15103 142.386
R11561 VSS.n15205 VSS.n15110 142.386
R11562 VSS.n15193 VSS.n15113 142.386
R11563 VSS.n15189 VSS.n15122 142.386
R11564 VSS.n15183 VSS.n15129 142.386
R11565 VSS.n15171 VSS.n15132 142.386
R11566 VSS.n15167 VSS.n15141 142.386
R11567 VSS.n15160 VSS.n15148 142.386
R11568 VSS.n15446 VSS.n14141 142.386
R11569 VSS.n15320 VSS.n14979 142.386
R11570 VSS.n15308 VSS.n14982 142.386
R11571 VSS.n15304 VSS.n14991 142.386
R11572 VSS.n15297 VSS.n14998 142.386
R11573 VSS.n15285 VSS.n15001 142.386
R11574 VSS.n15281 VSS.n15010 142.386
R11575 VSS.n15275 VSS.n15017 142.386
R11576 VSS.n15263 VSS.n15020 142.386
R11577 VSS.n15259 VSS.n15029 142.386
R11578 VSS.n15252 VSS.n15036 142.386
R11579 VSS.n15240 VSS.n15039 142.386
R11580 VSS.n15887 VSS.n15564 142.386
R11581 VSS.n15875 VSS.n15569 142.386
R11582 VSS.n15871 VSS.n15578 142.386
R11583 VSS.n15864 VSS.n15585 142.386
R11584 VSS.n15852 VSS.n15588 142.386
R11585 VSS.n15848 VSS.n15597 142.386
R11586 VSS.n15842 VSS.n15604 142.386
R11587 VSS.n15830 VSS.n15607 142.386
R11588 VSS.n15826 VSS.n15616 142.386
R11589 VSS.n15819 VSS.n15623 142.386
R11590 VSS.n15807 VSS.n15626 142.386
R11591 VSS.n15463 VSS.n14131 142.386
R11592 VSS.n15470 VSS.n14123 142.386
R11593 VSS.n15482 VSS.n14119 142.386
R11594 VSS.n15486 VSS.n14112 142.386
R11595 VSS.n15498 VSS.n14110 142.386
R11596 VSS.n15505 VSS.n14102 142.386
R11597 VSS.n15516 VSS.n14098 142.386
R11598 VSS.n15520 VSS.n14091 142.386
R11599 VSS.n15532 VSS.n14089 142.386
R11600 VSS.n15539 VSS.n14081 142.386
R11601 VSS.n15551 VSS.n14077 142.386
R11602 VSS.n15795 VSS.n15675 142.386
R11603 VSS.n15783 VSS.n15681 142.386
R11604 VSS.n15779 VSS.n15690 142.386
R11605 VSS.n15772 VSS.n15697 142.386
R11606 VSS.n15760 VSS.n15700 142.386
R11607 VSS.n15756 VSS.n15709 142.386
R11608 VSS.n15750 VSS.n15716 142.386
R11609 VSS.n15738 VSS.n15719 142.386
R11610 VSS.n15734 VSS.n15728 142.386
R11611 VSS.n16020 VSS.n14000 142.386
R11612 VSS.n16008 VSS.n14003 142.386
R11613 VSS.n12798 VSS.n12716 142.386
R11614 VSS.n12810 VSS.n12714 142.386
R11615 VSS.n12817 VSS.n12706 142.386
R11616 VSS.n12829 VSS.n12702 142.386
R11617 VSS.n12833 VSS.n12695 142.386
R11618 VSS.n12845 VSS.n12693 142.386
R11619 VSS.n12851 VSS.n12685 142.386
R11620 VSS.n12863 VSS.n12681 142.386
R11621 VSS.n12867 VSS.n12674 142.386
R11622 VSS.n12880 VSS.n12671 142.386
R11623 VSS.n12889 VSS.n12666 142.386
R11624 VSS.n13155 VSS.n12575 142.386
R11625 VSS.n13167 VSS.n12573 142.386
R11626 VSS.n13174 VSS.n12565 142.386
R11627 VSS.n13186 VSS.n12561 142.386
R11628 VSS.n13190 VSS.n12554 142.386
R11629 VSS.n13202 VSS.n12552 142.386
R11630 VSS.n13208 VSS.n12544 142.386
R11631 VSS.n13220 VSS.n12540 142.386
R11632 VSS.n13224 VSS.n12533 142.386
R11633 VSS.n13237 VSS.n12530 142.386
R11634 VSS.n13246 VSS.n12525 142.386
R11635 VSS.n13046 VSS.n12893 142.386
R11636 VSS.n13042 VSS.n12900 142.386
R11637 VSS.n13035 VSS.n12907 142.386
R11638 VSS.n13023 VSS.n12910 142.386
R11639 VSS.n13019 VSS.n12919 142.386
R11640 VSS.n13012 VSS.n12926 142.386
R11641 VSS.n13001 VSS.n12929 142.386
R11642 VSS.n12997 VSS.n12938 142.386
R11643 VSS.n12990 VSS.n12945 142.386
R11644 VSS.n12978 VSS.n12948 142.386
R11645 VSS.n12974 VSS.n12957 142.386
R11646 VSS.n11676 VSS.n11666 142.386
R11647 VSS.n11688 VSS.n11664 142.386
R11648 VSS.n11695 VSS.n11656 142.386
R11649 VSS.n11707 VSS.n11652 142.386
R11650 VSS.n11711 VSS.n11645 142.386
R11651 VSS.n11723 VSS.n11643 142.386
R11652 VSS.n11729 VSS.n11635 142.386
R11653 VSS.n11741 VSS.n11631 142.386
R11654 VSS.n11745 VSS.n11624 142.386
R11655 VSS.n11757 VSS.n11622 142.386
R11656 VSS.n11764 VSS.n11613 142.386
R11657 VSS.n13295 VSS.n13250 142.386
R11658 VSS.n13291 VSS.n13257 142.386
R11659 VSS.n13284 VSS.n13264 142.386
R11660 VSS.n13270 VSS.n13267 142.386
R11661 VSS.n13454 VSS.n11434 142.386
R11662 VSS.n13442 VSS.n11437 142.386
R11663 VSS.n13438 VSS.n11446 142.386
R11664 VSS.n13432 VSS.n11453 142.386
R11665 VSS.n13420 VSS.n11456 142.386
R11666 VSS.n13416 VSS.n11465 142.386
R11667 VSS.n13409 VSS.n11472 142.386
R11668 VSS.n12395 VSS.n11913 142.386
R11669 VSS.n12383 VSS.n11916 142.386
R11670 VSS.n12379 VSS.n11925 142.386
R11671 VSS.n12372 VSS.n11932 142.386
R11672 VSS.n12360 VSS.n11935 142.386
R11673 VSS.n12356 VSS.n11944 142.386
R11674 VSS.n12350 VSS.n11951 142.386
R11675 VSS.n12338 VSS.n11954 142.386
R11676 VSS.n12334 VSS.n11963 142.386
R11677 VSS.n12327 VSS.n11970 142.386
R11678 VSS.n12315 VSS.n11973 142.386
R11679 VSS.n11818 VSS.n11601 142.386
R11680 VSS.n11822 VSS.n11594 142.386
R11681 VSS.n11834 VSS.n11592 142.386
R11682 VSS.n11841 VSS.n11584 142.386
R11683 VSS.n11853 VSS.n11580 142.386
R11684 VSS.n11857 VSS.n11573 142.386
R11685 VSS.n11868 VSS.n11571 142.386
R11686 VSS.n11875 VSS.n11563 142.386
R11687 VSS.n11887 VSS.n11559 142.386
R11688 VSS.n11891 VSS.n11552 142.386
R11689 VSS.n11903 VSS.n11550 142.386
R11690 VSS.n12303 VSS.n11989 142.386
R11691 VSS.n12291 VSS.n11995 142.386
R11692 VSS.n12287 VSS.n12004 142.386
R11693 VSS.n12280 VSS.n12011 142.386
R11694 VSS.n12268 VSS.n12014 142.386
R11695 VSS.n12264 VSS.n12023 142.386
R11696 VSS.n12258 VSS.n12030 142.386
R11697 VSS.n12246 VSS.n12033 142.386
R11698 VSS.n12242 VSS.n12042 142.386
R11699 VSS.n12235 VSS.n12049 142.386
R11700 VSS.n12223 VSS.n12052 142.386
R11701 VSS.n7833 VSS.n7677 142.386
R11702 VSS.n7821 VSS.n7679 142.386
R11703 VSS.n7817 VSS.n7689 142.386
R11704 VSS.n7810 VSS.n7696 142.386
R11705 VSS.n7798 VSS.n7699 142.386
R11706 VSS.n7794 VSS.n7708 142.386
R11707 VSS.n7788 VSS.n7715 142.386
R11708 VSS.n7776 VSS.n7718 142.386
R11709 VSS.n7772 VSS.n7727 142.386
R11710 VSS.n7765 VSS.n7734 142.386
R11711 VSS.n7753 VSS.n7737 142.386
R11712 VSS.n8177 VSS.n8020 142.386
R11713 VSS.n8173 VSS.n8031 142.386
R11714 VSS.n8161 VSS.n8033 142.386
R11715 VSS.n8157 VSS.n8043 142.386
R11716 VSS.n8150 VSS.n8050 142.386
R11717 VSS.n8138 VSS.n8053 142.386
R11718 VSS.n8134 VSS.n8062 142.386
R11719 VSS.n8128 VSS.n8069 142.386
R11720 VSS.n8116 VSS.n8072 142.386
R11721 VSS.n8112 VSS.n8081 142.386
R11722 VSS.n8105 VSS.n8088 142.386
R11723 VSS.n7929 VSS.n7595 142.386
R11724 VSS.n7933 VSS.n7588 142.386
R11725 VSS.n7945 VSS.n7586 142.386
R11726 VSS.n7952 VSS.n7578 142.386
R11727 VSS.n7964 VSS.n7574 142.386
R11728 VSS.n7968 VSS.n7567 142.386
R11729 VSS.n7979 VSS.n7565 142.386
R11730 VSS.n7986 VSS.n7557 142.386
R11731 VSS.n7998 VSS.n7553 142.386
R11732 VSS.n8002 VSS.n7546 142.386
R11733 VSS.n8014 VSS.n7544 142.386
R11734 VSS.n8535 VSS.n8378 142.386
R11735 VSS.n8531 VSS.n8389 142.386
R11736 VSS.n8519 VSS.n8391 142.386
R11737 VSS.n8515 VSS.n8401 142.386
R11738 VSS.n8508 VSS.n8408 142.386
R11739 VSS.n8496 VSS.n8411 142.386
R11740 VSS.n8492 VSS.n8420 142.386
R11741 VSS.n8486 VSS.n8427 142.386
R11742 VSS.n8474 VSS.n8430 142.386
R11743 VSS.n8470 VSS.n8439 142.386
R11744 VSS.n8463 VSS.n8446 142.386
R11745 VSS.n8287 VSS.n7455 142.386
R11746 VSS.n8291 VSS.n7448 142.386
R11747 VSS.n8303 VSS.n7446 142.386
R11748 VSS.n8310 VSS.n7438 142.386
R11749 VSS.n8322 VSS.n7434 142.386
R11750 VSS.n8326 VSS.n7427 142.386
R11751 VSS.n8337 VSS.n7425 142.386
R11752 VSS.n8344 VSS.n7417 142.386
R11753 VSS.n8356 VSS.n7413 142.386
R11754 VSS.n8360 VSS.n7406 142.386
R11755 VSS.n8372 VSS.n7404 142.386
R11756 VSS.n8757 VSS.n8736 142.386
R11757 VSS.n8753 VSS.n8750 142.386
R11758 VSS.n8926 VSS.n6906 142.386
R11759 VSS.n8914 VSS.n6909 142.386
R11760 VSS.n8910 VSS.n6918 142.386
R11761 VSS.n8903 VSS.n6925 142.386
R11762 VSS.n8892 VSS.n6928 142.386
R11763 VSS.n8888 VSS.n6937 142.386
R11764 VSS.n8881 VSS.n6944 142.386
R11765 VSS.n8869 VSS.n6947 142.386
R11766 VSS.n8865 VSS.n6956 142.386
R11767 VSS.n8645 VSS.n7315 142.386
R11768 VSS.n8649 VSS.n7308 142.386
R11769 VSS.n8661 VSS.n7306 142.386
R11770 VSS.n8668 VSS.n7298 142.386
R11771 VSS.n8680 VSS.n7294 142.386
R11772 VSS.n8684 VSS.n7287 142.386
R11773 VSS.n8695 VSS.n7285 142.386
R11774 VSS.n8702 VSS.n7277 142.386
R11775 VSS.n8714 VSS.n7273 142.386
R11776 VSS.n8718 VSS.n7266 142.386
R11777 VSS.n8730 VSS.n7264 142.386
R11778 VSS.n7079 VSS.n7066 142.386
R11779 VSS.n7086 VSS.n7058 142.386
R11780 VSS.n7098 VSS.n7054 142.386
R11781 VSS.n7102 VSS.n7047 142.386
R11782 VSS.n7114 VSS.n7045 142.386
R11783 VSS.n7121 VSS.n7037 142.386
R11784 VSS.n7132 VSS.n7033 142.386
R11785 VSS.n7136 VSS.n7026 142.386
R11786 VSS.n7148 VSS.n7024 142.386
R11787 VSS.n7155 VSS.n7016 142.386
R11788 VSS.n7167 VSS.n7012 142.386
R11789 VSS.n4251 VSS.n4169 142.386
R11790 VSS.n4263 VSS.n4167 142.386
R11791 VSS.n4270 VSS.n4159 142.386
R11792 VSS.n4282 VSS.n4155 142.386
R11793 VSS.n4286 VSS.n4148 142.386
R11794 VSS.n4298 VSS.n4146 142.386
R11795 VSS.n4304 VSS.n4138 142.386
R11796 VSS.n4316 VSS.n4134 142.386
R11797 VSS.n4320 VSS.n4127 142.386
R11798 VSS.n4333 VSS.n4124 142.386
R11799 VSS.n4342 VSS.n4119 142.386
R11800 VSS.n4608 VSS.n4028 142.386
R11801 VSS.n4620 VSS.n4026 142.386
R11802 VSS.n4627 VSS.n4018 142.386
R11803 VSS.n4639 VSS.n4014 142.386
R11804 VSS.n4643 VSS.n4007 142.386
R11805 VSS.n4655 VSS.n4005 142.386
R11806 VSS.n4661 VSS.n3997 142.386
R11807 VSS.n4673 VSS.n3993 142.386
R11808 VSS.n4677 VSS.n3986 142.386
R11809 VSS.n4690 VSS.n3983 142.386
R11810 VSS.n4699 VSS.n3978 142.386
R11811 VSS.n4499 VSS.n4346 142.386
R11812 VSS.n4495 VSS.n4353 142.386
R11813 VSS.n4488 VSS.n4360 142.386
R11814 VSS.n4476 VSS.n4363 142.386
R11815 VSS.n4472 VSS.n4372 142.386
R11816 VSS.n4465 VSS.n4379 142.386
R11817 VSS.n4454 VSS.n4382 142.386
R11818 VSS.n4450 VSS.n4391 142.386
R11819 VSS.n4443 VSS.n4398 142.386
R11820 VSS.n4431 VSS.n4401 142.386
R11821 VSS.n4427 VSS.n4410 142.386
R11822 VSS.n4965 VSS.n3887 142.386
R11823 VSS.n4977 VSS.n3885 142.386
R11824 VSS.n4984 VSS.n3877 142.386
R11825 VSS.n4996 VSS.n3873 142.386
R11826 VSS.n5000 VSS.n3866 142.386
R11827 VSS.n5012 VSS.n3864 142.386
R11828 VSS.n5018 VSS.n3856 142.386
R11829 VSS.n5030 VSS.n3852 142.386
R11830 VSS.n5034 VSS.n3845 142.386
R11831 VSS.n5047 VSS.n3842 142.386
R11832 VSS.n5056 VSS.n3837 142.386
R11833 VSS.n4856 VSS.n4703 142.386
R11834 VSS.n4852 VSS.n4710 142.386
R11835 VSS.n4845 VSS.n4717 142.386
R11836 VSS.n4833 VSS.n4720 142.386
R11837 VSS.n4829 VSS.n4729 142.386
R11838 VSS.n4822 VSS.n4736 142.386
R11839 VSS.n4811 VSS.n4739 142.386
R11840 VSS.n4807 VSS.n4748 142.386
R11841 VSS.n4800 VSS.n4755 142.386
R11842 VSS.n4788 VSS.n4758 142.386
R11843 VSS.n4784 VSS.n4767 142.386
R11844 VSS.n5322 VSS.n3746 142.386
R11845 VSS.n5334 VSS.n3744 142.386
R11846 VSS.n5341 VSS.n3736 142.386
R11847 VSS.n5353 VSS.n3732 142.386
R11848 VSS.n5357 VSS.n3725 142.386
R11849 VSS.n5369 VSS.n3723 142.386
R11850 VSS.n5375 VSS.n3715 142.386
R11851 VSS.n5387 VSS.n3711 142.386
R11852 VSS.n5391 VSS.n3704 142.386
R11853 VSS.n5404 VSS.n3701 142.386
R11854 VSS.n5413 VSS.n3696 142.386
R11855 VSS.n5213 VSS.n5060 142.386
R11856 VSS.n5209 VSS.n5067 142.386
R11857 VSS.n5202 VSS.n5074 142.386
R11858 VSS.n5190 VSS.n5077 142.386
R11859 VSS.n5186 VSS.n5086 142.386
R11860 VSS.n5179 VSS.n5093 142.386
R11861 VSS.n5168 VSS.n5096 142.386
R11862 VSS.n5164 VSS.n5105 142.386
R11863 VSS.n5157 VSS.n5112 142.386
R11864 VSS.n5145 VSS.n5115 142.386
R11865 VSS.n5141 VSS.n5124 142.386
R11866 VSS.n5559 VSS.n5417 142.386
R11867 VSS.n5555 VSS.n5424 142.386
R11868 VSS.n5548 VSS.n5431 142.386
R11869 VSS.n5536 VSS.n5434 142.386
R11870 VSS.n5532 VSS.n5443 142.386
R11871 VSS.n5525 VSS.n5450 142.386
R11872 VSS.n5514 VSS.n5453 142.386
R11873 VSS.n5510 VSS.n5462 142.386
R11874 VSS.n5503 VSS.n5469 142.386
R11875 VSS.n5491 VSS.n5472 142.386
R11876 VSS.n5487 VSS.n5481 142.386
R11877 VSS.n1960 VSS.n1611 142.386
R11878 VSS.n1948 VSS.n1613 142.386
R11879 VSS.n1944 VSS.n1623 142.386
R11880 VSS.n1937 VSS.n1630 142.386
R11881 VSS.n1925 VSS.n1633 142.386
R11882 VSS.n1921 VSS.n1642 142.386
R11883 VSS.n1915 VSS.n1649 142.386
R11884 VSS.n1903 VSS.n1652 142.386
R11885 VSS.n1899 VSS.n1661 142.386
R11886 VSS.n1892 VSS.n1668 142.386
R11887 VSS.n1880 VSS.n1671 142.386
R11888 VSS.n2125 VSS.n1537 142.386
R11889 VSS.n2129 VSS.n1530 142.386
R11890 VSS.n2141 VSS.n1528 142.386
R11891 VSS.n2148 VSS.n1520 142.386
R11892 VSS.n2160 VSS.n1516 142.386
R11893 VSS.n2164 VSS.n1509 142.386
R11894 VSS.n2175 VSS.n1507 142.386
R11895 VSS.n2182 VSS.n1499 142.386
R11896 VSS.n2194 VSS.n1495 142.386
R11897 VSS.n2198 VSS.n1488 142.386
R11898 VSS.n2210 VSS.n1486 142.386
R11899 VSS.n1868 VSS.n1720 142.386
R11900 VSS.n1856 VSS.n1726 142.386
R11901 VSS.n1852 VSS.n1735 142.386
R11902 VSS.n1845 VSS.n1742 142.386
R11903 VSS.n1833 VSS.n1745 142.386
R11904 VSS.n1829 VSS.n1754 142.386
R11905 VSS.n1823 VSS.n1761 142.386
R11906 VSS.n1811 VSS.n1764 142.386
R11907 VSS.n1807 VSS.n1773 142.386
R11908 VSS.n1800 VSS.n1780 142.386
R11909 VSS.n1786 VSS.n1783 142.386
R11910 VSS.n2469 VSS.n2329 142.386
R11911 VSS.n2457 VSS.n2335 142.386
R11912 VSS.n2453 VSS.n2344 142.386
R11913 VSS.n2446 VSS.n2351 142.386
R11914 VSS.n2434 VSS.n2354 142.386
R11915 VSS.n2430 VSS.n2363 142.386
R11916 VSS.n2424 VSS.n2370 142.386
R11917 VSS.n2412 VSS.n2373 142.386
R11918 VSS.n2408 VSS.n2382 142.386
R11919 VSS.n2401 VSS.n2389 142.386
R11920 VSS.n2687 VSS.n1382 142.386
R11921 VSS.n2561 VSS.n2220 142.386
R11922 VSS.n2549 VSS.n2223 142.386
R11923 VSS.n2545 VSS.n2232 142.386
R11924 VSS.n2538 VSS.n2239 142.386
R11925 VSS.n2526 VSS.n2242 142.386
R11926 VSS.n2522 VSS.n2251 142.386
R11927 VSS.n2516 VSS.n2258 142.386
R11928 VSS.n2504 VSS.n2261 142.386
R11929 VSS.n2500 VSS.n2270 142.386
R11930 VSS.n2493 VSS.n2277 142.386
R11931 VSS.n2481 VSS.n2280 142.386
R11932 VSS.n2704 VSS.n1372 142.386
R11933 VSS.n2711 VSS.n1364 142.386
R11934 VSS.n2723 VSS.n1360 142.386
R11935 VSS.n2727 VSS.n1353 142.386
R11936 VSS.n2739 VSS.n1351 142.386
R11937 VSS.n2746 VSS.n1343 142.386
R11938 VSS.n2757 VSS.n1339 142.386
R11939 VSS.n2761 VSS.n1332 142.386
R11940 VSS.n2773 VSS.n1330 142.386
R11941 VSS.n2780 VSS.n1322 142.386
R11942 VSS.n2792 VSS.n1318 142.386
R11943 VSS.n2961 VSS.n2805 142.386
R11944 VSS.n2949 VSS.n2810 142.386
R11945 VSS.n2945 VSS.n2819 142.386
R11946 VSS.n2938 VSS.n2826 142.386
R11947 VSS.n2926 VSS.n2829 142.386
R11948 VSS.n2922 VSS.n2838 142.386
R11949 VSS.n2916 VSS.n2845 142.386
R11950 VSS.n2904 VSS.n2848 142.386
R11951 VSS.n2900 VSS.n2857 142.386
R11952 VSS.n2893 VSS.n2864 142.386
R11953 VSS.n2881 VSS.n2867 142.386
R11954 sky130_asc_nfet_01v8_lvt_9_0/SOURCE VSS.t0 137.313
R11955 VSS.n1267 VSS.t13 130.913
R11956 VSS.n17658 sky130_asc_nfet_01v8_lvt_1_0/SOURCE 130.062
R11957 VSS.n15996 VSS.n14012 126.781
R11958 VSS.n12211 VSS.n12061 126.781
R11959 VSS.n7010 VSS.n7004 126.781
R11960 VSS.n6802 VSS.n6772 126.781
R11961 VSS.n5656 VSS.n3640 126.781
R11962 VSS.n3043 VSS.n1271 126.781
R11963 VSS.n10436 VSS.n10434 126.563
R11964 VSS.n10433 VSS.n10432 126.563
R11965 VSS.n14727 VSS.n14363 124.831
R11966 VSS.n12788 VSS.n12723 124.831
R11967 VSS.n7672 VSS.n7670 124.831
R11968 VSS.n6830 VSS.n6757 124.831
R11969 VSS.n4241 VSS.n4176 124.831
R11970 VSS.n1968 VSS.n1604 124.831
R11971 VSS.n10438 VSS.n10437 123.662
R11972 VSS.n14338 VSS.n14334 97.524
R11973 VSS.n15361 VSS.n14222 97.524
R11974 VSS.n14833 VSS.n14324 97.524
R11975 VSS.n14192 VSS.n14158 97.524
R11976 VSS.n14209 VSS.n14205 97.524
R11977 VSS.n15921 VSS.n14055 97.524
R11978 VSS.n14042 VSS.n14038 97.524
R11979 VSS.n12644 VSS.n12640 97.524
R11980 VSS.n12503 VSS.n12499 97.524
R11981 VSS.n12627 VSS.n12598 97.524
R11982 VSS.n12457 VSS.n11513 97.524
R11983 VSS.n12486 VSS.n11497 97.524
R11984 VSS.n12136 VSS.n11527 97.524
R11985 VSS.n12091 VSS.n12087 97.524
R11986 VSS.n7645 VSS.n7616 97.524
R11987 VSS.n7505 VSS.n7476 97.524
R11988 VSS.n7522 VSS.n7518 97.524
R11989 VSS.n7365 VSS.n7336 97.524
R11990 VSS.n7382 VSS.n7378 97.524
R11991 VSS.n7242 VSS.n7238 97.524
R11992 VSS.n7225 VSS.n6980 97.524
R11993 VSS.n4097 VSS.n4093 97.524
R11994 VSS.n3956 VSS.n3952 97.524
R11995 VSS.n4080 VSS.n4051 97.524
R11996 VSS.n3815 VSS.n3811 97.524
R11997 VSS.n3939 VSS.n3910 97.524
R11998 VSS.n3798 VSS.n3769 97.524
R11999 VSS.n3674 VSS.n3670 97.524
R12000 VSS.n1579 VSS.n1575 97.524
R12001 VSS.n2602 VSS.n1463 97.524
R12002 VSS.n2074 VSS.n1565 97.524
R12003 VSS.n1433 VSS.n1399 97.524
R12004 VSS.n1450 VSS.n1446 97.524
R12005 VSS.n2995 VSS.n1296 97.524
R12006 VSS.n16035 VSS.n16029 92.501
R12007 VSS.n17224 VSS.n16074 92.501
R12008 VSS.n17134 VSS.n16164 92.501
R12009 VSS.n17044 VSS.n16254 92.501
R12010 VSS.n16954 VSS.n16344 92.501
R12011 VSS.n16864 VSS.n16434 92.501
R12012 VSS.n16774 VSS.n16524 92.501
R12013 VSS.n16684 VSS.n16614 92.501
R12014 VSS.n11180 VSS.n11081 92.501
R12015 VSS.n11270 VSS.n10991 92.501
R12016 VSS.n11360 VSS.n10901 92.501
R12017 VSS.n13479 VSS.n10811 92.501
R12018 VSS.n13570 VSS.n10721 92.501
R12019 VSS.n13660 VSS.n10631 92.501
R12020 VSS.n13750 VSS.n10541 92.501
R12021 VSS.n13954 VSS.n10496 92.501
R12022 VSS.n10179 VSS.n9209 92.501
R12023 VSS.n10089 VSS.n9299 92.501
R12024 VSS.n9999 VSS.n9389 92.501
R12025 VSS.n9909 VSS.n9479 92.501
R12026 VSS.n9819 VSS.n9569 92.501
R12027 VSS.n9729 VSS.n9659 92.501
R12028 VSS.n9178 VSS.n8934 92.501
R12029 VSS.n5733 VSS.n3581 92.501
R12030 VSS.n5855 VSS.n3523 92.501
R12031 VSS.n5977 VSS.n3465 92.501
R12032 VSS.n6099 VSS.n3407 92.501
R12033 VSS.n6221 VSS.n3349 92.501
R12034 VSS.n6343 VSS.n3291 92.501
R12035 VSS.n6465 VSS.n3233 92.501
R12036 VSS.n6535 VSS.n3145 92.501
R12037 VSS.n1177 VSS.n26 92.501
R12038 VSS.n1087 VSS.n117 92.501
R12039 VSS.n997 VSS.n207 92.501
R12040 VSS.n907 VSS.n297 92.501
R12041 VSS.n817 VSS.n387 92.501
R12042 VSS.n727 VSS.n477 92.501
R12043 VSS.n637 VSS.n567 92.501
R12044 VSS.n17351 VSS.n17350 92.5
R12045 VSS.n17337 VSS.n17336 92.5
R12046 VSS.n17339 VSS.n17338 92.5
R12047 VSS.n17341 VSS.n17340 92.5
R12048 VSS.n17343 VSS.n17342 92.5
R12049 VSS.n17345 VSS.n17344 92.5
R12050 VSS.n17347 VSS.n17346 92.5
R12051 VSS.n17349 VSS.n17348 92.5
R12052 VSS.n17335 VSS.n16030 92.5
R12053 VSS.t30 VSS.n16030 92.5
R12054 VSS.n17366 VSS.n17365 92.5
R12055 VSS.n17364 VSS.n17363 92.5
R12056 VSS.n17362 VSS.n17361 92.5
R12057 VSS.n17360 VSS.n17359 92.5
R12058 VSS.n17358 VSS.n17357 92.5
R12059 VSS.n17356 VSS.n17355 92.5
R12060 VSS.n17354 VSS.n17353 92.5
R12061 VSS.n17352 VSS.n17321 92.5
R12062 VSS.t30 VSS.n17321 92.5
R12063 VSS.n17368 VSS.n17367 92.5
R12064 VSS.n17370 VSS.n17369 92.5
R12065 VSS.n17372 VSS.n17371 92.5
R12066 VSS.n17374 VSS.n17373 92.5
R12067 VSS.n17376 VSS.n17375 92.5
R12068 VSS.n17378 VSS.n17377 92.5
R12069 VSS.n17380 VSS.n17379 92.5
R12070 VSS.n17381 VSS.n17326 92.5
R12071 VSS.n17383 VSS.n17382 92.5
R12072 VSS.n17330 VSS.n17313 92.5
R12073 VSS.t30 VSS.n17313 92.5
R12074 VSS.n16029 VSS.n16027 92.5
R12075 VSS.n17385 VSS.n17312 92.5
R12076 VSS.n17394 VSS.n16034 92.5
R12077 VSS.n17456 VSS.n16037 92.5
R12078 VSS.n17447 VSS.n16033 92.5
R12079 VSS.n17404 VSS.n16038 92.5
R12080 VSS.n17408 VSS.n16032 92.5
R12081 VSS.n17412 VSS.n16039 92.5
R12082 VSS.n17415 VSS.n16031 92.5
R12083 VSS.n16107 VSS.n16106 92.5
R12084 VSS.n16056 VSS.n16054 92.5
R12085 VSS.n16095 VSS.n16094 92.5
R12086 VSS.n16097 VSS.n16096 92.5
R12087 VSS.n16099 VSS.n16098 92.5
R12088 VSS.n16101 VSS.n16100 92.5
R12089 VSS.n16103 VSS.n16102 92.5
R12090 VSS.n16105 VSS.n16104 92.5
R12091 VSS.n17308 VSS.n17307 92.5
R12092 VSS.n17307 VSS.t54 92.5
R12093 VSS.n16122 VSS.n16121 92.5
R12094 VSS.n16120 VSS.n16119 92.5
R12095 VSS.n16118 VSS.n16117 92.5
R12096 VSS.n16116 VSS.n16115 92.5
R12097 VSS.n16114 VSS.n16113 92.5
R12098 VSS.n16112 VSS.n16111 92.5
R12099 VSS.n16110 VSS.n16109 92.5
R12100 VSS.n16108 VSS.n16065 92.5
R12101 VSS.t54 VSS.n16065 92.5
R12102 VSS.n16124 VSS.n16123 92.5
R12103 VSS.n16126 VSS.n16125 92.5
R12104 VSS.n16128 VSS.n16127 92.5
R12105 VSS.n16130 VSS.n16129 92.5
R12106 VSS.n16132 VSS.n16131 92.5
R12107 VSS.n16134 VSS.n16133 92.5
R12108 VSS.n16136 VSS.n16135 92.5
R12109 VSS.n16138 VSS.n16137 92.5
R12110 VSS.n16140 VSS.n16139 92.5
R12111 VSS.n16141 VSS.n16057 92.5
R12112 VSS.t54 VSS.n16057 92.5
R12113 VSS.n17225 VSS.n17224 92.5
R12114 VSS.n17300 VSS.n16076 92.5
R12115 VSS.n17291 VSS.n16073 92.5
R12116 VSS.n17235 VSS.n16077 92.5
R12117 VSS.n17239 VSS.n16072 92.5
R12118 VSS.n17243 VSS.n16078 92.5
R12119 VSS.n17247 VSS.n16071 92.5
R12120 VSS.n17306 VSS.n16081 92.5
R12121 VSS.n17253 VSS.n16075 92.5
R12122 VSS.n16197 VSS.n16196 92.5
R12123 VSS.n16146 VSS.n16144 92.5
R12124 VSS.n16185 VSS.n16184 92.5
R12125 VSS.n16187 VSS.n16186 92.5
R12126 VSS.n16189 VSS.n16188 92.5
R12127 VSS.n16191 VSS.n16190 92.5
R12128 VSS.n16193 VSS.n16192 92.5
R12129 VSS.n16195 VSS.n16194 92.5
R12130 VSS.n17218 VSS.n17217 92.5
R12131 VSS.n17217 VSS.t50 92.5
R12132 VSS.n16212 VSS.n16211 92.5
R12133 VSS.n16210 VSS.n16209 92.5
R12134 VSS.n16208 VSS.n16207 92.5
R12135 VSS.n16206 VSS.n16205 92.5
R12136 VSS.n16204 VSS.n16203 92.5
R12137 VSS.n16202 VSS.n16201 92.5
R12138 VSS.n16200 VSS.n16199 92.5
R12139 VSS.n16198 VSS.n16155 92.5
R12140 VSS.t50 VSS.n16155 92.5
R12141 VSS.n16214 VSS.n16213 92.5
R12142 VSS.n16216 VSS.n16215 92.5
R12143 VSS.n16218 VSS.n16217 92.5
R12144 VSS.n16220 VSS.n16219 92.5
R12145 VSS.n16222 VSS.n16221 92.5
R12146 VSS.n16224 VSS.n16223 92.5
R12147 VSS.n16226 VSS.n16225 92.5
R12148 VSS.n16228 VSS.n16227 92.5
R12149 VSS.n16230 VSS.n16229 92.5
R12150 VSS.n16231 VSS.n16147 92.5
R12151 VSS.t50 VSS.n16147 92.5
R12152 VSS.n17135 VSS.n17134 92.5
R12153 VSS.n17210 VSS.n16166 92.5
R12154 VSS.n17201 VSS.n16163 92.5
R12155 VSS.n17145 VSS.n16167 92.5
R12156 VSS.n17149 VSS.n16162 92.5
R12157 VSS.n17153 VSS.n16168 92.5
R12158 VSS.n17157 VSS.n16161 92.5
R12159 VSS.n17216 VSS.n16171 92.5
R12160 VSS.n17163 VSS.n16165 92.5
R12161 VSS.n16287 VSS.n16286 92.5
R12162 VSS.n16236 VSS.n16234 92.5
R12163 VSS.n16275 VSS.n16274 92.5
R12164 VSS.n16277 VSS.n16276 92.5
R12165 VSS.n16279 VSS.n16278 92.5
R12166 VSS.n16281 VSS.n16280 92.5
R12167 VSS.n16283 VSS.n16282 92.5
R12168 VSS.n16285 VSS.n16284 92.5
R12169 VSS.n17128 VSS.n17127 92.5
R12170 VSS.n17127 VSS.t42 92.5
R12171 VSS.n16302 VSS.n16301 92.5
R12172 VSS.n16300 VSS.n16299 92.5
R12173 VSS.n16298 VSS.n16297 92.5
R12174 VSS.n16296 VSS.n16295 92.5
R12175 VSS.n16294 VSS.n16293 92.5
R12176 VSS.n16292 VSS.n16291 92.5
R12177 VSS.n16290 VSS.n16289 92.5
R12178 VSS.n16288 VSS.n16245 92.5
R12179 VSS.t42 VSS.n16245 92.5
R12180 VSS.n16304 VSS.n16303 92.5
R12181 VSS.n16306 VSS.n16305 92.5
R12182 VSS.n16308 VSS.n16307 92.5
R12183 VSS.n16310 VSS.n16309 92.5
R12184 VSS.n16312 VSS.n16311 92.5
R12185 VSS.n16314 VSS.n16313 92.5
R12186 VSS.n16316 VSS.n16315 92.5
R12187 VSS.n16318 VSS.n16317 92.5
R12188 VSS.n16320 VSS.n16319 92.5
R12189 VSS.n16321 VSS.n16237 92.5
R12190 VSS.t42 VSS.n16237 92.5
R12191 VSS.n17045 VSS.n17044 92.5
R12192 VSS.n17120 VSS.n16256 92.5
R12193 VSS.n17111 VSS.n16253 92.5
R12194 VSS.n17055 VSS.n16257 92.5
R12195 VSS.n17059 VSS.n16252 92.5
R12196 VSS.n17063 VSS.n16258 92.5
R12197 VSS.n17067 VSS.n16251 92.5
R12198 VSS.n17126 VSS.n16261 92.5
R12199 VSS.n17073 VSS.n16255 92.5
R12200 VSS.n16377 VSS.n16376 92.5
R12201 VSS.n16326 VSS.n16324 92.5
R12202 VSS.n16365 VSS.n16364 92.5
R12203 VSS.n16367 VSS.n16366 92.5
R12204 VSS.n16369 VSS.n16368 92.5
R12205 VSS.n16371 VSS.n16370 92.5
R12206 VSS.n16373 VSS.n16372 92.5
R12207 VSS.n16375 VSS.n16374 92.5
R12208 VSS.n17038 VSS.n17037 92.5
R12209 VSS.n17037 VSS.t68 92.5
R12210 VSS.n16392 VSS.n16391 92.5
R12211 VSS.n16390 VSS.n16389 92.5
R12212 VSS.n16388 VSS.n16387 92.5
R12213 VSS.n16386 VSS.n16385 92.5
R12214 VSS.n16384 VSS.n16383 92.5
R12215 VSS.n16382 VSS.n16381 92.5
R12216 VSS.n16380 VSS.n16379 92.5
R12217 VSS.n16378 VSS.n16335 92.5
R12218 VSS.t68 VSS.n16335 92.5
R12219 VSS.n16394 VSS.n16393 92.5
R12220 VSS.n16396 VSS.n16395 92.5
R12221 VSS.n16398 VSS.n16397 92.5
R12222 VSS.n16400 VSS.n16399 92.5
R12223 VSS.n16402 VSS.n16401 92.5
R12224 VSS.n16404 VSS.n16403 92.5
R12225 VSS.n16406 VSS.n16405 92.5
R12226 VSS.n16408 VSS.n16407 92.5
R12227 VSS.n16410 VSS.n16409 92.5
R12228 VSS.n16411 VSS.n16327 92.5
R12229 VSS.t68 VSS.n16327 92.5
R12230 VSS.n16955 VSS.n16954 92.5
R12231 VSS.n17030 VSS.n16346 92.5
R12232 VSS.n17021 VSS.n16343 92.5
R12233 VSS.n16965 VSS.n16347 92.5
R12234 VSS.n16969 VSS.n16342 92.5
R12235 VSS.n16973 VSS.n16348 92.5
R12236 VSS.n16977 VSS.n16341 92.5
R12237 VSS.n17036 VSS.n16351 92.5
R12238 VSS.n16983 VSS.n16345 92.5
R12239 VSS.n16467 VSS.n16466 92.5
R12240 VSS.n16416 VSS.n16414 92.5
R12241 VSS.n16455 VSS.n16454 92.5
R12242 VSS.n16457 VSS.n16456 92.5
R12243 VSS.n16459 VSS.n16458 92.5
R12244 VSS.n16461 VSS.n16460 92.5
R12245 VSS.n16463 VSS.n16462 92.5
R12246 VSS.n16465 VSS.n16464 92.5
R12247 VSS.n16948 VSS.n16947 92.5
R12248 VSS.n16947 VSS.t74 92.5
R12249 VSS.n16482 VSS.n16481 92.5
R12250 VSS.n16480 VSS.n16479 92.5
R12251 VSS.n16478 VSS.n16477 92.5
R12252 VSS.n16476 VSS.n16475 92.5
R12253 VSS.n16474 VSS.n16473 92.5
R12254 VSS.n16472 VSS.n16471 92.5
R12255 VSS.n16470 VSS.n16469 92.5
R12256 VSS.n16468 VSS.n16425 92.5
R12257 VSS.t74 VSS.n16425 92.5
R12258 VSS.n16484 VSS.n16483 92.5
R12259 VSS.n16486 VSS.n16485 92.5
R12260 VSS.n16488 VSS.n16487 92.5
R12261 VSS.n16490 VSS.n16489 92.5
R12262 VSS.n16492 VSS.n16491 92.5
R12263 VSS.n16494 VSS.n16493 92.5
R12264 VSS.n16496 VSS.n16495 92.5
R12265 VSS.n16498 VSS.n16497 92.5
R12266 VSS.n16500 VSS.n16499 92.5
R12267 VSS.n16501 VSS.n16417 92.5
R12268 VSS.t74 VSS.n16417 92.5
R12269 VSS.n16865 VSS.n16864 92.5
R12270 VSS.n16940 VSS.n16436 92.5
R12271 VSS.n16931 VSS.n16433 92.5
R12272 VSS.n16875 VSS.n16437 92.5
R12273 VSS.n16879 VSS.n16432 92.5
R12274 VSS.n16883 VSS.n16438 92.5
R12275 VSS.n16887 VSS.n16431 92.5
R12276 VSS.n16946 VSS.n16441 92.5
R12277 VSS.n16893 VSS.n16435 92.5
R12278 VSS.n16557 VSS.n16556 92.5
R12279 VSS.n16506 VSS.n16504 92.5
R12280 VSS.n16545 VSS.n16544 92.5
R12281 VSS.n16547 VSS.n16546 92.5
R12282 VSS.n16549 VSS.n16548 92.5
R12283 VSS.n16551 VSS.n16550 92.5
R12284 VSS.n16553 VSS.n16552 92.5
R12285 VSS.n16555 VSS.n16554 92.5
R12286 VSS.n16858 VSS.n16857 92.5
R12287 VSS.n16857 VSS.t90 92.5
R12288 VSS.n16572 VSS.n16571 92.5
R12289 VSS.n16570 VSS.n16569 92.5
R12290 VSS.n16568 VSS.n16567 92.5
R12291 VSS.n16566 VSS.n16565 92.5
R12292 VSS.n16564 VSS.n16563 92.5
R12293 VSS.n16562 VSS.n16561 92.5
R12294 VSS.n16560 VSS.n16559 92.5
R12295 VSS.n16558 VSS.n16515 92.5
R12296 VSS.t90 VSS.n16515 92.5
R12297 VSS.n16574 VSS.n16573 92.5
R12298 VSS.n16576 VSS.n16575 92.5
R12299 VSS.n16578 VSS.n16577 92.5
R12300 VSS.n16580 VSS.n16579 92.5
R12301 VSS.n16582 VSS.n16581 92.5
R12302 VSS.n16584 VSS.n16583 92.5
R12303 VSS.n16586 VSS.n16585 92.5
R12304 VSS.n16588 VSS.n16587 92.5
R12305 VSS.n16590 VSS.n16589 92.5
R12306 VSS.n16591 VSS.n16507 92.5
R12307 VSS.t90 VSS.n16507 92.5
R12308 VSS.n16775 VSS.n16774 92.5
R12309 VSS.n16850 VSS.n16526 92.5
R12310 VSS.n16841 VSS.n16523 92.5
R12311 VSS.n16785 VSS.n16527 92.5
R12312 VSS.n16789 VSS.n16522 92.5
R12313 VSS.n16793 VSS.n16528 92.5
R12314 VSS.n16797 VSS.n16521 92.5
R12315 VSS.n16856 VSS.n16531 92.5
R12316 VSS.n16803 VSS.n16525 92.5
R12317 VSS.n16647 VSS.n16646 92.5
R12318 VSS.n16596 VSS.n16594 92.5
R12319 VSS.n16635 VSS.n16634 92.5
R12320 VSS.n16637 VSS.n16636 92.5
R12321 VSS.n16639 VSS.n16638 92.5
R12322 VSS.n16641 VSS.n16640 92.5
R12323 VSS.n16643 VSS.n16642 92.5
R12324 VSS.n16645 VSS.n16644 92.5
R12325 VSS.n16768 VSS.n16767 92.5
R12326 VSS.n16767 VSS.t28 92.5
R12327 VSS.n16662 VSS.n16661 92.5
R12328 VSS.n16660 VSS.n16659 92.5
R12329 VSS.n16658 VSS.n16657 92.5
R12330 VSS.n16656 VSS.n16655 92.5
R12331 VSS.n16654 VSS.n16653 92.5
R12332 VSS.n16652 VSS.n16651 92.5
R12333 VSS.n16650 VSS.n16649 92.5
R12334 VSS.n16648 VSS.n16605 92.5
R12335 VSS.t28 VSS.n16605 92.5
R12336 VSS.n16664 VSS.n16663 92.5
R12337 VSS.n16666 VSS.n16665 92.5
R12338 VSS.n16668 VSS.n16667 92.5
R12339 VSS.n16670 VSS.n16669 92.5
R12340 VSS.n16672 VSS.n16671 92.5
R12341 VSS.n16674 VSS.n16673 92.5
R12342 VSS.n16676 VSS.n16675 92.5
R12343 VSS.n16678 VSS.n16677 92.5
R12344 VSS.n16680 VSS.n16679 92.5
R12345 VSS.n16681 VSS.n16597 92.5
R12346 VSS.t28 VSS.n16597 92.5
R12347 VSS.n16685 VSS.n16684 92.5
R12348 VSS.n16760 VSS.n16616 92.5
R12349 VSS.n16751 VSS.n16613 92.5
R12350 VSS.n16695 VSS.n16617 92.5
R12351 VSS.n16699 VSS.n16612 92.5
R12352 VSS.n16703 VSS.n16618 92.5
R12353 VSS.n16707 VSS.n16611 92.5
R12354 VSS.n16766 VSS.n16621 92.5
R12355 VSS.n16713 VSS.n16615 92.5
R12356 VSS.n11114 VSS.n11113 92.5
R12357 VSS.n11063 VSS.n11061 92.5
R12358 VSS.n11102 VSS.n11101 92.5
R12359 VSS.n11104 VSS.n11103 92.5
R12360 VSS.n11106 VSS.n11105 92.5
R12361 VSS.n11108 VSS.n11107 92.5
R12362 VSS.n11110 VSS.n11109 92.5
R12363 VSS.n11112 VSS.n11111 92.5
R12364 VSS.n11235 VSS.n11234 92.5
R12365 VSS.n11234 VSS.t58 92.5
R12366 VSS.n11129 VSS.n11128 92.5
R12367 VSS.n11127 VSS.n11126 92.5
R12368 VSS.n11125 VSS.n11124 92.5
R12369 VSS.n11123 VSS.n11122 92.5
R12370 VSS.n11121 VSS.n11120 92.5
R12371 VSS.n11119 VSS.n11118 92.5
R12372 VSS.n11117 VSS.n11116 92.5
R12373 VSS.n11115 VSS.n11072 92.5
R12374 VSS.t58 VSS.n11072 92.5
R12375 VSS.n11131 VSS.n11130 92.5
R12376 VSS.n11133 VSS.n11132 92.5
R12377 VSS.n11135 VSS.n11134 92.5
R12378 VSS.n11137 VSS.n11136 92.5
R12379 VSS.n11139 VSS.n11138 92.5
R12380 VSS.n11141 VSS.n11140 92.5
R12381 VSS.n11143 VSS.n11142 92.5
R12382 VSS.n11145 VSS.n11144 92.5
R12383 VSS.n11147 VSS.n11146 92.5
R12384 VSS.n11148 VSS.n11064 92.5
R12385 VSS.t58 VSS.n11064 92.5
R12386 VSS.n11181 VSS.n11180 92.5
R12387 VSS.n11152 VSS.n11083 92.5
R12388 VSS.n11228 VSS.n11080 92.5
R12389 VSS.n11219 VSS.n11084 92.5
R12390 VSS.n11162 VSS.n11079 92.5
R12391 VSS.n11166 VSS.n11085 92.5
R12392 VSS.n11170 VSS.n11078 92.5
R12393 VSS.n11233 VSS.n11088 92.5
R12394 VSS.n11176 VSS.n11082 92.5
R12395 VSS.n11024 VSS.n11023 92.5
R12396 VSS.n10973 VSS.n10971 92.5
R12397 VSS.n11012 VSS.n11011 92.5
R12398 VSS.n11014 VSS.n11013 92.5
R12399 VSS.n11016 VSS.n11015 92.5
R12400 VSS.n11018 VSS.n11017 92.5
R12401 VSS.n11020 VSS.n11019 92.5
R12402 VSS.n11022 VSS.n11021 92.5
R12403 VSS.n11325 VSS.n11324 92.5
R12404 VSS.n11324 VSS.t32 92.5
R12405 VSS.n11039 VSS.n11038 92.5
R12406 VSS.n11037 VSS.n11036 92.5
R12407 VSS.n11035 VSS.n11034 92.5
R12408 VSS.n11033 VSS.n11032 92.5
R12409 VSS.n11031 VSS.n11030 92.5
R12410 VSS.n11029 VSS.n11028 92.5
R12411 VSS.n11027 VSS.n11026 92.5
R12412 VSS.n11025 VSS.n10982 92.5
R12413 VSS.t32 VSS.n10982 92.5
R12414 VSS.n11041 VSS.n11040 92.5
R12415 VSS.n11043 VSS.n11042 92.5
R12416 VSS.n11045 VSS.n11044 92.5
R12417 VSS.n11047 VSS.n11046 92.5
R12418 VSS.n11049 VSS.n11048 92.5
R12419 VSS.n11051 VSS.n11050 92.5
R12420 VSS.n11053 VSS.n11052 92.5
R12421 VSS.n11055 VSS.n11054 92.5
R12422 VSS.n11057 VSS.n11056 92.5
R12423 VSS.n11058 VSS.n10974 92.5
R12424 VSS.t32 VSS.n10974 92.5
R12425 VSS.n11271 VSS.n11270 92.5
R12426 VSS.n11242 VSS.n10993 92.5
R12427 VSS.n11318 VSS.n10990 92.5
R12428 VSS.n11309 VSS.n10994 92.5
R12429 VSS.n11252 VSS.n10989 92.5
R12430 VSS.n11256 VSS.n10995 92.5
R12431 VSS.n11260 VSS.n10988 92.5
R12432 VSS.n11323 VSS.n10998 92.5
R12433 VSS.n11266 VSS.n10992 92.5
R12434 VSS.n10934 VSS.n10933 92.5
R12435 VSS.n10883 VSS.n10881 92.5
R12436 VSS.n10922 VSS.n10921 92.5
R12437 VSS.n10924 VSS.n10923 92.5
R12438 VSS.n10926 VSS.n10925 92.5
R12439 VSS.n10928 VSS.n10927 92.5
R12440 VSS.n10930 VSS.n10929 92.5
R12441 VSS.n10932 VSS.n10931 92.5
R12442 VSS.n11415 VSS.n11414 92.5
R12443 VSS.n11414 VSS.t92 92.5
R12444 VSS.n10949 VSS.n10948 92.5
R12445 VSS.n10947 VSS.n10946 92.5
R12446 VSS.n10945 VSS.n10944 92.5
R12447 VSS.n10943 VSS.n10942 92.5
R12448 VSS.n10941 VSS.n10940 92.5
R12449 VSS.n10939 VSS.n10938 92.5
R12450 VSS.n10937 VSS.n10936 92.5
R12451 VSS.n10935 VSS.n10892 92.5
R12452 VSS.t92 VSS.n10892 92.5
R12453 VSS.n10951 VSS.n10950 92.5
R12454 VSS.n10953 VSS.n10952 92.5
R12455 VSS.n10955 VSS.n10954 92.5
R12456 VSS.n10957 VSS.n10956 92.5
R12457 VSS.n10959 VSS.n10958 92.5
R12458 VSS.n10961 VSS.n10960 92.5
R12459 VSS.n10963 VSS.n10962 92.5
R12460 VSS.n10965 VSS.n10964 92.5
R12461 VSS.n10967 VSS.n10966 92.5
R12462 VSS.n10968 VSS.n10884 92.5
R12463 VSS.t92 VSS.n10884 92.5
R12464 VSS.n11361 VSS.n11360 92.5
R12465 VSS.n11332 VSS.n10903 92.5
R12466 VSS.n11408 VSS.n10900 92.5
R12467 VSS.n11399 VSS.n10904 92.5
R12468 VSS.n11342 VSS.n10899 92.5
R12469 VSS.n11346 VSS.n10905 92.5
R12470 VSS.n11350 VSS.n10898 92.5
R12471 VSS.n11413 VSS.n10908 92.5
R12472 VSS.n11356 VSS.n10902 92.5
R12473 VSS.n10844 VSS.n10843 92.5
R12474 VSS.n10793 VSS.n10791 92.5
R12475 VSS.n10832 VSS.n10831 92.5
R12476 VSS.n10834 VSS.n10833 92.5
R12477 VSS.n10836 VSS.n10835 92.5
R12478 VSS.n10838 VSS.n10837 92.5
R12479 VSS.n10840 VSS.n10839 92.5
R12480 VSS.n10842 VSS.n10841 92.5
R12481 VSS.n13535 VSS.n13534 92.5
R12482 VSS.n13534 VSS.t88 92.5
R12483 VSS.n10859 VSS.n10858 92.5
R12484 VSS.n10857 VSS.n10856 92.5
R12485 VSS.n10855 VSS.n10854 92.5
R12486 VSS.n10853 VSS.n10852 92.5
R12487 VSS.n10851 VSS.n10850 92.5
R12488 VSS.n10849 VSS.n10848 92.5
R12489 VSS.n10847 VSS.n10846 92.5
R12490 VSS.n10845 VSS.n10802 92.5
R12491 VSS.t88 VSS.n10802 92.5
R12492 VSS.n10861 VSS.n10860 92.5
R12493 VSS.n10863 VSS.n10862 92.5
R12494 VSS.n10865 VSS.n10864 92.5
R12495 VSS.n10867 VSS.n10866 92.5
R12496 VSS.n10869 VSS.n10868 92.5
R12497 VSS.n10871 VSS.n10870 92.5
R12498 VSS.n10873 VSS.n10872 92.5
R12499 VSS.n10875 VSS.n10874 92.5
R12500 VSS.n10877 VSS.n10876 92.5
R12501 VSS.n10878 VSS.n10794 92.5
R12502 VSS.t88 VSS.n10794 92.5
R12503 VSS.n13480 VSS.n13479 92.5
R12504 VSS.n11422 VSS.n10813 92.5
R12505 VSS.n13528 VSS.n10810 92.5
R12506 VSS.n13519 VSS.n10814 92.5
R12507 VSS.n13461 VSS.n10809 92.5
R12508 VSS.n13465 VSS.n10815 92.5
R12509 VSS.n13469 VSS.n10808 92.5
R12510 VSS.n13533 VSS.n10818 92.5
R12511 VSS.n13475 VSS.n10812 92.5
R12512 VSS.n10754 VSS.n10753 92.5
R12513 VSS.n10703 VSS.n10701 92.5
R12514 VSS.n10742 VSS.n10741 92.5
R12515 VSS.n10744 VSS.n10743 92.5
R12516 VSS.n10746 VSS.n10745 92.5
R12517 VSS.n10748 VSS.n10747 92.5
R12518 VSS.n10750 VSS.n10749 92.5
R12519 VSS.n10752 VSS.n10751 92.5
R12520 VSS.n13625 VSS.n13624 92.5
R12521 VSS.n13624 VSS.t72 92.5
R12522 VSS.n10769 VSS.n10768 92.5
R12523 VSS.n10767 VSS.n10766 92.5
R12524 VSS.n10765 VSS.n10764 92.5
R12525 VSS.n10763 VSS.n10762 92.5
R12526 VSS.n10761 VSS.n10760 92.5
R12527 VSS.n10759 VSS.n10758 92.5
R12528 VSS.n10757 VSS.n10756 92.5
R12529 VSS.n10755 VSS.n10712 92.5
R12530 VSS.t72 VSS.n10712 92.5
R12531 VSS.n10771 VSS.n10770 92.5
R12532 VSS.n10773 VSS.n10772 92.5
R12533 VSS.n10775 VSS.n10774 92.5
R12534 VSS.n10777 VSS.n10776 92.5
R12535 VSS.n10779 VSS.n10778 92.5
R12536 VSS.n10781 VSS.n10780 92.5
R12537 VSS.n10783 VSS.n10782 92.5
R12538 VSS.n10785 VSS.n10784 92.5
R12539 VSS.n10787 VSS.n10786 92.5
R12540 VSS.n10788 VSS.n10704 92.5
R12541 VSS.t72 VSS.n10704 92.5
R12542 VSS.n13571 VSS.n13570 92.5
R12543 VSS.n13542 VSS.n10723 92.5
R12544 VSS.n13618 VSS.n10720 92.5
R12545 VSS.n13609 VSS.n10724 92.5
R12546 VSS.n13552 VSS.n10719 92.5
R12547 VSS.n13556 VSS.n10725 92.5
R12548 VSS.n13560 VSS.n10718 92.5
R12549 VSS.n13623 VSS.n10728 92.5
R12550 VSS.n13566 VSS.n10722 92.5
R12551 VSS.n10664 VSS.n10663 92.5
R12552 VSS.n10613 VSS.n10611 92.5
R12553 VSS.n10652 VSS.n10651 92.5
R12554 VSS.n10654 VSS.n10653 92.5
R12555 VSS.n10656 VSS.n10655 92.5
R12556 VSS.n10658 VSS.n10657 92.5
R12557 VSS.n10660 VSS.n10659 92.5
R12558 VSS.n10662 VSS.n10661 92.5
R12559 VSS.n13715 VSS.n13714 92.5
R12560 VSS.n13714 VSS.t78 92.5
R12561 VSS.n10679 VSS.n10678 92.5
R12562 VSS.n10677 VSS.n10676 92.5
R12563 VSS.n10675 VSS.n10674 92.5
R12564 VSS.n10673 VSS.n10672 92.5
R12565 VSS.n10671 VSS.n10670 92.5
R12566 VSS.n10669 VSS.n10668 92.5
R12567 VSS.n10667 VSS.n10666 92.5
R12568 VSS.n10665 VSS.n10622 92.5
R12569 VSS.t78 VSS.n10622 92.5
R12570 VSS.n10681 VSS.n10680 92.5
R12571 VSS.n10683 VSS.n10682 92.5
R12572 VSS.n10685 VSS.n10684 92.5
R12573 VSS.n10687 VSS.n10686 92.5
R12574 VSS.n10689 VSS.n10688 92.5
R12575 VSS.n10691 VSS.n10690 92.5
R12576 VSS.n10693 VSS.n10692 92.5
R12577 VSS.n10695 VSS.n10694 92.5
R12578 VSS.n10697 VSS.n10696 92.5
R12579 VSS.n10698 VSS.n10614 92.5
R12580 VSS.t78 VSS.n10614 92.5
R12581 VSS.n13661 VSS.n13660 92.5
R12582 VSS.n13632 VSS.n10633 92.5
R12583 VSS.n13708 VSS.n10630 92.5
R12584 VSS.n13699 VSS.n10634 92.5
R12585 VSS.n13642 VSS.n10629 92.5
R12586 VSS.n13646 VSS.n10635 92.5
R12587 VSS.n13650 VSS.n10628 92.5
R12588 VSS.n13713 VSS.n10638 92.5
R12589 VSS.n13656 VSS.n10632 92.5
R12590 VSS.n10574 VSS.n10573 92.5
R12591 VSS.n10523 VSS.n10521 92.5
R12592 VSS.n10562 VSS.n10561 92.5
R12593 VSS.n10564 VSS.n10563 92.5
R12594 VSS.n10566 VSS.n10565 92.5
R12595 VSS.n10568 VSS.n10567 92.5
R12596 VSS.n10570 VSS.n10569 92.5
R12597 VSS.n10572 VSS.n10571 92.5
R12598 VSS.n13805 VSS.n13804 92.5
R12599 VSS.n13804 VSS.t82 92.5
R12600 VSS.n10589 VSS.n10588 92.5
R12601 VSS.n10587 VSS.n10586 92.5
R12602 VSS.n10585 VSS.n10584 92.5
R12603 VSS.n10583 VSS.n10582 92.5
R12604 VSS.n10581 VSS.n10580 92.5
R12605 VSS.n10579 VSS.n10578 92.5
R12606 VSS.n10577 VSS.n10576 92.5
R12607 VSS.n10575 VSS.n10532 92.5
R12608 VSS.t82 VSS.n10532 92.5
R12609 VSS.n10591 VSS.n10590 92.5
R12610 VSS.n10593 VSS.n10592 92.5
R12611 VSS.n10595 VSS.n10594 92.5
R12612 VSS.n10597 VSS.n10596 92.5
R12613 VSS.n10599 VSS.n10598 92.5
R12614 VSS.n10601 VSS.n10600 92.5
R12615 VSS.n10603 VSS.n10602 92.5
R12616 VSS.n10605 VSS.n10604 92.5
R12617 VSS.n10607 VSS.n10606 92.5
R12618 VSS.n10608 VSS.n10524 92.5
R12619 VSS.t82 VSS.n10524 92.5
R12620 VSS.n13751 VSS.n13750 92.5
R12621 VSS.n13722 VSS.n10543 92.5
R12622 VSS.n13798 VSS.n10540 92.5
R12623 VSS.n13789 VSS.n10544 92.5
R12624 VSS.n13732 VSS.n10539 92.5
R12625 VSS.n13736 VSS.n10545 92.5
R12626 VSS.n13740 VSS.n10538 92.5
R12627 VSS.n13803 VSS.n10548 92.5
R12628 VSS.n13746 VSS.n10542 92.5
R12629 VSS.n13851 VSS.n13850 92.5
R12630 VSS.n13837 VSS.n13836 92.5
R12631 VSS.n13839 VSS.n13838 92.5
R12632 VSS.n13841 VSS.n13840 92.5
R12633 VSS.n13843 VSS.n13842 92.5
R12634 VSS.n13845 VSS.n13844 92.5
R12635 VSS.n13847 VSS.n13846 92.5
R12636 VSS.n13849 VSS.n13848 92.5
R12637 VSS.n13835 VSS.n10497 92.5
R12638 VSS.t62 VSS.n10497 92.5
R12639 VSS.n13866 VSS.n13865 92.5
R12640 VSS.n13864 VSS.n13863 92.5
R12641 VSS.n13862 VSS.n13861 92.5
R12642 VSS.n13860 VSS.n13859 92.5
R12643 VSS.n13858 VSS.n13857 92.5
R12644 VSS.n13856 VSS.n13855 92.5
R12645 VSS.n13854 VSS.n13853 92.5
R12646 VSS.n13852 VSS.n13818 92.5
R12647 VSS.t62 VSS.n13818 92.5
R12648 VSS.n13868 VSS.n13867 92.5
R12649 VSS.n13870 VSS.n13869 92.5
R12650 VSS.n13872 VSS.n13871 92.5
R12651 VSS.n13874 VSS.n13873 92.5
R12652 VSS.n13876 VSS.n13875 92.5
R12653 VSS.n13878 VSS.n13877 92.5
R12654 VSS.n13880 VSS.n13879 92.5
R12655 VSS.n13881 VSS.n13823 92.5
R12656 VSS.n13883 VSS.n13882 92.5
R12657 VSS.n13827 VSS.n13810 92.5
R12658 VSS.t62 VSS.n13810 92.5
R12659 VSS.n13954 VSS.n10494 92.5
R12660 VSS.n13885 VSS.n13809 92.5
R12661 VSS.n13894 VSS.n10503 92.5
R12662 VSS.n13948 VSS.n10505 92.5
R12663 VSS.n13939 VSS.n10502 92.5
R12664 VSS.n13904 VSS.n10506 92.5
R12665 VSS.n13908 VSS.n10501 92.5
R12666 VSS.n13912 VSS.n10507 92.5
R12667 VSS.n13913 VSS.n10500 92.5
R12668 VSS.n9132 VSS.n9131 92.5
R12669 VSS.n9146 VSS.n9145 92.5
R12670 VSS.n9144 VSS.n9143 92.5
R12671 VSS.n9142 VSS.n9141 92.5
R12672 VSS.n9140 VSS.n9139 92.5
R12673 VSS.n9138 VSS.n9137 92.5
R12674 VSS.n9136 VSS.n9135 92.5
R12675 VSS.n9134 VSS.n9133 92.5
R12676 VSS.n9147 VSS.n9016 92.5
R12677 VSS.n9116 VSS.n9115 92.5
R12678 VSS.n9118 VSS.n9117 92.5
R12679 VSS.n9120 VSS.n9119 92.5
R12680 VSS.n9122 VSS.n9121 92.5
R12681 VSS.n9124 VSS.n9123 92.5
R12682 VSS.n9126 VSS.n9125 92.5
R12683 VSS.n9128 VSS.n9127 92.5
R12684 VSS.n9130 VSS.n9129 92.5
R12685 VSS.n9114 VSS.n9113 92.5
R12686 VSS.n8984 VSS.n8982 92.5
R12687 VSS.n9099 VSS.n9098 92.5
R12688 VSS.n9101 VSS.n9100 92.5
R12689 VSS.n9103 VSS.n9102 92.5
R12690 VSS.n9105 VSS.n9104 92.5
R12691 VSS.n9107 VSS.n9106 92.5
R12692 VSS.n9109 VSS.n9108 92.5
R12693 VSS.n9111 VSS.n9110 92.5
R12694 VSS.n9112 VSS.n8993 92.5
R12695 VSS.t20 VSS.n8993 92.5
R12696 VSS.n8985 VSS.n8983 92.5
R12697 VSS.n9032 VSS.n8989 92.5
R12698 VSS.t20 VSS.n8989 92.5
R12699 VSS.n9030 VSS.n8988 92.5
R12700 VSS.t20 VSS.n8988 92.5
R12701 VSS.n9028 VSS.n8990 92.5
R12702 VSS.t20 VSS.n8990 92.5
R12703 VSS.n9026 VSS.n8987 92.5
R12704 VSS.t20 VSS.n8987 92.5
R12705 VSS.n9024 VSS.n8991 92.5
R12706 VSS.t20 VSS.n8991 92.5
R12707 VSS.n9022 VSS.n8986 92.5
R12708 VSS.t20 VSS.n8986 92.5
R12709 VSS.n9020 VSS.n8992 92.5
R12710 VSS.t20 VSS.n8992 92.5
R12711 VSS.n9017 VSS.n9015 92.5
R12712 VSS.n9242 VSS.n9241 92.5
R12713 VSS.n9191 VSS.n9189 92.5
R12714 VSS.n9230 VSS.n9229 92.5
R12715 VSS.n9232 VSS.n9231 92.5
R12716 VSS.n9234 VSS.n9233 92.5
R12717 VSS.n9236 VSS.n9235 92.5
R12718 VSS.n9238 VSS.n9237 92.5
R12719 VSS.n9240 VSS.n9239 92.5
R12720 VSS.n10263 VSS.n10262 92.5
R12721 VSS.n10262 VSS.t34 92.5
R12722 VSS.n9257 VSS.n9256 92.5
R12723 VSS.n9255 VSS.n9254 92.5
R12724 VSS.n9253 VSS.n9252 92.5
R12725 VSS.n9251 VSS.n9250 92.5
R12726 VSS.n9249 VSS.n9248 92.5
R12727 VSS.n9247 VSS.n9246 92.5
R12728 VSS.n9245 VSS.n9244 92.5
R12729 VSS.n9243 VSS.n9200 92.5
R12730 VSS.t34 VSS.n9200 92.5
R12731 VSS.n9259 VSS.n9258 92.5
R12732 VSS.n9261 VSS.n9260 92.5
R12733 VSS.n9263 VSS.n9262 92.5
R12734 VSS.n9265 VSS.n9264 92.5
R12735 VSS.n9267 VSS.n9266 92.5
R12736 VSS.n9269 VSS.n9268 92.5
R12737 VSS.n9271 VSS.n9270 92.5
R12738 VSS.n9273 VSS.n9272 92.5
R12739 VSS.n9275 VSS.n9274 92.5
R12740 VSS.n9276 VSS.n9192 92.5
R12741 VSS.t34 VSS.n9192 92.5
R12742 VSS.n10180 VSS.n10179 92.5
R12743 VSS.n10255 VSS.n9211 92.5
R12744 VSS.n10246 VSS.n9208 92.5
R12745 VSS.n10190 VSS.n9212 92.5
R12746 VSS.n10194 VSS.n9207 92.5
R12747 VSS.n10198 VSS.n9213 92.5
R12748 VSS.n10202 VSS.n9206 92.5
R12749 VSS.n10261 VSS.n9216 92.5
R12750 VSS.n10208 VSS.n9210 92.5
R12751 VSS.n9332 VSS.n9331 92.5
R12752 VSS.n9281 VSS.n9279 92.5
R12753 VSS.n9320 VSS.n9319 92.5
R12754 VSS.n9322 VSS.n9321 92.5
R12755 VSS.n9324 VSS.n9323 92.5
R12756 VSS.n9326 VSS.n9325 92.5
R12757 VSS.n9328 VSS.n9327 92.5
R12758 VSS.n9330 VSS.n9329 92.5
R12759 VSS.n10173 VSS.n10172 92.5
R12760 VSS.n10172 VSS.t26 92.5
R12761 VSS.n9347 VSS.n9346 92.5
R12762 VSS.n9345 VSS.n9344 92.5
R12763 VSS.n9343 VSS.n9342 92.5
R12764 VSS.n9341 VSS.n9340 92.5
R12765 VSS.n9339 VSS.n9338 92.5
R12766 VSS.n9337 VSS.n9336 92.5
R12767 VSS.n9335 VSS.n9334 92.5
R12768 VSS.n9333 VSS.n9290 92.5
R12769 VSS.t26 VSS.n9290 92.5
R12770 VSS.n9349 VSS.n9348 92.5
R12771 VSS.n9351 VSS.n9350 92.5
R12772 VSS.n9353 VSS.n9352 92.5
R12773 VSS.n9355 VSS.n9354 92.5
R12774 VSS.n9357 VSS.n9356 92.5
R12775 VSS.n9359 VSS.n9358 92.5
R12776 VSS.n9361 VSS.n9360 92.5
R12777 VSS.n9363 VSS.n9362 92.5
R12778 VSS.n9365 VSS.n9364 92.5
R12779 VSS.n9366 VSS.n9282 92.5
R12780 VSS.t26 VSS.n9282 92.5
R12781 VSS.n10090 VSS.n10089 92.5
R12782 VSS.n10165 VSS.n9301 92.5
R12783 VSS.n10156 VSS.n9298 92.5
R12784 VSS.n10100 VSS.n9302 92.5
R12785 VSS.n10104 VSS.n9297 92.5
R12786 VSS.n10108 VSS.n9303 92.5
R12787 VSS.n10112 VSS.n9296 92.5
R12788 VSS.n10171 VSS.n9306 92.5
R12789 VSS.n10118 VSS.n9300 92.5
R12790 VSS.n9422 VSS.n9421 92.5
R12791 VSS.n9371 VSS.n9369 92.5
R12792 VSS.n9410 VSS.n9409 92.5
R12793 VSS.n9412 VSS.n9411 92.5
R12794 VSS.n9414 VSS.n9413 92.5
R12795 VSS.n9416 VSS.n9415 92.5
R12796 VSS.n9418 VSS.n9417 92.5
R12797 VSS.n9420 VSS.n9419 92.5
R12798 VSS.n10083 VSS.n10082 92.5
R12799 VSS.n10082 VSS.t52 92.5
R12800 VSS.n9437 VSS.n9436 92.5
R12801 VSS.n9435 VSS.n9434 92.5
R12802 VSS.n9433 VSS.n9432 92.5
R12803 VSS.n9431 VSS.n9430 92.5
R12804 VSS.n9429 VSS.n9428 92.5
R12805 VSS.n9427 VSS.n9426 92.5
R12806 VSS.n9425 VSS.n9424 92.5
R12807 VSS.n9423 VSS.n9380 92.5
R12808 VSS.t52 VSS.n9380 92.5
R12809 VSS.n9439 VSS.n9438 92.5
R12810 VSS.n9441 VSS.n9440 92.5
R12811 VSS.n9443 VSS.n9442 92.5
R12812 VSS.n9445 VSS.n9444 92.5
R12813 VSS.n9447 VSS.n9446 92.5
R12814 VSS.n9449 VSS.n9448 92.5
R12815 VSS.n9451 VSS.n9450 92.5
R12816 VSS.n9453 VSS.n9452 92.5
R12817 VSS.n9455 VSS.n9454 92.5
R12818 VSS.n9456 VSS.n9372 92.5
R12819 VSS.t52 VSS.n9372 92.5
R12820 VSS.n10000 VSS.n9999 92.5
R12821 VSS.n10075 VSS.n9391 92.5
R12822 VSS.n10066 VSS.n9388 92.5
R12823 VSS.n10010 VSS.n9392 92.5
R12824 VSS.n10014 VSS.n9387 92.5
R12825 VSS.n10018 VSS.n9393 92.5
R12826 VSS.n10022 VSS.n9386 92.5
R12827 VSS.n10081 VSS.n9396 92.5
R12828 VSS.n10028 VSS.n9390 92.5
R12829 VSS.n9512 VSS.n9511 92.5
R12830 VSS.n9461 VSS.n9459 92.5
R12831 VSS.n9500 VSS.n9499 92.5
R12832 VSS.n9502 VSS.n9501 92.5
R12833 VSS.n9504 VSS.n9503 92.5
R12834 VSS.n9506 VSS.n9505 92.5
R12835 VSS.n9508 VSS.n9507 92.5
R12836 VSS.n9510 VSS.n9509 92.5
R12837 VSS.n9993 VSS.n9992 92.5
R12838 VSS.n9992 VSS.t56 92.5
R12839 VSS.n9527 VSS.n9526 92.5
R12840 VSS.n9525 VSS.n9524 92.5
R12841 VSS.n9523 VSS.n9522 92.5
R12842 VSS.n9521 VSS.n9520 92.5
R12843 VSS.n9519 VSS.n9518 92.5
R12844 VSS.n9517 VSS.n9516 92.5
R12845 VSS.n9515 VSS.n9514 92.5
R12846 VSS.n9513 VSS.n9470 92.5
R12847 VSS.t56 VSS.n9470 92.5
R12848 VSS.n9529 VSS.n9528 92.5
R12849 VSS.n9531 VSS.n9530 92.5
R12850 VSS.n9533 VSS.n9532 92.5
R12851 VSS.n9535 VSS.n9534 92.5
R12852 VSS.n9537 VSS.n9536 92.5
R12853 VSS.n9539 VSS.n9538 92.5
R12854 VSS.n9541 VSS.n9540 92.5
R12855 VSS.n9543 VSS.n9542 92.5
R12856 VSS.n9545 VSS.n9544 92.5
R12857 VSS.n9546 VSS.n9462 92.5
R12858 VSS.t56 VSS.n9462 92.5
R12859 VSS.n9910 VSS.n9909 92.5
R12860 VSS.n9985 VSS.n9481 92.5
R12861 VSS.n9976 VSS.n9478 92.5
R12862 VSS.n9920 VSS.n9482 92.5
R12863 VSS.n9924 VSS.n9477 92.5
R12864 VSS.n9928 VSS.n9483 92.5
R12865 VSS.n9932 VSS.n9476 92.5
R12866 VSS.n9991 VSS.n9486 92.5
R12867 VSS.n9938 VSS.n9480 92.5
R12868 VSS.n9602 VSS.n9601 92.5
R12869 VSS.n9551 VSS.n9549 92.5
R12870 VSS.n9590 VSS.n9589 92.5
R12871 VSS.n9592 VSS.n9591 92.5
R12872 VSS.n9594 VSS.n9593 92.5
R12873 VSS.n9596 VSS.n9595 92.5
R12874 VSS.n9598 VSS.n9597 92.5
R12875 VSS.n9600 VSS.n9599 92.5
R12876 VSS.n9903 VSS.n9902 92.5
R12877 VSS.n9902 VSS.t80 92.5
R12878 VSS.n9617 VSS.n9616 92.5
R12879 VSS.n9615 VSS.n9614 92.5
R12880 VSS.n9613 VSS.n9612 92.5
R12881 VSS.n9611 VSS.n9610 92.5
R12882 VSS.n9609 VSS.n9608 92.5
R12883 VSS.n9607 VSS.n9606 92.5
R12884 VSS.n9605 VSS.n9604 92.5
R12885 VSS.n9603 VSS.n9560 92.5
R12886 VSS.t80 VSS.n9560 92.5
R12887 VSS.n9619 VSS.n9618 92.5
R12888 VSS.n9621 VSS.n9620 92.5
R12889 VSS.n9623 VSS.n9622 92.5
R12890 VSS.n9625 VSS.n9624 92.5
R12891 VSS.n9627 VSS.n9626 92.5
R12892 VSS.n9629 VSS.n9628 92.5
R12893 VSS.n9631 VSS.n9630 92.5
R12894 VSS.n9633 VSS.n9632 92.5
R12895 VSS.n9635 VSS.n9634 92.5
R12896 VSS.n9636 VSS.n9552 92.5
R12897 VSS.t80 VSS.n9552 92.5
R12898 VSS.n9820 VSS.n9819 92.5
R12899 VSS.n9895 VSS.n9571 92.5
R12900 VSS.n9886 VSS.n9568 92.5
R12901 VSS.n9830 VSS.n9572 92.5
R12902 VSS.n9834 VSS.n9567 92.5
R12903 VSS.n9838 VSS.n9573 92.5
R12904 VSS.n9842 VSS.n9566 92.5
R12905 VSS.n9901 VSS.n9576 92.5
R12906 VSS.n9848 VSS.n9570 92.5
R12907 VSS.n9692 VSS.n9691 92.5
R12908 VSS.n9641 VSS.n9639 92.5
R12909 VSS.n9680 VSS.n9679 92.5
R12910 VSS.n9682 VSS.n9681 92.5
R12911 VSS.n9684 VSS.n9683 92.5
R12912 VSS.n9686 VSS.n9685 92.5
R12913 VSS.n9688 VSS.n9687 92.5
R12914 VSS.n9690 VSS.n9689 92.5
R12915 VSS.n9813 VSS.n9812 92.5
R12916 VSS.n9812 VSS.t18 92.5
R12917 VSS.n9707 VSS.n9706 92.5
R12918 VSS.n9705 VSS.n9704 92.5
R12919 VSS.n9703 VSS.n9702 92.5
R12920 VSS.n9701 VSS.n9700 92.5
R12921 VSS.n9699 VSS.n9698 92.5
R12922 VSS.n9697 VSS.n9696 92.5
R12923 VSS.n9695 VSS.n9694 92.5
R12924 VSS.n9693 VSS.n9650 92.5
R12925 VSS.t18 VSS.n9650 92.5
R12926 VSS.n9709 VSS.n9708 92.5
R12927 VSS.n9711 VSS.n9710 92.5
R12928 VSS.n9713 VSS.n9712 92.5
R12929 VSS.n9715 VSS.n9714 92.5
R12930 VSS.n9717 VSS.n9716 92.5
R12931 VSS.n9719 VSS.n9718 92.5
R12932 VSS.n9721 VSS.n9720 92.5
R12933 VSS.n9723 VSS.n9722 92.5
R12934 VSS.n9725 VSS.n9724 92.5
R12935 VSS.n9726 VSS.n9642 92.5
R12936 VSS.t18 VSS.n9642 92.5
R12937 VSS.n9730 VSS.n9729 92.5
R12938 VSS.n9805 VSS.n9661 92.5
R12939 VSS.n9796 VSS.n9658 92.5
R12940 VSS.n9740 VSS.n9662 92.5
R12941 VSS.n9744 VSS.n9657 92.5
R12942 VSS.n9748 VSS.n9663 92.5
R12943 VSS.n9752 VSS.n9656 92.5
R12944 VSS.n9811 VSS.n9666 92.5
R12945 VSS.n9758 VSS.n9660 92.5
R12946 VSS.n10280 VSS.n10279 92.5
R12947 VSS.n10266 VSS.n9164 92.5
R12948 VSS.n10268 VSS.n10267 92.5
R12949 VSS.n10270 VSS.n10269 92.5
R12950 VSS.n10272 VSS.n10271 92.5
R12951 VSS.n10274 VSS.n10273 92.5
R12952 VSS.n10276 VSS.n10275 92.5
R12953 VSS.n10278 VSS.n10277 92.5
R12954 VSS.n10325 VSS.n9163 92.5
R12955 VSS.n10296 VSS.n10295 92.5
R12956 VSS.n10294 VSS.n10293 92.5
R12957 VSS.n10292 VSS.n10291 92.5
R12958 VSS.n10290 VSS.n10289 92.5
R12959 VSS.n10288 VSS.n10287 92.5
R12960 VSS.n10286 VSS.n10285 92.5
R12961 VSS.n10284 VSS.n10283 92.5
R12962 VSS.n10282 VSS.n10281 92.5
R12963 VSS.n10298 VSS.n10297 92.5
R12964 VSS.n10316 VSS.n10315 92.5
R12965 VSS.n10313 VSS.n10312 92.5
R12966 VSS.n10311 VSS.n10310 92.5
R12967 VSS.n10309 VSS.n10308 92.5
R12968 VSS.n10307 VSS.n10306 92.5
R12969 VSS.n10305 VSS.n10304 92.5
R12970 VSS.n10303 VSS.n10302 92.5
R12971 VSS.n10301 VSS.n10300 92.5
R12972 VSS.n10299 VSS.n9165 92.5
R12973 VSS.t38 VSS.n9165 92.5
R12974 VSS.n8934 VSS.n8932 92.5
R12975 VSS.n10364 VSS.n8936 92.5
R12976 VSS.n10358 VSS.n8941 92.5
R12977 VSS.n10352 VSS.n8947 92.5
R12978 VSS.n10346 VSS.n8953 92.5
R12979 VSS.n10340 VSS.n8958 92.5
R12980 VSS.n10334 VSS.n8965 92.5
R12981 VSS.n10328 VSS.n8971 92.5
R12982 VSS.n10323 VSS.n10322 92.5
R12983 VSS.n6691 VSS.n6659 92.5
R12984 VSS.n6678 VSS.n6677 92.5
R12985 VSS.n6680 VSS.n6679 92.5
R12986 VSS.n6682 VSS.n6681 92.5
R12987 VSS.n6684 VSS.n6683 92.5
R12988 VSS.n6686 VSS.n6685 92.5
R12989 VSS.n6688 VSS.n6687 92.5
R12990 VSS.n6690 VSS.n6689 92.5
R12991 VSS.n6676 VSS.n6675 92.5
R12992 VSS.n6693 VSS.n6692 92.5
R12993 VSS.n6695 VSS.n6694 92.5
R12994 VSS.n6697 VSS.n6696 92.5
R12995 VSS.n6699 VSS.n6698 92.5
R12996 VSS.n6701 VSS.n6700 92.5
R12997 VSS.n6703 VSS.n6702 92.5
R12998 VSS.n6705 VSS.n6704 92.5
R12999 VSS.n6707 VSS.n6706 92.5
R13000 VSS.n6709 VSS.n6708 92.5
R13001 VSS.n6711 VSS.n6710 92.5
R13002 VSS.n6713 VSS.n6712 92.5
R13003 VSS.n6715 VSS.n6714 92.5
R13004 VSS.n6717 VSS.n6716 92.5
R13005 VSS.n6719 VSS.n6718 92.5
R13006 VSS.n6720 VSS.n6658 92.5
R13007 VSS.n6723 VSS.n6722 92.5
R13008 VSS.n6721 VSS.n6638 92.5
R13009 VSS.n6725 VSS.n6635 92.5
R13010 VSS.n6725 VSS.t14 92.5
R13011 VSS.n6674 VSS.n6673 92.5
R13012 VSS.n6672 VSS.n6671 92.5
R13013 VSS.n6670 VSS.n6669 92.5
R13014 VSS.n6668 VSS.n6667 92.5
R13015 VSS.n6666 VSS.n6665 92.5
R13016 VSS.n6664 VSS.n6663 92.5
R13017 VSS.n6662 VSS.n6661 92.5
R13018 VSS.n6660 VSS.n6636 92.5
R13019 VSS.n6727 VSS.n6726 92.5
R13020 VSS.n5699 VSS.n5698 92.5
R13021 VSS.n5685 VSS.n3631 92.5
R13022 VSS.n5687 VSS.n5686 92.5
R13023 VSS.n5689 VSS.n5688 92.5
R13024 VSS.n5691 VSS.n5690 92.5
R13025 VSS.n5693 VSS.n5692 92.5
R13026 VSS.n5695 VSS.n5694 92.5
R13027 VSS.n5697 VSS.n5696 92.5
R13028 VSS.n5734 VSS.n5667 92.5
R13029 VSS.n5734 VSS.t46 92.5
R13030 VSS.n5714 VSS.n5713 92.5
R13031 VSS.n5712 VSS.n5711 92.5
R13032 VSS.n5710 VSS.n5709 92.5
R13033 VSS.n5708 VSS.n5707 92.5
R13034 VSS.n5706 VSS.n5705 92.5
R13035 VSS.n5704 VSS.n5703 92.5
R13036 VSS.n5702 VSS.n5701 92.5
R13037 VSS.n5700 VSS.n5678 92.5
R13038 VSS.t46 VSS.n5678 92.5
R13039 VSS.n5716 VSS.n5715 92.5
R13040 VSS.n5718 VSS.n5717 92.5
R13041 VSS.n5720 VSS.n5719 92.5
R13042 VSS.n5722 VSS.n5721 92.5
R13043 VSS.n5724 VSS.n5723 92.5
R13044 VSS.n5726 VSS.n5725 92.5
R13045 VSS.n5728 VSS.n5727 92.5
R13046 VSS.n5729 VSS.n5683 92.5
R13047 VSS.n5731 VSS.n5730 92.5
R13048 VSS.n5684 VSS.n5670 92.5
R13049 VSS.t46 VSS.n5670 92.5
R13050 VSS.n3581 VSS.n3579 92.5
R13051 VSS.n5779 VSS.n3583 92.5
R13052 VSS.n5773 VSS.n3588 92.5
R13053 VSS.n5767 VSS.n3594 92.5
R13054 VSS.n5761 VSS.n3600 92.5
R13055 VSS.n5755 VSS.n3606 92.5
R13056 VSS.n5749 VSS.n3611 92.5
R13057 VSS.n5743 VSS.n3618 92.5
R13058 VSS.n5737 VSS.n3624 92.5
R13059 VSS.n5821 VSS.n5820 92.5
R13060 VSS.n5807 VSS.n3573 92.5
R13061 VSS.n5809 VSS.n5808 92.5
R13062 VSS.n5811 VSS.n5810 92.5
R13063 VSS.n5813 VSS.n5812 92.5
R13064 VSS.n5815 VSS.n5814 92.5
R13065 VSS.n5817 VSS.n5816 92.5
R13066 VSS.n5819 VSS.n5818 92.5
R13067 VSS.n5856 VSS.n5789 92.5
R13068 VSS.n5856 VSS.t70 92.5
R13069 VSS.n5836 VSS.n5835 92.5
R13070 VSS.n5834 VSS.n5833 92.5
R13071 VSS.n5832 VSS.n5831 92.5
R13072 VSS.n5830 VSS.n5829 92.5
R13073 VSS.n5828 VSS.n5827 92.5
R13074 VSS.n5826 VSS.n5825 92.5
R13075 VSS.n5824 VSS.n5823 92.5
R13076 VSS.n5822 VSS.n5800 92.5
R13077 VSS.t70 VSS.n5800 92.5
R13078 VSS.n5838 VSS.n5837 92.5
R13079 VSS.n5840 VSS.n5839 92.5
R13080 VSS.n5842 VSS.n5841 92.5
R13081 VSS.n5844 VSS.n5843 92.5
R13082 VSS.n5846 VSS.n5845 92.5
R13083 VSS.n5848 VSS.n5847 92.5
R13084 VSS.n5850 VSS.n5849 92.5
R13085 VSS.n5851 VSS.n5805 92.5
R13086 VSS.n5853 VSS.n5852 92.5
R13087 VSS.n5806 VSS.n5792 92.5
R13088 VSS.t70 VSS.n5792 92.5
R13089 VSS.n3523 VSS.n3521 92.5
R13090 VSS.n5901 VSS.n3525 92.5
R13091 VSS.n5895 VSS.n3530 92.5
R13092 VSS.n5889 VSS.n3536 92.5
R13093 VSS.n5883 VSS.n3542 92.5
R13094 VSS.n5877 VSS.n3548 92.5
R13095 VSS.n5871 VSS.n3553 92.5
R13096 VSS.n5865 VSS.n3560 92.5
R13097 VSS.n5859 VSS.n3566 92.5
R13098 VSS.n5943 VSS.n5942 92.5
R13099 VSS.n5929 VSS.n3515 92.5
R13100 VSS.n5931 VSS.n5930 92.5
R13101 VSS.n5933 VSS.n5932 92.5
R13102 VSS.n5935 VSS.n5934 92.5
R13103 VSS.n5937 VSS.n5936 92.5
R13104 VSS.n5939 VSS.n5938 92.5
R13105 VSS.n5941 VSS.n5940 92.5
R13106 VSS.n5978 VSS.n5911 92.5
R13107 VSS.n5978 VSS.t66 92.5
R13108 VSS.n5958 VSS.n5957 92.5
R13109 VSS.n5956 VSS.n5955 92.5
R13110 VSS.n5954 VSS.n5953 92.5
R13111 VSS.n5952 VSS.n5951 92.5
R13112 VSS.n5950 VSS.n5949 92.5
R13113 VSS.n5948 VSS.n5947 92.5
R13114 VSS.n5946 VSS.n5945 92.5
R13115 VSS.n5944 VSS.n5922 92.5
R13116 VSS.t66 VSS.n5922 92.5
R13117 VSS.n5960 VSS.n5959 92.5
R13118 VSS.n5962 VSS.n5961 92.5
R13119 VSS.n5964 VSS.n5963 92.5
R13120 VSS.n5966 VSS.n5965 92.5
R13121 VSS.n5968 VSS.n5967 92.5
R13122 VSS.n5970 VSS.n5969 92.5
R13123 VSS.n5972 VSS.n5971 92.5
R13124 VSS.n5973 VSS.n5927 92.5
R13125 VSS.n5975 VSS.n5974 92.5
R13126 VSS.n5928 VSS.n5914 92.5
R13127 VSS.t66 VSS.n5914 92.5
R13128 VSS.n3465 VSS.n3463 92.5
R13129 VSS.n6023 VSS.n3467 92.5
R13130 VSS.n6017 VSS.n3472 92.5
R13131 VSS.n6011 VSS.n3478 92.5
R13132 VSS.n6005 VSS.n3484 92.5
R13133 VSS.n5999 VSS.n3490 92.5
R13134 VSS.n5993 VSS.n3495 92.5
R13135 VSS.n5987 VSS.n3502 92.5
R13136 VSS.n5981 VSS.n3508 92.5
R13137 VSS.n6065 VSS.n6064 92.5
R13138 VSS.n6051 VSS.n3457 92.5
R13139 VSS.n6053 VSS.n6052 92.5
R13140 VSS.n6055 VSS.n6054 92.5
R13141 VSS.n6057 VSS.n6056 92.5
R13142 VSS.n6059 VSS.n6058 92.5
R13143 VSS.n6061 VSS.n6060 92.5
R13144 VSS.n6063 VSS.n6062 92.5
R13145 VSS.n6100 VSS.n6033 92.5
R13146 VSS.n6100 VSS.t64 92.5
R13147 VSS.n6080 VSS.n6079 92.5
R13148 VSS.n6078 VSS.n6077 92.5
R13149 VSS.n6076 VSS.n6075 92.5
R13150 VSS.n6074 VSS.n6073 92.5
R13151 VSS.n6072 VSS.n6071 92.5
R13152 VSS.n6070 VSS.n6069 92.5
R13153 VSS.n6068 VSS.n6067 92.5
R13154 VSS.n6066 VSS.n6044 92.5
R13155 VSS.t64 VSS.n6044 92.5
R13156 VSS.n6082 VSS.n6081 92.5
R13157 VSS.n6084 VSS.n6083 92.5
R13158 VSS.n6086 VSS.n6085 92.5
R13159 VSS.n6088 VSS.n6087 92.5
R13160 VSS.n6090 VSS.n6089 92.5
R13161 VSS.n6092 VSS.n6091 92.5
R13162 VSS.n6094 VSS.n6093 92.5
R13163 VSS.n6095 VSS.n6049 92.5
R13164 VSS.n6097 VSS.n6096 92.5
R13165 VSS.n6050 VSS.n6036 92.5
R13166 VSS.t64 VSS.n6036 92.5
R13167 VSS.n3407 VSS.n3405 92.5
R13168 VSS.n6145 VSS.n3409 92.5
R13169 VSS.n6139 VSS.n3414 92.5
R13170 VSS.n6133 VSS.n3420 92.5
R13171 VSS.n6127 VSS.n3426 92.5
R13172 VSS.n6121 VSS.n3432 92.5
R13173 VSS.n6115 VSS.n3437 92.5
R13174 VSS.n6109 VSS.n3444 92.5
R13175 VSS.n6103 VSS.n3450 92.5
R13176 VSS.n6187 VSS.n6186 92.5
R13177 VSS.n6173 VSS.n3399 92.5
R13178 VSS.n6175 VSS.n6174 92.5
R13179 VSS.n6177 VSS.n6176 92.5
R13180 VSS.n6179 VSS.n6178 92.5
R13181 VSS.n6181 VSS.n6180 92.5
R13182 VSS.n6183 VSS.n6182 92.5
R13183 VSS.n6185 VSS.n6184 92.5
R13184 VSS.n6222 VSS.n6155 92.5
R13185 VSS.n6222 VSS.t84 92.5
R13186 VSS.n6202 VSS.n6201 92.5
R13187 VSS.n6200 VSS.n6199 92.5
R13188 VSS.n6198 VSS.n6197 92.5
R13189 VSS.n6196 VSS.n6195 92.5
R13190 VSS.n6194 VSS.n6193 92.5
R13191 VSS.n6192 VSS.n6191 92.5
R13192 VSS.n6190 VSS.n6189 92.5
R13193 VSS.n6188 VSS.n6166 92.5
R13194 VSS.t84 VSS.n6166 92.5
R13195 VSS.n6204 VSS.n6203 92.5
R13196 VSS.n6206 VSS.n6205 92.5
R13197 VSS.n6208 VSS.n6207 92.5
R13198 VSS.n6210 VSS.n6209 92.5
R13199 VSS.n6212 VSS.n6211 92.5
R13200 VSS.n6214 VSS.n6213 92.5
R13201 VSS.n6216 VSS.n6215 92.5
R13202 VSS.n6217 VSS.n6171 92.5
R13203 VSS.n6219 VSS.n6218 92.5
R13204 VSS.n6172 VSS.n6158 92.5
R13205 VSS.t84 VSS.n6158 92.5
R13206 VSS.n3349 VSS.n3347 92.5
R13207 VSS.n6267 VSS.n3351 92.5
R13208 VSS.n6261 VSS.n3356 92.5
R13209 VSS.n6255 VSS.n3362 92.5
R13210 VSS.n6249 VSS.n3368 92.5
R13211 VSS.n6243 VSS.n3374 92.5
R13212 VSS.n6237 VSS.n3379 92.5
R13213 VSS.n6231 VSS.n3386 92.5
R13214 VSS.n6225 VSS.n3392 92.5
R13215 VSS.n6309 VSS.n6308 92.5
R13216 VSS.n6295 VSS.n3341 92.5
R13217 VSS.n6297 VSS.n6296 92.5
R13218 VSS.n6299 VSS.n6298 92.5
R13219 VSS.n6301 VSS.n6300 92.5
R13220 VSS.n6303 VSS.n6302 92.5
R13221 VSS.n6305 VSS.n6304 92.5
R13222 VSS.n6307 VSS.n6306 92.5
R13223 VSS.n6344 VSS.n6277 92.5
R13224 VSS.n6344 VSS.t86 92.5
R13225 VSS.n6324 VSS.n6323 92.5
R13226 VSS.n6322 VSS.n6321 92.5
R13227 VSS.n6320 VSS.n6319 92.5
R13228 VSS.n6318 VSS.n6317 92.5
R13229 VSS.n6316 VSS.n6315 92.5
R13230 VSS.n6314 VSS.n6313 92.5
R13231 VSS.n6312 VSS.n6311 92.5
R13232 VSS.n6310 VSS.n6288 92.5
R13233 VSS.t86 VSS.n6288 92.5
R13234 VSS.n6326 VSS.n6325 92.5
R13235 VSS.n6328 VSS.n6327 92.5
R13236 VSS.n6330 VSS.n6329 92.5
R13237 VSS.n6332 VSS.n6331 92.5
R13238 VSS.n6334 VSS.n6333 92.5
R13239 VSS.n6336 VSS.n6335 92.5
R13240 VSS.n6338 VSS.n6337 92.5
R13241 VSS.n6339 VSS.n6293 92.5
R13242 VSS.n6341 VSS.n6340 92.5
R13243 VSS.n6294 VSS.n6280 92.5
R13244 VSS.t86 VSS.n6280 92.5
R13245 VSS.n3291 VSS.n3289 92.5
R13246 VSS.n6389 VSS.n3293 92.5
R13247 VSS.n6383 VSS.n3298 92.5
R13248 VSS.n6377 VSS.n3304 92.5
R13249 VSS.n6371 VSS.n3310 92.5
R13250 VSS.n6365 VSS.n3316 92.5
R13251 VSS.n6359 VSS.n3321 92.5
R13252 VSS.n6353 VSS.n3328 92.5
R13253 VSS.n6347 VSS.n3334 92.5
R13254 VSS.n6431 VSS.n6430 92.5
R13255 VSS.n6417 VSS.n3283 92.5
R13256 VSS.n6419 VSS.n6418 92.5
R13257 VSS.n6421 VSS.n6420 92.5
R13258 VSS.n6423 VSS.n6422 92.5
R13259 VSS.n6425 VSS.n6424 92.5
R13260 VSS.n6427 VSS.n6426 92.5
R13261 VSS.n6429 VSS.n6428 92.5
R13262 VSS.n6466 VSS.n6399 92.5
R13263 VSS.n6466 VSS.t24 92.5
R13264 VSS.n6446 VSS.n6445 92.5
R13265 VSS.n6444 VSS.n6443 92.5
R13266 VSS.n6442 VSS.n6441 92.5
R13267 VSS.n6440 VSS.n6439 92.5
R13268 VSS.n6438 VSS.n6437 92.5
R13269 VSS.n6436 VSS.n6435 92.5
R13270 VSS.n6434 VSS.n6433 92.5
R13271 VSS.n6432 VSS.n6410 92.5
R13272 VSS.t24 VSS.n6410 92.5
R13273 VSS.n6448 VSS.n6447 92.5
R13274 VSS.n6450 VSS.n6449 92.5
R13275 VSS.n6452 VSS.n6451 92.5
R13276 VSS.n6454 VSS.n6453 92.5
R13277 VSS.n6456 VSS.n6455 92.5
R13278 VSS.n6458 VSS.n6457 92.5
R13279 VSS.n6460 VSS.n6459 92.5
R13280 VSS.n6461 VSS.n6415 92.5
R13281 VSS.n6463 VSS.n6462 92.5
R13282 VSS.n6416 VSS.n6402 92.5
R13283 VSS.t24 VSS.n6402 92.5
R13284 VSS.n3233 VSS.n3231 92.5
R13285 VSS.n6511 VSS.n3235 92.5
R13286 VSS.n6505 VSS.n3240 92.5
R13287 VSS.n6499 VSS.n3246 92.5
R13288 VSS.n6493 VSS.n3252 92.5
R13289 VSS.n6487 VSS.n3258 92.5
R13290 VSS.n6481 VSS.n3263 92.5
R13291 VSS.n6475 VSS.n3270 92.5
R13292 VSS.n6469 VSS.n3276 92.5
R13293 VSS.n6575 VSS.n6525 92.5
R13294 VSS.n6588 VSS.n6587 92.5
R13295 VSS.n6585 VSS.n6520 92.5
R13296 VSS.n6584 VSS.n6583 92.5
R13297 VSS.n6582 VSS.n6581 92.5
R13298 VSS.n6580 VSS.n6522 92.5
R13299 VSS.n6578 VSS.n6577 92.5
R13300 VSS.n6576 VSS.n6523 92.5
R13301 VSS.n6589 VSS.n3158 92.5
R13302 VSS.n3158 VSS.t44 92.5
R13303 VSS.n6560 VSS.n6529 92.5
R13304 VSS.n6562 VSS.n6561 92.5
R13305 VSS.n6564 VSS.n6528 92.5
R13306 VSS.n6567 VSS.n6566 92.5
R13307 VSS.n6568 VSS.n6527 92.5
R13308 VSS.n6570 VSS.n6569 92.5
R13309 VSS.n6572 VSS.n6526 92.5
R13310 VSS.n6574 VSS.n6573 92.5
R13311 VSS.n6573 VSS.t44 92.5
R13312 VSS.n6559 VSS.n6558 92.5
R13313 VSS.n6556 VSS.n6530 92.5
R13314 VSS.n6554 VSS.n6553 92.5
R13315 VSS.n6552 VSS.n6531 92.5
R13316 VSS.n6551 VSS.n6550 92.5
R13317 VSS.n6548 VSS.n6532 92.5
R13318 VSS.n6546 VSS.n6545 92.5
R13319 VSS.n6544 VSS.n6533 92.5
R13320 VSS.n6543 VSS.n6542 92.5
R13321 VSS.n6540 VSS.n6539 92.5
R13322 VSS.n6540 VSS.t44 92.5
R13323 VSS.n6536 VSS.n6535 92.5
R13324 VSS.n6599 VSS.n3139 92.5
R13325 VSS.n3172 VSS.n3144 92.5
R13326 VSS.n3170 VSS.n3146 92.5
R13327 VSS.n3168 VSS.n3143 92.5
R13328 VSS.n3166 VSS.n3147 92.5
R13329 VSS.n3164 VSS.n3142 92.5
R13330 VSS.n3162 VSS.n3148 92.5
R13331 VSS.n3159 VSS.n3157 92.5
R13332 VSS.n60 VSS.n59 92.5
R13333 VSS.n46 VSS.n8 92.5
R13334 VSS.n48 VSS.n47 92.5
R13335 VSS.n50 VSS.n49 92.5
R13336 VSS.n52 VSS.n51 92.5
R13337 VSS.n54 VSS.n53 92.5
R13338 VSS.n56 VSS.n55 92.5
R13339 VSS.n58 VSS.n57 92.5
R13340 VSS.n1254 VSS.n3 92.5
R13341 VSS.n1254 VSS.t60 92.5
R13342 VSS.n75 VSS.n74 92.5
R13343 VSS.n73 VSS.n72 92.5
R13344 VSS.n71 VSS.n70 92.5
R13345 VSS.n69 VSS.n68 92.5
R13346 VSS.n67 VSS.n66 92.5
R13347 VSS.n65 VSS.n64 92.5
R13348 VSS.n63 VSS.n62 92.5
R13349 VSS.n61 VSS.n17 92.5
R13350 VSS.t60 VSS.n17 92.5
R13351 VSS.n77 VSS.n76 92.5
R13352 VSS.n79 VSS.n78 92.5
R13353 VSS.n81 VSS.n80 92.5
R13354 VSS.n83 VSS.n82 92.5
R13355 VSS.n85 VSS.n84 92.5
R13356 VSS.n87 VSS.n86 92.5
R13357 VSS.n89 VSS.n88 92.5
R13358 VSS.n91 VSS.n90 92.5
R13359 VSS.n93 VSS.n92 92.5
R13360 VSS.n94 VSS.n9 92.5
R13361 VSS.t60 VSS.n9 92.5
R13362 VSS.n1178 VSS.n1177 92.5
R13363 VSS.n1248 VSS.n28 92.5
R13364 VSS.n1239 VSS.n25 92.5
R13365 VSS.n1188 VSS.n29 92.5
R13366 VSS.n1192 VSS.n24 92.5
R13367 VSS.n1196 VSS.n30 92.5
R13368 VSS.n1200 VSS.n23 92.5
R13369 VSS.n1253 VSS.n33 92.5
R13370 VSS.n27 VSS.n6 92.5
R13371 VSS.n150 VSS.n149 92.5
R13372 VSS.n99 VSS.n97 92.5
R13373 VSS.n138 VSS.n137 92.5
R13374 VSS.n140 VSS.n139 92.5
R13375 VSS.n142 VSS.n141 92.5
R13376 VSS.n144 VSS.n143 92.5
R13377 VSS.n146 VSS.n145 92.5
R13378 VSS.n148 VSS.n147 92.5
R13379 VSS.n1171 VSS.n1170 92.5
R13380 VSS.n1170 VSS.t48 92.5
R13381 VSS.n165 VSS.n164 92.5
R13382 VSS.n163 VSS.n162 92.5
R13383 VSS.n161 VSS.n160 92.5
R13384 VSS.n159 VSS.n158 92.5
R13385 VSS.n157 VSS.n156 92.5
R13386 VSS.n155 VSS.n154 92.5
R13387 VSS.n153 VSS.n152 92.5
R13388 VSS.n151 VSS.n108 92.5
R13389 VSS.t48 VSS.n108 92.5
R13390 VSS.n167 VSS.n166 92.5
R13391 VSS.n169 VSS.n168 92.5
R13392 VSS.n171 VSS.n170 92.5
R13393 VSS.n173 VSS.n172 92.5
R13394 VSS.n175 VSS.n174 92.5
R13395 VSS.n177 VSS.n176 92.5
R13396 VSS.n179 VSS.n178 92.5
R13397 VSS.n181 VSS.n180 92.5
R13398 VSS.n183 VSS.n182 92.5
R13399 VSS.n184 VSS.n100 92.5
R13400 VSS.t48 VSS.n100 92.5
R13401 VSS.n1088 VSS.n1087 92.5
R13402 VSS.n1163 VSS.n119 92.5
R13403 VSS.n1154 VSS.n116 92.5
R13404 VSS.n1098 VSS.n120 92.5
R13405 VSS.n1102 VSS.n115 92.5
R13406 VSS.n1106 VSS.n121 92.5
R13407 VSS.n1110 VSS.n114 92.5
R13408 VSS.n1169 VSS.n124 92.5
R13409 VSS.n1116 VSS.n118 92.5
R13410 VSS.n240 VSS.n239 92.5
R13411 VSS.n189 VSS.n187 92.5
R13412 VSS.n228 VSS.n227 92.5
R13413 VSS.n230 VSS.n229 92.5
R13414 VSS.n232 VSS.n231 92.5
R13415 VSS.n234 VSS.n233 92.5
R13416 VSS.n236 VSS.n235 92.5
R13417 VSS.n238 VSS.n237 92.5
R13418 VSS.n1081 VSS.n1080 92.5
R13419 VSS.n1080 VSS.t76 92.5
R13420 VSS.n255 VSS.n254 92.5
R13421 VSS.n253 VSS.n252 92.5
R13422 VSS.n251 VSS.n250 92.5
R13423 VSS.n249 VSS.n248 92.5
R13424 VSS.n247 VSS.n246 92.5
R13425 VSS.n245 VSS.n244 92.5
R13426 VSS.n243 VSS.n242 92.5
R13427 VSS.n241 VSS.n198 92.5
R13428 VSS.t76 VSS.n198 92.5
R13429 VSS.n257 VSS.n256 92.5
R13430 VSS.n259 VSS.n258 92.5
R13431 VSS.n261 VSS.n260 92.5
R13432 VSS.n263 VSS.n262 92.5
R13433 VSS.n265 VSS.n264 92.5
R13434 VSS.n267 VSS.n266 92.5
R13435 VSS.n269 VSS.n268 92.5
R13436 VSS.n271 VSS.n270 92.5
R13437 VSS.n273 VSS.n272 92.5
R13438 VSS.n274 VSS.n190 92.5
R13439 VSS.t76 VSS.n190 92.5
R13440 VSS.n998 VSS.n997 92.5
R13441 VSS.n1073 VSS.n209 92.5
R13442 VSS.n1064 VSS.n206 92.5
R13443 VSS.n1008 VSS.n210 92.5
R13444 VSS.n1012 VSS.n205 92.5
R13445 VSS.n1016 VSS.n211 92.5
R13446 VSS.n1020 VSS.n204 92.5
R13447 VSS.n1079 VSS.n214 92.5
R13448 VSS.n1026 VSS.n208 92.5
R13449 VSS.n330 VSS.n329 92.5
R13450 VSS.n279 VSS.n277 92.5
R13451 VSS.n318 VSS.n317 92.5
R13452 VSS.n320 VSS.n319 92.5
R13453 VSS.n322 VSS.n321 92.5
R13454 VSS.n324 VSS.n323 92.5
R13455 VSS.n326 VSS.n325 92.5
R13456 VSS.n328 VSS.n327 92.5
R13457 VSS.n991 VSS.n990 92.5
R13458 VSS.n990 VSS.t22 92.5
R13459 VSS.n345 VSS.n344 92.5
R13460 VSS.n343 VSS.n342 92.5
R13461 VSS.n341 VSS.n340 92.5
R13462 VSS.n339 VSS.n338 92.5
R13463 VSS.n337 VSS.n336 92.5
R13464 VSS.n335 VSS.n334 92.5
R13465 VSS.n333 VSS.n332 92.5
R13466 VSS.n331 VSS.n288 92.5
R13467 VSS.t22 VSS.n288 92.5
R13468 VSS.n347 VSS.n346 92.5
R13469 VSS.n349 VSS.n348 92.5
R13470 VSS.n351 VSS.n350 92.5
R13471 VSS.n353 VSS.n352 92.5
R13472 VSS.n355 VSS.n354 92.5
R13473 VSS.n357 VSS.n356 92.5
R13474 VSS.n359 VSS.n358 92.5
R13475 VSS.n361 VSS.n360 92.5
R13476 VSS.n363 VSS.n362 92.5
R13477 VSS.n364 VSS.n280 92.5
R13478 VSS.t22 VSS.n280 92.5
R13479 VSS.n908 VSS.n907 92.5
R13480 VSS.n983 VSS.n299 92.5
R13481 VSS.n974 VSS.n296 92.5
R13482 VSS.n918 VSS.n300 92.5
R13483 VSS.n922 VSS.n295 92.5
R13484 VSS.n926 VSS.n301 92.5
R13485 VSS.n930 VSS.n294 92.5
R13486 VSS.n989 VSS.n304 92.5
R13487 VSS.n936 VSS.n298 92.5
R13488 VSS.n420 VSS.n419 92.5
R13489 VSS.n369 VSS.n367 92.5
R13490 VSS.n408 VSS.n407 92.5
R13491 VSS.n410 VSS.n409 92.5
R13492 VSS.n412 VSS.n411 92.5
R13493 VSS.n414 VSS.n413 92.5
R13494 VSS.n416 VSS.n415 92.5
R13495 VSS.n418 VSS.n417 92.5
R13496 VSS.n901 VSS.n900 92.5
R13497 VSS.n900 VSS.t16 92.5
R13498 VSS.n435 VSS.n434 92.5
R13499 VSS.n433 VSS.n432 92.5
R13500 VSS.n431 VSS.n430 92.5
R13501 VSS.n429 VSS.n428 92.5
R13502 VSS.n427 VSS.n426 92.5
R13503 VSS.n425 VSS.n424 92.5
R13504 VSS.n423 VSS.n422 92.5
R13505 VSS.n421 VSS.n378 92.5
R13506 VSS.t16 VSS.n378 92.5
R13507 VSS.n437 VSS.n436 92.5
R13508 VSS.n439 VSS.n438 92.5
R13509 VSS.n441 VSS.n440 92.5
R13510 VSS.n443 VSS.n442 92.5
R13511 VSS.n445 VSS.n444 92.5
R13512 VSS.n447 VSS.n446 92.5
R13513 VSS.n449 VSS.n448 92.5
R13514 VSS.n451 VSS.n450 92.5
R13515 VSS.n453 VSS.n452 92.5
R13516 VSS.n454 VSS.n370 92.5
R13517 VSS.t16 VSS.n370 92.5
R13518 VSS.n818 VSS.n817 92.5
R13519 VSS.n893 VSS.n389 92.5
R13520 VSS.n884 VSS.n386 92.5
R13521 VSS.n828 VSS.n390 92.5
R13522 VSS.n832 VSS.n385 92.5
R13523 VSS.n836 VSS.n391 92.5
R13524 VSS.n840 VSS.n384 92.5
R13525 VSS.n899 VSS.n394 92.5
R13526 VSS.n846 VSS.n388 92.5
R13527 VSS.n510 VSS.n509 92.5
R13528 VSS.n459 VSS.n457 92.5
R13529 VSS.n498 VSS.n497 92.5
R13530 VSS.n500 VSS.n499 92.5
R13531 VSS.n502 VSS.n501 92.5
R13532 VSS.n504 VSS.n503 92.5
R13533 VSS.n506 VSS.n505 92.5
R13534 VSS.n508 VSS.n507 92.5
R13535 VSS.n811 VSS.n810 92.5
R13536 VSS.n810 VSS.t36 92.5
R13537 VSS.n525 VSS.n524 92.5
R13538 VSS.n523 VSS.n522 92.5
R13539 VSS.n521 VSS.n520 92.5
R13540 VSS.n519 VSS.n518 92.5
R13541 VSS.n517 VSS.n516 92.5
R13542 VSS.n515 VSS.n514 92.5
R13543 VSS.n513 VSS.n512 92.5
R13544 VSS.n511 VSS.n468 92.5
R13545 VSS.t36 VSS.n468 92.5
R13546 VSS.n527 VSS.n526 92.5
R13547 VSS.n529 VSS.n528 92.5
R13548 VSS.n531 VSS.n530 92.5
R13549 VSS.n533 VSS.n532 92.5
R13550 VSS.n535 VSS.n534 92.5
R13551 VSS.n537 VSS.n536 92.5
R13552 VSS.n539 VSS.n538 92.5
R13553 VSS.n541 VSS.n540 92.5
R13554 VSS.n543 VSS.n542 92.5
R13555 VSS.n544 VSS.n460 92.5
R13556 VSS.t36 VSS.n460 92.5
R13557 VSS.n728 VSS.n727 92.5
R13558 VSS.n803 VSS.n479 92.5
R13559 VSS.n794 VSS.n476 92.5
R13560 VSS.n738 VSS.n480 92.5
R13561 VSS.n742 VSS.n475 92.5
R13562 VSS.n746 VSS.n481 92.5
R13563 VSS.n750 VSS.n474 92.5
R13564 VSS.n809 VSS.n484 92.5
R13565 VSS.n756 VSS.n478 92.5
R13566 VSS.n600 VSS.n599 92.5
R13567 VSS.n549 VSS.n547 92.5
R13568 VSS.n588 VSS.n587 92.5
R13569 VSS.n590 VSS.n589 92.5
R13570 VSS.n592 VSS.n591 92.5
R13571 VSS.n594 VSS.n593 92.5
R13572 VSS.n596 VSS.n595 92.5
R13573 VSS.n598 VSS.n597 92.5
R13574 VSS.n721 VSS.n720 92.5
R13575 VSS.n720 VSS.t40 92.5
R13576 VSS.n615 VSS.n614 92.5
R13577 VSS.n613 VSS.n612 92.5
R13578 VSS.n611 VSS.n610 92.5
R13579 VSS.n609 VSS.n608 92.5
R13580 VSS.n607 VSS.n606 92.5
R13581 VSS.n605 VSS.n604 92.5
R13582 VSS.n603 VSS.n602 92.5
R13583 VSS.n601 VSS.n558 92.5
R13584 VSS.t40 VSS.n558 92.5
R13585 VSS.n617 VSS.n616 92.5
R13586 VSS.n619 VSS.n618 92.5
R13587 VSS.n621 VSS.n620 92.5
R13588 VSS.n623 VSS.n622 92.5
R13589 VSS.n625 VSS.n624 92.5
R13590 VSS.n627 VSS.n626 92.5
R13591 VSS.n629 VSS.n628 92.5
R13592 VSS.n631 VSS.n630 92.5
R13593 VSS.n633 VSS.n632 92.5
R13594 VSS.n634 VSS.n550 92.5
R13595 VSS.t40 VSS.n550 92.5
R13596 VSS.n638 VSS.n637 92.5
R13597 VSS.n713 VSS.n569 92.5
R13598 VSS.n704 VSS.n566 92.5
R13599 VSS.n648 VSS.n570 92.5
R13600 VSS.n652 VSS.n565 92.5
R13601 VSS.n656 VSS.n571 92.5
R13602 VSS.n660 VSS.n564 92.5
R13603 VSS.n719 VSS.n574 92.5
R13604 VSS.n666 VSS.n568 92.5
R13605 VSS.n14837 VSS.n14324 89.722
R13606 VSS.n14773 VSS.n14338 89.722
R13607 VSS.n15383 VSS.n14209 89.722
R13608 VSS.n14812 VSS.n14222 89.722
R13609 VSS.n14170 VSS.n14055 89.722
R13610 VSS.n15412 VSS.n14158 89.722
R13611 VSS.n15943 VSS.n14042 89.722
R13612 VSS.n13119 VSS.n12598 89.722
R13613 VSS.n13094 VSS.n12644 89.722
R13614 VSS.n13368 VSS.n11497 89.722
R13615 VSS.n13343 VSS.n12503 89.722
R13616 VSS.n12436 VSS.n11527 89.722
R13617 VSS.n11513 VSS.n11509 89.722
R13618 VSS.n12158 VSS.n12091 89.722
R13619 VSS.n8221 VSS.n7522 89.722
R13620 VSS.n7888 VSS.n7616 89.722
R13621 VSS.n8579 VSS.n7382 89.722
R13622 VSS.n8246 VSS.n7476 89.722
R13623 VSS.n8801 VSS.n7242 89.722
R13624 VSS.n8604 VSS.n7336 89.722
R13625 VSS.n8826 VSS.n6980 89.722
R13626 VSS.n4572 VSS.n4051 89.722
R13627 VSS.n4547 VSS.n4097 89.722
R13628 VSS.n4929 VSS.n3910 89.722
R13629 VSS.n4904 VSS.n3956 89.722
R13630 VSS.n5286 VSS.n3769 89.722
R13631 VSS.n5261 VSS.n3815 89.722
R13632 VSS.n5607 VSS.n3674 89.722
R13633 VSS.n2078 VSS.n1565 89.722
R13634 VSS.n2014 VSS.n1579 89.722
R13635 VSS.n2624 VSS.n1450 89.722
R13636 VSS.n2053 VSS.n1463 89.722
R13637 VSS.n1411 VSS.n1296 89.722
R13638 VSS.n2653 VSS.n1399 89.722
R13639 VSS.n17460 VSS.n16036 89.673
R13640 VSS.n11232 VSS.n11089 89.673
R13641 VSS.n11322 VSS.n10999 89.673
R13642 VSS.n11412 VSS.n10909 89.673
R13643 VSS.n13532 VSS.n10819 89.673
R13644 VSS.n13622 VSS.n10729 89.673
R13645 VSS.n13712 VSS.n10639 89.673
R13646 VSS.n13802 VSS.n10549 89.673
R13647 VSS.n13952 VSS.n10504 89.673
R13648 VSS.n9179 VSS.n8935 89.673
R13649 VSS.n6899 VSS.n6882 89.209
R13650 VSS.n14304 VSS.n14300 83.871
R13651 VSS.n14481 VSS.n14439 83.871
R13652 VSS.n15090 VSS.n15048 83.871
R13653 VSS.n14977 VSS.n14237 83.871
R13654 VSS.n15565 VSS.n14070 83.871
R13655 VSS.n15441 VSS.n14133 83.871
R13656 VSS.n15677 VSS.n15635 83.871
R13657 VSS.n13151 VSS.n12582 83.871
R13658 VSS.n13055 VSS.n12664 83.871
R13659 VSS.n11672 VSS.n11483 83.871
R13660 VSS.n13304 VSS.n12523 83.871
R13661 VSS.n11911 VSS.n11542 83.871
R13662 VSS.n11608 VSS.n11605 83.871
R13663 VSS.n11991 VSS.n11982 83.871
R13664 VSS.n8182 VSS.n7539 83.871
R13665 VSS.n7602 VSS.n7599 83.871
R13666 VSS.n8540 VSS.n7399 83.871
R13667 VSS.n7462 VSS.n7459 83.871
R13668 VSS.n8762 VSS.n7259 83.871
R13669 VSS.n7322 VSS.n7319 83.871
R13670 VSS.n7067 VSS.n6963 83.871
R13671 VSS.n4604 VSS.n4035 83.871
R13672 VSS.n4508 VSS.n4117 83.871
R13673 VSS.n4961 VSS.n3894 83.871
R13674 VSS.n4865 VSS.n3976 83.871
R13675 VSS.n5318 VSS.n3753 83.871
R13676 VSS.n5222 VSS.n3835 83.871
R13677 VSS.n5568 VSS.n3694 83.871
R13678 VSS.n1545 VSS.n1541 83.871
R13679 VSS.n1722 VSS.n1680 83.871
R13680 VSS.n2331 VSS.n2289 83.871
R13681 VSS.n2218 VSS.n1478 83.871
R13682 VSS.n2682 VSS.n1374 83.871
R13683 VSS.n2806 VSS.n1311 83.871
R13684 VSS.n17392 VSS.n16041 71.237
R13685 VSS.n17459 VSS.n17458 71.237
R13686 VSS.n17448 VSS.n16042 71.237
R13687 VSS.n17402 VSS.n16046 71.237
R13688 VSS.n17405 VSS.n16043 71.237
R13689 VSS.n17409 VSS.n16045 71.237
R13690 VSS.n17413 VSS.n16044 71.237
R13691 VSS.n17416 VSS.n16040 71.237
R13692 VSS.n17303 VSS.n17302 71.237
R13693 VSS.n17292 VSS.n16083 71.237
R13694 VSS.n17233 VSS.n16089 71.237
R13695 VSS.n17236 VSS.n16084 71.237
R13696 VSS.n17240 VSS.n16088 71.237
R13697 VSS.n17244 VSS.n16085 71.237
R13698 VSS.n16087 VSS.n16079 71.237
R13699 VSS.n17250 VSS.n16086 71.237
R13700 VSS.n17213 VSS.n17212 71.237
R13701 VSS.n17202 VSS.n16173 71.237
R13702 VSS.n17143 VSS.n16179 71.237
R13703 VSS.n17146 VSS.n16174 71.237
R13704 VSS.n17150 VSS.n16178 71.237
R13705 VSS.n17154 VSS.n16175 71.237
R13706 VSS.n16177 VSS.n16169 71.237
R13707 VSS.n17160 VSS.n16176 71.237
R13708 VSS.n17123 VSS.n17122 71.237
R13709 VSS.n17112 VSS.n16263 71.237
R13710 VSS.n17053 VSS.n16269 71.237
R13711 VSS.n17056 VSS.n16264 71.237
R13712 VSS.n17060 VSS.n16268 71.237
R13713 VSS.n17064 VSS.n16265 71.237
R13714 VSS.n16267 VSS.n16259 71.237
R13715 VSS.n17070 VSS.n16266 71.237
R13716 VSS.n17033 VSS.n17032 71.237
R13717 VSS.n17022 VSS.n16353 71.237
R13718 VSS.n16963 VSS.n16359 71.237
R13719 VSS.n16966 VSS.n16354 71.237
R13720 VSS.n16970 VSS.n16358 71.237
R13721 VSS.n16974 VSS.n16355 71.237
R13722 VSS.n16357 VSS.n16349 71.237
R13723 VSS.n16980 VSS.n16356 71.237
R13724 VSS.n16943 VSS.n16942 71.237
R13725 VSS.n16932 VSS.n16443 71.237
R13726 VSS.n16873 VSS.n16449 71.237
R13727 VSS.n16876 VSS.n16444 71.237
R13728 VSS.n16880 VSS.n16448 71.237
R13729 VSS.n16884 VSS.n16445 71.237
R13730 VSS.n16447 VSS.n16439 71.237
R13731 VSS.n16890 VSS.n16446 71.237
R13732 VSS.n16853 VSS.n16852 71.237
R13733 VSS.n16842 VSS.n16533 71.237
R13734 VSS.n16783 VSS.n16539 71.237
R13735 VSS.n16786 VSS.n16534 71.237
R13736 VSS.n16790 VSS.n16538 71.237
R13737 VSS.n16794 VSS.n16535 71.237
R13738 VSS.n16537 VSS.n16529 71.237
R13739 VSS.n16800 VSS.n16536 71.237
R13740 VSS.n16763 VSS.n16762 71.237
R13741 VSS.n16752 VSS.n16623 71.237
R13742 VSS.n16693 VSS.n16629 71.237
R13743 VSS.n16696 VSS.n16624 71.237
R13744 VSS.n16700 VSS.n16628 71.237
R13745 VSS.n16704 VSS.n16625 71.237
R13746 VSS.n16627 VSS.n16619 71.237
R13747 VSS.n16710 VSS.n16626 71.237
R13748 VSS.n11231 VSS.n11230 71.237
R13749 VSS.n11220 VSS.n11090 71.237
R13750 VSS.n11160 VSS.n11096 71.237
R13751 VSS.n11163 VSS.n11091 71.237
R13752 VSS.n11167 VSS.n11095 71.237
R13753 VSS.n11094 VSS.n11086 71.237
R13754 VSS.n11173 VSS.n11093 71.237
R13755 VSS.n11179 VSS.n11092 71.237
R13756 VSS.n11321 VSS.n11320 71.237
R13757 VSS.n11310 VSS.n11000 71.237
R13758 VSS.n11250 VSS.n11006 71.237
R13759 VSS.n11253 VSS.n11001 71.237
R13760 VSS.n11257 VSS.n11005 71.237
R13761 VSS.n11004 VSS.n10996 71.237
R13762 VSS.n11263 VSS.n11003 71.237
R13763 VSS.n11269 VSS.n11002 71.237
R13764 VSS.n11411 VSS.n11410 71.237
R13765 VSS.n11400 VSS.n10910 71.237
R13766 VSS.n11340 VSS.n10916 71.237
R13767 VSS.n11343 VSS.n10911 71.237
R13768 VSS.n11347 VSS.n10915 71.237
R13769 VSS.n10914 VSS.n10906 71.237
R13770 VSS.n11353 VSS.n10913 71.237
R13771 VSS.n11359 VSS.n10912 71.237
R13772 VSS.n13531 VSS.n13530 71.237
R13773 VSS.n13520 VSS.n10820 71.237
R13774 VSS.n13459 VSS.n10826 71.237
R13775 VSS.n13462 VSS.n10821 71.237
R13776 VSS.n13466 VSS.n10825 71.237
R13777 VSS.n10824 VSS.n10816 71.237
R13778 VSS.n13472 VSS.n10823 71.237
R13779 VSS.n13478 VSS.n10822 71.237
R13780 VSS.n13621 VSS.n13620 71.237
R13781 VSS.n13610 VSS.n10730 71.237
R13782 VSS.n13550 VSS.n10736 71.237
R13783 VSS.n13553 VSS.n10731 71.237
R13784 VSS.n13557 VSS.n10735 71.237
R13785 VSS.n10734 VSS.n10726 71.237
R13786 VSS.n13563 VSS.n10733 71.237
R13787 VSS.n13569 VSS.n10732 71.237
R13788 VSS.n13711 VSS.n13710 71.237
R13789 VSS.n13700 VSS.n10640 71.237
R13790 VSS.n13640 VSS.n10646 71.237
R13791 VSS.n13643 VSS.n10641 71.237
R13792 VSS.n13647 VSS.n10645 71.237
R13793 VSS.n10644 VSS.n10636 71.237
R13794 VSS.n13653 VSS.n10643 71.237
R13795 VSS.n13659 VSS.n10642 71.237
R13796 VSS.n13801 VSS.n13800 71.237
R13797 VSS.n13790 VSS.n10550 71.237
R13798 VSS.n13730 VSS.n10556 71.237
R13799 VSS.n13733 VSS.n10551 71.237
R13800 VSS.n13737 VSS.n10555 71.237
R13801 VSS.n10554 VSS.n10546 71.237
R13802 VSS.n13743 VSS.n10553 71.237
R13803 VSS.n13749 VSS.n10552 71.237
R13804 VSS.n13892 VSS.n10508 71.237
R13805 VSS.n13951 VSS.n13950 71.237
R13806 VSS.n13940 VSS.n10509 71.237
R13807 VSS.n13902 VSS.n10513 71.237
R13808 VSS.n13905 VSS.n10510 71.237
R13809 VSS.n13909 VSS.n10512 71.237
R13810 VSS.n13914 VSS.n10511 71.237
R13811 VSS.n13955 VSS.n10495 71.237
R13812 VSS.n9037 VSS.n9013 71.237
R13813 VSS.n9045 VSS.n9012 71.237
R13814 VSS.n9053 VSS.n9008 71.237
R13815 VSS.n9061 VSS.n9009 71.237
R13816 VSS.n9069 VSS.n9014 71.237
R13817 VSS.n9077 VSS.n9011 71.237
R13818 VSS.n9085 VSS.n9007 71.237
R13819 VSS.n9093 VSS.n9010 71.237
R13820 VSS.n10258 VSS.n10257 71.237
R13821 VSS.n10247 VSS.n9218 71.237
R13822 VSS.n10188 VSS.n9224 71.237
R13823 VSS.n10191 VSS.n9219 71.237
R13824 VSS.n10195 VSS.n9223 71.237
R13825 VSS.n10199 VSS.n9220 71.237
R13826 VSS.n9222 VSS.n9214 71.237
R13827 VSS.n10205 VSS.n9221 71.237
R13828 VSS.n10168 VSS.n10167 71.237
R13829 VSS.n10157 VSS.n9308 71.237
R13830 VSS.n10098 VSS.n9314 71.237
R13831 VSS.n10101 VSS.n9309 71.237
R13832 VSS.n10105 VSS.n9313 71.237
R13833 VSS.n10109 VSS.n9310 71.237
R13834 VSS.n9312 VSS.n9304 71.237
R13835 VSS.n10115 VSS.n9311 71.237
R13836 VSS.n10078 VSS.n10077 71.237
R13837 VSS.n10067 VSS.n9398 71.237
R13838 VSS.n10008 VSS.n9404 71.237
R13839 VSS.n10011 VSS.n9399 71.237
R13840 VSS.n10015 VSS.n9403 71.237
R13841 VSS.n10019 VSS.n9400 71.237
R13842 VSS.n9402 VSS.n9394 71.237
R13843 VSS.n10025 VSS.n9401 71.237
R13844 VSS.n9988 VSS.n9987 71.237
R13845 VSS.n9977 VSS.n9488 71.237
R13846 VSS.n9918 VSS.n9494 71.237
R13847 VSS.n9921 VSS.n9489 71.237
R13848 VSS.n9925 VSS.n9493 71.237
R13849 VSS.n9929 VSS.n9490 71.237
R13850 VSS.n9492 VSS.n9484 71.237
R13851 VSS.n9935 VSS.n9491 71.237
R13852 VSS.n9898 VSS.n9897 71.237
R13853 VSS.n9887 VSS.n9578 71.237
R13854 VSS.n9828 VSS.n9584 71.237
R13855 VSS.n9831 VSS.n9579 71.237
R13856 VSS.n9835 VSS.n9583 71.237
R13857 VSS.n9839 VSS.n9580 71.237
R13858 VSS.n9582 VSS.n9574 71.237
R13859 VSS.n9845 VSS.n9581 71.237
R13860 VSS.n9808 VSS.n9807 71.237
R13861 VSS.n9797 VSS.n9668 71.237
R13862 VSS.n9738 VSS.n9674 71.237
R13863 VSS.n9741 VSS.n9669 71.237
R13864 VSS.n9745 VSS.n9673 71.237
R13865 VSS.n9749 VSS.n9670 71.237
R13866 VSS.n9672 VSS.n9664 71.237
R13867 VSS.n9755 VSS.n9671 71.237
R13868 VSS.n9183 VSS.n9182 71.237
R13869 VSS.n10367 VSS.n10366 71.237
R13870 VSS.n10361 VSS.n10360 71.237
R13871 VSS.n10355 VSS.n10354 71.237
R13872 VSS.n10349 VSS.n10348 71.237
R13873 VSS.n10343 VSS.n10342 71.237
R13874 VSS.n10337 VSS.n10336 71.237
R13875 VSS.n10331 VSS.n10330 71.237
R13876 VSS.n5782 VSS.n5781 71.237
R13877 VSS.n5776 VSS.n5775 71.237
R13878 VSS.n5770 VSS.n5769 71.237
R13879 VSS.n5764 VSS.n5763 71.237
R13880 VSS.n5758 VSS.n5757 71.237
R13881 VSS.n5752 VSS.n5751 71.237
R13882 VSS.n5746 VSS.n5745 71.237
R13883 VSS.n5740 VSS.n5739 71.237
R13884 VSS.n5904 VSS.n5903 71.237
R13885 VSS.n5898 VSS.n5897 71.237
R13886 VSS.n5892 VSS.n5891 71.237
R13887 VSS.n5886 VSS.n5885 71.237
R13888 VSS.n5880 VSS.n5879 71.237
R13889 VSS.n5874 VSS.n5873 71.237
R13890 VSS.n5868 VSS.n5867 71.237
R13891 VSS.n5862 VSS.n5861 71.237
R13892 VSS.n6026 VSS.n6025 71.237
R13893 VSS.n6020 VSS.n6019 71.237
R13894 VSS.n6014 VSS.n6013 71.237
R13895 VSS.n6008 VSS.n6007 71.237
R13896 VSS.n6002 VSS.n6001 71.237
R13897 VSS.n5996 VSS.n5995 71.237
R13898 VSS.n5990 VSS.n5989 71.237
R13899 VSS.n5984 VSS.n5983 71.237
R13900 VSS.n6148 VSS.n6147 71.237
R13901 VSS.n6142 VSS.n6141 71.237
R13902 VSS.n6136 VSS.n6135 71.237
R13903 VSS.n6130 VSS.n6129 71.237
R13904 VSS.n6124 VSS.n6123 71.237
R13905 VSS.n6118 VSS.n6117 71.237
R13906 VSS.n6112 VSS.n6111 71.237
R13907 VSS.n6106 VSS.n6105 71.237
R13908 VSS.n6270 VSS.n6269 71.237
R13909 VSS.n6264 VSS.n6263 71.237
R13910 VSS.n6258 VSS.n6257 71.237
R13911 VSS.n6252 VSS.n6251 71.237
R13912 VSS.n6246 VSS.n6245 71.237
R13913 VSS.n6240 VSS.n6239 71.237
R13914 VSS.n6234 VSS.n6233 71.237
R13915 VSS.n6228 VSS.n6227 71.237
R13916 VSS.n6392 VSS.n6391 71.237
R13917 VSS.n6386 VSS.n6385 71.237
R13918 VSS.n6380 VSS.n6379 71.237
R13919 VSS.n6374 VSS.n6373 71.237
R13920 VSS.n6368 VSS.n6367 71.237
R13921 VSS.n6362 VSS.n6361 71.237
R13922 VSS.n6356 VSS.n6355 71.237
R13923 VSS.n6350 VSS.n6349 71.237
R13924 VSS.n6514 VSS.n6513 71.237
R13925 VSS.n6508 VSS.n6507 71.237
R13926 VSS.n6502 VSS.n6501 71.237
R13927 VSS.n6496 VSS.n6495 71.237
R13928 VSS.n6490 VSS.n6489 71.237
R13929 VSS.n6484 VSS.n6483 71.237
R13930 VSS.n6478 VSS.n6477 71.237
R13931 VSS.n6472 VSS.n6471 71.237
R13932 VSS.n6600 VSS.n3140 71.237
R13933 VSS.n3177 VSS.n3150 71.237
R13934 VSS.n3185 VSS.n3156 71.237
R13935 VSS.n3193 VSS.n3151 71.237
R13936 VSS.n3201 VSS.n3155 71.237
R13937 VSS.n3209 VSS.n3152 71.237
R13938 VSS.n3217 VSS.n3154 71.237
R13939 VSS.n3225 VSS.n3153 71.237
R13940 VSS.n1251 VSS.n1250 71.237
R13941 VSS.n1240 VSS.n35 71.237
R13942 VSS.n1186 VSS.n41 71.237
R13943 VSS.n1189 VSS.n36 71.237
R13944 VSS.n1193 VSS.n40 71.237
R13945 VSS.n1197 VSS.n37 71.237
R13946 VSS.n39 VSS.n31 71.237
R13947 VSS.n1203 VSS.n38 71.237
R13948 VSS.n1166 VSS.n1165 71.237
R13949 VSS.n1155 VSS.n126 71.237
R13950 VSS.n1096 VSS.n132 71.237
R13951 VSS.n1099 VSS.n127 71.237
R13952 VSS.n1103 VSS.n131 71.237
R13953 VSS.n1107 VSS.n128 71.237
R13954 VSS.n130 VSS.n122 71.237
R13955 VSS.n1113 VSS.n129 71.237
R13956 VSS.n1076 VSS.n1075 71.237
R13957 VSS.n1065 VSS.n216 71.237
R13958 VSS.n1006 VSS.n222 71.237
R13959 VSS.n1009 VSS.n217 71.237
R13960 VSS.n1013 VSS.n221 71.237
R13961 VSS.n1017 VSS.n218 71.237
R13962 VSS.n220 VSS.n212 71.237
R13963 VSS.n1023 VSS.n219 71.237
R13964 VSS.n986 VSS.n985 71.237
R13965 VSS.n975 VSS.n306 71.237
R13966 VSS.n916 VSS.n312 71.237
R13967 VSS.n919 VSS.n307 71.237
R13968 VSS.n923 VSS.n311 71.237
R13969 VSS.n927 VSS.n308 71.237
R13970 VSS.n310 VSS.n302 71.237
R13971 VSS.n933 VSS.n309 71.237
R13972 VSS.n896 VSS.n895 71.237
R13973 VSS.n885 VSS.n396 71.237
R13974 VSS.n826 VSS.n402 71.237
R13975 VSS.n829 VSS.n397 71.237
R13976 VSS.n833 VSS.n401 71.237
R13977 VSS.n837 VSS.n398 71.237
R13978 VSS.n400 VSS.n392 71.237
R13979 VSS.n843 VSS.n399 71.237
R13980 VSS.n806 VSS.n805 71.237
R13981 VSS.n795 VSS.n486 71.237
R13982 VSS.n736 VSS.n492 71.237
R13983 VSS.n739 VSS.n487 71.237
R13984 VSS.n743 VSS.n491 71.237
R13985 VSS.n747 VSS.n488 71.237
R13986 VSS.n490 VSS.n482 71.237
R13987 VSS.n753 VSS.n489 71.237
R13988 VSS.n716 VSS.n715 71.237
R13989 VSS.n705 VSS.n576 71.237
R13990 VSS.n646 VSS.n582 71.237
R13991 VSS.n649 VSS.n577 71.237
R13992 VSS.n653 VSS.n581 71.237
R13993 VSS.n657 VSS.n578 71.237
R13994 VSS.n580 VSS.n572 71.237
R13995 VSS.n663 VSS.n579 71.237
R13996 VSS.n14635 VSS.n14439 70.217
R13997 VSS.n15329 VSS.n14237 70.217
R13998 VSS.n14871 VSS.n14304 70.217
R13999 VSS.n15442 VSS.n15441 70.217
R14000 VSS.n15236 VSS.n15048 70.217
R14001 VSS.n15803 VSS.n15635 70.217
R14002 VSS.n15555 VSS.n14070 70.217
R14003 VSS.n13059 VSS.n12664 70.217
R14004 VSS.n13308 VSS.n12523 70.217
R14005 VSS.n12967 VSS.n12582 70.217
R14006 VSS.n11769 VSS.n11608 70.217
R14007 VSS.n11483 VSS.n11475 70.217
R14008 VSS.n12311 VSS.n11982 70.217
R14009 VSS.n12404 VSS.n11542 70.217
R14010 VSS.n7749 VSS.n7602 70.217
R14011 VSS.n8090 VSS.n7462 70.217
R14012 VSS.n8190 VSS.n7539 70.217
R14013 VSS.n8448 VSS.n7322 70.217
R14014 VSS.n8548 VSS.n7399 70.217
R14015 VSS.n8858 VSS.n6963 70.217
R14016 VSS.n8770 VSS.n7259 70.217
R14017 VSS.n4512 VSS.n4117 70.217
R14018 VSS.n4869 VSS.n3976 70.217
R14019 VSS.n4420 VSS.n4035 70.217
R14020 VSS.n5226 VSS.n3835 70.217
R14021 VSS.n4777 VSS.n3894 70.217
R14022 VSS.n5572 VSS.n3694 70.217
R14023 VSS.n5134 VSS.n3753 70.217
R14024 VSS.n1876 VSS.n1680 70.217
R14025 VSS.n2570 VSS.n1478 70.217
R14026 VSS.n2112 VSS.n1545 70.217
R14027 VSS.n2683 VSS.n2682 70.217
R14028 VSS.n2477 VSS.n2289 70.217
R14029 VSS.n2796 VSS.n1311 70.217
R14030 VSS.n14472 VSS.n14442 69.803
R14031 VSS.n14468 VSS.n14442 69.803
R14032 VSS.n14468 VSS.n14444 69.803
R14033 VSS.n14464 VSS.n14444 69.803
R14034 VSS.n14464 VSS.n14446 69.803
R14035 VSS.n14460 VSS.n14446 69.803
R14036 VSS.n14460 VSS.n14448 69.803
R14037 VSS.n14456 VSS.n14448 69.803
R14038 VSS.n14456 VSS.n14450 69.803
R14039 VSS.n14452 VSS.n14450 69.803
R14040 VSS.n14452 VSS.n14337 69.803
R14041 VSS.n14777 VSS.n14337 69.803
R14042 VSS.n14863 VSS.n14862 69.803
R14043 VSS.n14862 VSS.n14309 69.803
R14044 VSS.n14858 VSS.n14309 69.803
R14045 VSS.n14858 VSS.n14311 69.803
R14046 VSS.n14854 VSS.n14311 69.803
R14047 VSS.n14854 VSS.n14314 69.803
R14048 VSS.n14850 VSS.n14314 69.803
R14049 VSS.n14850 VSS.n14316 69.803
R14050 VSS.n14846 VSS.n14316 69.803
R14051 VSS.n14846 VSS.n14318 69.803
R14052 VSS.n14842 VSS.n14318 69.803
R14053 VSS.n14842 VSS.n14320 69.803
R14054 VSS.n15333 VSS.n14235 69.803
R14055 VSS.n15337 VSS.n14235 69.803
R14056 VSS.n15337 VSS.n14233 69.803
R14057 VSS.n15341 VSS.n14233 69.803
R14058 VSS.n15341 VSS.n14231 69.803
R14059 VSS.n15345 VSS.n14231 69.803
R14060 VSS.n15345 VSS.n14229 69.803
R14061 VSS.n15349 VSS.n14229 69.803
R14062 VSS.n15349 VSS.n14227 69.803
R14063 VSS.n15353 VSS.n14227 69.803
R14064 VSS.n15353 VSS.n14225 69.803
R14065 VSS.n15357 VSS.n14225 69.803
R14066 VSS.n15081 VSS.n15051 69.803
R14067 VSS.n15077 VSS.n15051 69.803
R14068 VSS.n15077 VSS.n15053 69.803
R14069 VSS.n15073 VSS.n15053 69.803
R14070 VSS.n15073 VSS.n15055 69.803
R14071 VSS.n15069 VSS.n15055 69.803
R14072 VSS.n15069 VSS.n15057 69.803
R14073 VSS.n15065 VSS.n15057 69.803
R14074 VSS.n15065 VSS.n15059 69.803
R14075 VSS.n15061 VSS.n15059 69.803
R14076 VSS.n15061 VSS.n14208 69.803
R14077 VSS.n15387 VSS.n14208 69.803
R14078 VSS.n15440 VSS.n14145 69.803
R14079 VSS.n15436 VSS.n14145 69.803
R14080 VSS.n15436 VSS.n14147 69.803
R14081 VSS.n15432 VSS.n14147 69.803
R14082 VSS.n15432 VSS.n14150 69.803
R14083 VSS.n15428 VSS.n14150 69.803
R14084 VSS.n15428 VSS.n14152 69.803
R14085 VSS.n15424 VSS.n14152 69.803
R14086 VSS.n15424 VSS.n14154 69.803
R14087 VSS.n15420 VSS.n14154 69.803
R14088 VSS.n15420 VSS.n14156 69.803
R14089 VSS.n15416 VSS.n14156 69.803
R14090 VSS.n15893 VSS.n14068 69.803
R14091 VSS.n15897 VSS.n14068 69.803
R14092 VSS.n15897 VSS.n14066 69.803
R14093 VSS.n15901 VSS.n14066 69.803
R14094 VSS.n15901 VSS.n14064 69.803
R14095 VSS.n15905 VSS.n14064 69.803
R14096 VSS.n15905 VSS.n14062 69.803
R14097 VSS.n15909 VSS.n14062 69.803
R14098 VSS.n15909 VSS.n14060 69.803
R14099 VSS.n15913 VSS.n14060 69.803
R14100 VSS.n15913 VSS.n14058 69.803
R14101 VSS.n15917 VSS.n14058 69.803
R14102 VSS.n15668 VSS.n15638 69.803
R14103 VSS.n15664 VSS.n15638 69.803
R14104 VSS.n15664 VSS.n15640 69.803
R14105 VSS.n15660 VSS.n15640 69.803
R14106 VSS.n15660 VSS.n15642 69.803
R14107 VSS.n15656 VSS.n15642 69.803
R14108 VSS.n15656 VSS.n15644 69.803
R14109 VSS.n15652 VSS.n15644 69.803
R14110 VSS.n15652 VSS.n15646 69.803
R14111 VSS.n15648 VSS.n15646 69.803
R14112 VSS.n15648 VSS.n14041 69.803
R14113 VSS.n15947 VSS.n14041 69.803
R14114 VSS.n13068 VSS.n12657 69.803
R14115 VSS.n13068 VSS.n12655 69.803
R14116 VSS.n13072 VSS.n12655 69.803
R14117 VSS.n13072 VSS.n12653 69.803
R14118 VSS.n13076 VSS.n12653 69.803
R14119 VSS.n13076 VSS.n12651 69.803
R14120 VSS.n13080 VSS.n12651 69.803
R14121 VSS.n13080 VSS.n12649 69.803
R14122 VSS.n13085 VSS.n12649 69.803
R14123 VSS.n13085 VSS.n12647 69.803
R14124 VSS.n13089 VSS.n12647 69.803
R14125 VSS.n13090 VSS.n13089 69.803
R14126 VSS.n13147 VSS.n12586 69.803
R14127 VSS.n13143 VSS.n12586 69.803
R14128 VSS.n13143 VSS.n12588 69.803
R14129 VSS.n13139 VSS.n12588 69.803
R14130 VSS.n13139 VSS.n12590 69.803
R14131 VSS.n13135 VSS.n12590 69.803
R14132 VSS.n13135 VSS.n12592 69.803
R14133 VSS.n13131 VSS.n12592 69.803
R14134 VSS.n13131 VSS.n12594 69.803
R14135 VSS.n13127 VSS.n12594 69.803
R14136 VSS.n13127 VSS.n12596 69.803
R14137 VSS.n13123 VSS.n12596 69.803
R14138 VSS.n13317 VSS.n12516 69.803
R14139 VSS.n13317 VSS.n12514 69.803
R14140 VSS.n13321 VSS.n12514 69.803
R14141 VSS.n13321 VSS.n12512 69.803
R14142 VSS.n13325 VSS.n12512 69.803
R14143 VSS.n13325 VSS.n12510 69.803
R14144 VSS.n13329 VSS.n12510 69.803
R14145 VSS.n13329 VSS.n12508 69.803
R14146 VSS.n13334 VSS.n12508 69.803
R14147 VSS.n13334 VSS.n12506 69.803
R14148 VSS.n13338 VSS.n12506 69.803
R14149 VSS.n13339 VSS.n13338 69.803
R14150 VSS.n13396 VSS.n11484 69.803
R14151 VSS.n13392 VSS.n11484 69.803
R14152 VSS.n13392 VSS.n11487 69.803
R14153 VSS.n13388 VSS.n11487 69.803
R14154 VSS.n13388 VSS.n11489 69.803
R14155 VSS.n13384 VSS.n11489 69.803
R14156 VSS.n13384 VSS.n11491 69.803
R14157 VSS.n13380 VSS.n11491 69.803
R14158 VSS.n13380 VSS.n11493 69.803
R14159 VSS.n13376 VSS.n11493 69.803
R14160 VSS.n13376 VSS.n11495 69.803
R14161 VSS.n13372 VSS.n11495 69.803
R14162 VSS.n11805 VSS.n11609 69.803
R14163 VSS.n11801 VSS.n11609 69.803
R14164 VSS.n11801 VSS.n11777 69.803
R14165 VSS.n11797 VSS.n11777 69.803
R14166 VSS.n11797 VSS.n11779 69.803
R14167 VSS.n11793 VSS.n11779 69.803
R14168 VSS.n11793 VSS.n11781 69.803
R14169 VSS.n11789 VSS.n11781 69.803
R14170 VSS.n11789 VSS.n11783 69.803
R14171 VSS.n11785 VSS.n11783 69.803
R14172 VSS.n11785 VSS.n11512 69.803
R14173 VSS.n12461 VSS.n11512 69.803
R14174 VSS.n12408 VSS.n11540 69.803
R14175 VSS.n12412 VSS.n11540 69.803
R14176 VSS.n12412 VSS.n11538 69.803
R14177 VSS.n12416 VSS.n11538 69.803
R14178 VSS.n12416 VSS.n11536 69.803
R14179 VSS.n12420 VSS.n11536 69.803
R14180 VSS.n12420 VSS.n11534 69.803
R14181 VSS.n12424 VSS.n11534 69.803
R14182 VSS.n12424 VSS.n11532 69.803
R14183 VSS.n12428 VSS.n11532 69.803
R14184 VSS.n12428 VSS.n11530 69.803
R14185 VSS.n12432 VSS.n11530 69.803
R14186 VSS.n12103 VSS.n12101 69.803
R14187 VSS.n12107 VSS.n12101 69.803
R14188 VSS.n12107 VSS.n12099 69.803
R14189 VSS.n12111 VSS.n12099 69.803
R14190 VSS.n12111 VSS.n12097 69.803
R14191 VSS.n12115 VSS.n12097 69.803
R14192 VSS.n12115 VSS.n12095 69.803
R14193 VSS.n12119 VSS.n12095 69.803
R14194 VSS.n12119 VSS.n12093 69.803
R14195 VSS.n12123 VSS.n12093 69.803
R14196 VSS.n12123 VSS.n12090 69.803
R14197 VSS.n12162 VSS.n12090 69.803
R14198 VSS.n7916 VSS.n7603 69.803
R14199 VSS.n7912 VSS.n7603 69.803
R14200 VSS.n7912 VSS.n7606 69.803
R14201 VSS.n7908 VSS.n7606 69.803
R14202 VSS.n7908 VSS.n7608 69.803
R14203 VSS.n7904 VSS.n7608 69.803
R14204 VSS.n7904 VSS.n7610 69.803
R14205 VSS.n7900 VSS.n7610 69.803
R14206 VSS.n7900 VSS.n7612 69.803
R14207 VSS.n7896 VSS.n7612 69.803
R14208 VSS.n7896 VSS.n7614 69.803
R14209 VSS.n7892 VSS.n7614 69.803
R14210 VSS.n8195 VSS.n7535 69.803
R14211 VSS.n8195 VSS.n7533 69.803
R14212 VSS.n8199 VSS.n7533 69.803
R14213 VSS.n8199 VSS.n7531 69.803
R14214 VSS.n8203 VSS.n7531 69.803
R14215 VSS.n8203 VSS.n7529 69.803
R14216 VSS.n8207 VSS.n7529 69.803
R14217 VSS.n8207 VSS.n7527 69.803
R14218 VSS.n8212 VSS.n7527 69.803
R14219 VSS.n8212 VSS.n7525 69.803
R14220 VSS.n8216 VSS.n7525 69.803
R14221 VSS.n8217 VSS.n8216 69.803
R14222 VSS.n8274 VSS.n7463 69.803
R14223 VSS.n8270 VSS.n7463 69.803
R14224 VSS.n8270 VSS.n7466 69.803
R14225 VSS.n8266 VSS.n7466 69.803
R14226 VSS.n8266 VSS.n7468 69.803
R14227 VSS.n8262 VSS.n7468 69.803
R14228 VSS.n8262 VSS.n7470 69.803
R14229 VSS.n8258 VSS.n7470 69.803
R14230 VSS.n8258 VSS.n7472 69.803
R14231 VSS.n8254 VSS.n7472 69.803
R14232 VSS.n8254 VSS.n7474 69.803
R14233 VSS.n8250 VSS.n7474 69.803
R14234 VSS.n8553 VSS.n7395 69.803
R14235 VSS.n8553 VSS.n7393 69.803
R14236 VSS.n8557 VSS.n7393 69.803
R14237 VSS.n8557 VSS.n7391 69.803
R14238 VSS.n8561 VSS.n7391 69.803
R14239 VSS.n8561 VSS.n7389 69.803
R14240 VSS.n8565 VSS.n7389 69.803
R14241 VSS.n8565 VSS.n7387 69.803
R14242 VSS.n8570 VSS.n7387 69.803
R14243 VSS.n8570 VSS.n7385 69.803
R14244 VSS.n8574 VSS.n7385 69.803
R14245 VSS.n8575 VSS.n8574 69.803
R14246 VSS.n8632 VSS.n7323 69.803
R14247 VSS.n8628 VSS.n7323 69.803
R14248 VSS.n8628 VSS.n7326 69.803
R14249 VSS.n8624 VSS.n7326 69.803
R14250 VSS.n8624 VSS.n7328 69.803
R14251 VSS.n8620 VSS.n7328 69.803
R14252 VSS.n8620 VSS.n7330 69.803
R14253 VSS.n8616 VSS.n7330 69.803
R14254 VSS.n8616 VSS.n7332 69.803
R14255 VSS.n8612 VSS.n7332 69.803
R14256 VSS.n8612 VSS.n7334 69.803
R14257 VSS.n8608 VSS.n7334 69.803
R14258 VSS.n8775 VSS.n7255 69.803
R14259 VSS.n8775 VSS.n7253 69.803
R14260 VSS.n8779 VSS.n7253 69.803
R14261 VSS.n8779 VSS.n7251 69.803
R14262 VSS.n8783 VSS.n7251 69.803
R14263 VSS.n8783 VSS.n7249 69.803
R14264 VSS.n8787 VSS.n7249 69.803
R14265 VSS.n8787 VSS.n7247 69.803
R14266 VSS.n8792 VSS.n7247 69.803
R14267 VSS.n8792 VSS.n7245 69.803
R14268 VSS.n8796 VSS.n7245 69.803
R14269 VSS.n8797 VSS.n8796 69.803
R14270 VSS.n8854 VSS.n6967 69.803
R14271 VSS.n8850 VSS.n6967 69.803
R14272 VSS.n8850 VSS.n6970 69.803
R14273 VSS.n8846 VSS.n6970 69.803
R14274 VSS.n8846 VSS.n6972 69.803
R14275 VSS.n8842 VSS.n6972 69.803
R14276 VSS.n8842 VSS.n6974 69.803
R14277 VSS.n8838 VSS.n6974 69.803
R14278 VSS.n8838 VSS.n6976 69.803
R14279 VSS.n8834 VSS.n6976 69.803
R14280 VSS.n8834 VSS.n6978 69.803
R14281 VSS.n8830 VSS.n6978 69.803
R14282 VSS.n4521 VSS.n4110 69.803
R14283 VSS.n4521 VSS.n4108 69.803
R14284 VSS.n4525 VSS.n4108 69.803
R14285 VSS.n4525 VSS.n4106 69.803
R14286 VSS.n4529 VSS.n4106 69.803
R14287 VSS.n4529 VSS.n4104 69.803
R14288 VSS.n4533 VSS.n4104 69.803
R14289 VSS.n4533 VSS.n4102 69.803
R14290 VSS.n4538 VSS.n4102 69.803
R14291 VSS.n4538 VSS.n4100 69.803
R14292 VSS.n4542 VSS.n4100 69.803
R14293 VSS.n4543 VSS.n4542 69.803
R14294 VSS.n4600 VSS.n4039 69.803
R14295 VSS.n4596 VSS.n4039 69.803
R14296 VSS.n4596 VSS.n4041 69.803
R14297 VSS.n4592 VSS.n4041 69.803
R14298 VSS.n4592 VSS.n4043 69.803
R14299 VSS.n4588 VSS.n4043 69.803
R14300 VSS.n4588 VSS.n4045 69.803
R14301 VSS.n4584 VSS.n4045 69.803
R14302 VSS.n4584 VSS.n4047 69.803
R14303 VSS.n4580 VSS.n4047 69.803
R14304 VSS.n4580 VSS.n4049 69.803
R14305 VSS.n4576 VSS.n4049 69.803
R14306 VSS.n4878 VSS.n3969 69.803
R14307 VSS.n4878 VSS.n3967 69.803
R14308 VSS.n4882 VSS.n3967 69.803
R14309 VSS.n4882 VSS.n3965 69.803
R14310 VSS.n4886 VSS.n3965 69.803
R14311 VSS.n4886 VSS.n3963 69.803
R14312 VSS.n4890 VSS.n3963 69.803
R14313 VSS.n4890 VSS.n3961 69.803
R14314 VSS.n4895 VSS.n3961 69.803
R14315 VSS.n4895 VSS.n3959 69.803
R14316 VSS.n4899 VSS.n3959 69.803
R14317 VSS.n4900 VSS.n4899 69.803
R14318 VSS.n4957 VSS.n3898 69.803
R14319 VSS.n4953 VSS.n3898 69.803
R14320 VSS.n4953 VSS.n3900 69.803
R14321 VSS.n4949 VSS.n3900 69.803
R14322 VSS.n4949 VSS.n3902 69.803
R14323 VSS.n4945 VSS.n3902 69.803
R14324 VSS.n4945 VSS.n3904 69.803
R14325 VSS.n4941 VSS.n3904 69.803
R14326 VSS.n4941 VSS.n3906 69.803
R14327 VSS.n4937 VSS.n3906 69.803
R14328 VSS.n4937 VSS.n3908 69.803
R14329 VSS.n4933 VSS.n3908 69.803
R14330 VSS.n5235 VSS.n3828 69.803
R14331 VSS.n5235 VSS.n3826 69.803
R14332 VSS.n5239 VSS.n3826 69.803
R14333 VSS.n5239 VSS.n3824 69.803
R14334 VSS.n5243 VSS.n3824 69.803
R14335 VSS.n5243 VSS.n3822 69.803
R14336 VSS.n5247 VSS.n3822 69.803
R14337 VSS.n5247 VSS.n3820 69.803
R14338 VSS.n5252 VSS.n3820 69.803
R14339 VSS.n5252 VSS.n3818 69.803
R14340 VSS.n5256 VSS.n3818 69.803
R14341 VSS.n5257 VSS.n5256 69.803
R14342 VSS.n5314 VSS.n3757 69.803
R14343 VSS.n5310 VSS.n3757 69.803
R14344 VSS.n5310 VSS.n3759 69.803
R14345 VSS.n5306 VSS.n3759 69.803
R14346 VSS.n5306 VSS.n3761 69.803
R14347 VSS.n5302 VSS.n3761 69.803
R14348 VSS.n5302 VSS.n3763 69.803
R14349 VSS.n5298 VSS.n3763 69.803
R14350 VSS.n5298 VSS.n3765 69.803
R14351 VSS.n5294 VSS.n3765 69.803
R14352 VSS.n5294 VSS.n3767 69.803
R14353 VSS.n5290 VSS.n3767 69.803
R14354 VSS.n5581 VSS.n3687 69.803
R14355 VSS.n5581 VSS.n3685 69.803
R14356 VSS.n5585 VSS.n3685 69.803
R14357 VSS.n5585 VSS.n3683 69.803
R14358 VSS.n5589 VSS.n3683 69.803
R14359 VSS.n5589 VSS.n3681 69.803
R14360 VSS.n5593 VSS.n3681 69.803
R14361 VSS.n5593 VSS.n3679 69.803
R14362 VSS.n5598 VSS.n3679 69.803
R14363 VSS.n5598 VSS.n3677 69.803
R14364 VSS.n5602 VSS.n3677 69.803
R14365 VSS.n5603 VSS.n5602 69.803
R14366 VSS.n1713 VSS.n1683 69.803
R14367 VSS.n1709 VSS.n1683 69.803
R14368 VSS.n1709 VSS.n1685 69.803
R14369 VSS.n1705 VSS.n1685 69.803
R14370 VSS.n1705 VSS.n1687 69.803
R14371 VSS.n1701 VSS.n1687 69.803
R14372 VSS.n1701 VSS.n1689 69.803
R14373 VSS.n1697 VSS.n1689 69.803
R14374 VSS.n1697 VSS.n1691 69.803
R14375 VSS.n1693 VSS.n1691 69.803
R14376 VSS.n1693 VSS.n1578 69.803
R14377 VSS.n2018 VSS.n1578 69.803
R14378 VSS.n2104 VSS.n2103 69.803
R14379 VSS.n2103 VSS.n1550 69.803
R14380 VSS.n2099 VSS.n1550 69.803
R14381 VSS.n2099 VSS.n1552 69.803
R14382 VSS.n2095 VSS.n1552 69.803
R14383 VSS.n2095 VSS.n1555 69.803
R14384 VSS.n2091 VSS.n1555 69.803
R14385 VSS.n2091 VSS.n1557 69.803
R14386 VSS.n2087 VSS.n1557 69.803
R14387 VSS.n2087 VSS.n1559 69.803
R14388 VSS.n2083 VSS.n1559 69.803
R14389 VSS.n2083 VSS.n1561 69.803
R14390 VSS.n2574 VSS.n1476 69.803
R14391 VSS.n2578 VSS.n1476 69.803
R14392 VSS.n2578 VSS.n1474 69.803
R14393 VSS.n2582 VSS.n1474 69.803
R14394 VSS.n2582 VSS.n1472 69.803
R14395 VSS.n2586 VSS.n1472 69.803
R14396 VSS.n2586 VSS.n1470 69.803
R14397 VSS.n2590 VSS.n1470 69.803
R14398 VSS.n2590 VSS.n1468 69.803
R14399 VSS.n2594 VSS.n1468 69.803
R14400 VSS.n2594 VSS.n1466 69.803
R14401 VSS.n2598 VSS.n1466 69.803
R14402 VSS.n2322 VSS.n2292 69.803
R14403 VSS.n2318 VSS.n2292 69.803
R14404 VSS.n2318 VSS.n2294 69.803
R14405 VSS.n2314 VSS.n2294 69.803
R14406 VSS.n2314 VSS.n2296 69.803
R14407 VSS.n2310 VSS.n2296 69.803
R14408 VSS.n2310 VSS.n2298 69.803
R14409 VSS.n2306 VSS.n2298 69.803
R14410 VSS.n2306 VSS.n2300 69.803
R14411 VSS.n2302 VSS.n2300 69.803
R14412 VSS.n2302 VSS.n1449 69.803
R14413 VSS.n2628 VSS.n1449 69.803
R14414 VSS.n2681 VSS.n1386 69.803
R14415 VSS.n2677 VSS.n1386 69.803
R14416 VSS.n2677 VSS.n1388 69.803
R14417 VSS.n2673 VSS.n1388 69.803
R14418 VSS.n2673 VSS.n1391 69.803
R14419 VSS.n2669 VSS.n1391 69.803
R14420 VSS.n2669 VSS.n1393 69.803
R14421 VSS.n2665 VSS.n1393 69.803
R14422 VSS.n2665 VSS.n1395 69.803
R14423 VSS.n2661 VSS.n1395 69.803
R14424 VSS.n2661 VSS.n1397 69.803
R14425 VSS.n2657 VSS.n1397 69.803
R14426 VSS.n2967 VSS.n1309 69.803
R14427 VSS.n2971 VSS.n1309 69.803
R14428 VSS.n2971 VSS.n1307 69.803
R14429 VSS.n2975 VSS.n1307 69.803
R14430 VSS.n2975 VSS.n1305 69.803
R14431 VSS.n2979 VSS.n1305 69.803
R14432 VSS.n2979 VSS.n1303 69.803
R14433 VSS.n2983 VSS.n1303 69.803
R14434 VSS.n2983 VSS.n1301 69.803
R14435 VSS.n2987 VSS.n1301 69.803
R14436 VSS.n2987 VSS.n1299 69.803
R14437 VSS.n2991 VSS.n1299 69.803
R14438 VSS.n6659 VSS.n6642 68.545
R14439 VSS.t14 VSS.n6648 65.818
R14440 VSS.t14 VSS.n6647 65.818
R14441 VSS.t14 VSS.n6646 65.818
R14442 VSS.t14 VSS.n6645 65.818
R14443 VSS.t14 VSS.n6644 65.818
R14444 VSS.t14 VSS.n6643 65.818
R14445 VSS.n6679 VSS.n6649 64.913
R14446 VSS.n14777 VSS.n14338 64.374
R14447 VSS.n14324 VSS.n14320 64.374
R14448 VSS.n15357 VSS.n14222 64.374
R14449 VSS.n15387 VSS.n14209 64.374
R14450 VSS.n15416 VSS.n14158 64.374
R14451 VSS.n15917 VSS.n14055 64.374
R14452 VSS.n15947 VSS.n14042 64.374
R14453 VSS.n13090 VSS.n12644 64.374
R14454 VSS.n13123 VSS.n12598 64.374
R14455 VSS.n13339 VSS.n12503 64.374
R14456 VSS.n13372 VSS.n11497 64.374
R14457 VSS.n12461 VSS.n11513 64.374
R14458 VSS.n12432 VSS.n11527 64.374
R14459 VSS.n12162 VSS.n12091 64.374
R14460 VSS.n7892 VSS.n7616 64.374
R14461 VSS.n8217 VSS.n7522 64.374
R14462 VSS.n8250 VSS.n7476 64.374
R14463 VSS.n8575 VSS.n7382 64.374
R14464 VSS.n8608 VSS.n7336 64.374
R14465 VSS.n8797 VSS.n7242 64.374
R14466 VSS.n8830 VSS.n6980 64.374
R14467 VSS.n4543 VSS.n4097 64.374
R14468 VSS.n4576 VSS.n4051 64.374
R14469 VSS.n4900 VSS.n3956 64.374
R14470 VSS.n4933 VSS.n3910 64.374
R14471 VSS.n5257 VSS.n3815 64.374
R14472 VSS.n5290 VSS.n3769 64.374
R14473 VSS.n5603 VSS.n3674 64.374
R14474 VSS.n2018 VSS.n1579 64.374
R14475 VSS.n1565 VSS.n1561 64.374
R14476 VSS.n2598 VSS.n1463 64.374
R14477 VSS.n2628 VSS.n1450 64.374
R14478 VSS.n2657 VSS.n1399 64.374
R14479 VSS.n2991 VSS.n1296 64.374
R14480 VSS.n9156 VSS.t20 59.179
R14481 VSS.n9129 VSS.n8997 53.901
R14482 VSS.n9132 VSS.n8997 53.901
R14483 VSS.n10282 VSS.n9169 53.901
R14484 VSS.n10279 VSS.n9169 53.901
R14485 VSS.n6689 VSS.n6643 53.366
R14486 VSS.n6687 VSS.n6644 53.366
R14487 VSS.n6685 VSS.n6645 53.366
R14488 VSS.n6683 VSS.n6646 53.366
R14489 VSS.n6681 VSS.n6647 53.366
R14490 VSS.n6679 VSS.n6648 53.366
R14491 VSS.n6689 VSS.n6644 53.366
R14492 VSS.n6687 VSS.n6645 53.366
R14493 VSS.n6685 VSS.n6646 53.366
R14494 VSS.n6683 VSS.n6647 53.366
R14495 VSS.n6681 VSS.n6648 53.366
R14496 VSS.n6659 VSS.n6643 53.366
R14497 VSS.n6673 VSS.n6650 53.161
R14498 VSS.n6676 VSS.n6650 53.161
R14499 VSS.n17481 VSS.n13993 47.316
R14500 VSS.n13964 VSS.n10489 47.316
R14501 VSS.n17485 VSS.n13993 46.878
R14502 VSS.n13965 VSS.n13964 46.878
R14503 VSS.n17365 VSS.n17322 41.419
R14504 VSS.n17364 VSS.n17320 41.419
R14505 VSS.n17360 VSS.n17319 41.419
R14506 VSS.n17356 VSS.n17318 41.419
R14507 VSS.n16121 VSS.n16066 41.419
R14508 VSS.n16120 VSS.n16064 41.419
R14509 VSS.n16116 VSS.n16063 41.419
R14510 VSS.n16112 VSS.n16062 41.419
R14511 VSS.n16211 VSS.n16156 41.419
R14512 VSS.n16210 VSS.n16154 41.419
R14513 VSS.n16206 VSS.n16153 41.419
R14514 VSS.n16202 VSS.n16152 41.419
R14515 VSS.n16301 VSS.n16246 41.419
R14516 VSS.n16300 VSS.n16244 41.419
R14517 VSS.n16296 VSS.n16243 41.419
R14518 VSS.n16292 VSS.n16242 41.419
R14519 VSS.n16391 VSS.n16336 41.419
R14520 VSS.n16390 VSS.n16334 41.419
R14521 VSS.n16386 VSS.n16333 41.419
R14522 VSS.n16382 VSS.n16332 41.419
R14523 VSS.n16481 VSS.n16426 41.419
R14524 VSS.n16480 VSS.n16424 41.419
R14525 VSS.n16476 VSS.n16423 41.419
R14526 VSS.n16472 VSS.n16422 41.419
R14527 VSS.n16571 VSS.n16516 41.419
R14528 VSS.n16570 VSS.n16514 41.419
R14529 VSS.n16566 VSS.n16513 41.419
R14530 VSS.n16562 VSS.n16512 41.419
R14531 VSS.n16661 VSS.n16606 41.419
R14532 VSS.n16660 VSS.n16604 41.419
R14533 VSS.n16656 VSS.n16603 41.419
R14534 VSS.n16652 VSS.n16602 41.419
R14535 VSS.n11128 VSS.n11073 41.419
R14536 VSS.n11127 VSS.n11071 41.419
R14537 VSS.n11123 VSS.n11070 41.419
R14538 VSS.n11119 VSS.n11069 41.419
R14539 VSS.n11038 VSS.n10983 41.419
R14540 VSS.n11037 VSS.n10981 41.419
R14541 VSS.n11033 VSS.n10980 41.419
R14542 VSS.n11029 VSS.n10979 41.419
R14543 VSS.n10948 VSS.n10893 41.419
R14544 VSS.n10947 VSS.n10891 41.419
R14545 VSS.n10943 VSS.n10890 41.419
R14546 VSS.n10939 VSS.n10889 41.419
R14547 VSS.n10858 VSS.n10803 41.419
R14548 VSS.n10857 VSS.n10801 41.419
R14549 VSS.n10853 VSS.n10800 41.419
R14550 VSS.n10849 VSS.n10799 41.419
R14551 VSS.n10768 VSS.n10713 41.419
R14552 VSS.n10767 VSS.n10711 41.419
R14553 VSS.n10763 VSS.n10710 41.419
R14554 VSS.n10759 VSS.n10709 41.419
R14555 VSS.n10678 VSS.n10623 41.419
R14556 VSS.n10677 VSS.n10621 41.419
R14557 VSS.n10673 VSS.n10620 41.419
R14558 VSS.n10669 VSS.n10619 41.419
R14559 VSS.n10588 VSS.n10533 41.419
R14560 VSS.n10587 VSS.n10531 41.419
R14561 VSS.n10583 VSS.n10530 41.419
R14562 VSS.n10579 VSS.n10529 41.419
R14563 VSS.n13865 VSS.n13819 41.419
R14564 VSS.n13864 VSS.n13817 41.419
R14565 VSS.n13860 VSS.n13816 41.419
R14566 VSS.n13856 VSS.n13815 41.419
R14567 VSS.n9116 VSS.n8998 41.419
R14568 VSS.n9117 VSS.n8996 41.419
R14569 VSS.n9121 VSS.n8995 41.419
R14570 VSS.n9125 VSS.n8994 41.419
R14571 VSS.n9256 VSS.n9201 41.419
R14572 VSS.n9255 VSS.n9199 41.419
R14573 VSS.n9251 VSS.n9198 41.419
R14574 VSS.n9247 VSS.n9197 41.419
R14575 VSS.n9346 VSS.n9291 41.419
R14576 VSS.n9345 VSS.n9289 41.419
R14577 VSS.n9341 VSS.n9288 41.419
R14578 VSS.n9337 VSS.n9287 41.419
R14579 VSS.n9436 VSS.n9381 41.419
R14580 VSS.n9435 VSS.n9379 41.419
R14581 VSS.n9431 VSS.n9378 41.419
R14582 VSS.n9427 VSS.n9377 41.419
R14583 VSS.n9526 VSS.n9471 41.419
R14584 VSS.n9525 VSS.n9469 41.419
R14585 VSS.n9521 VSS.n9468 41.419
R14586 VSS.n9517 VSS.n9467 41.419
R14587 VSS.n9616 VSS.n9561 41.419
R14588 VSS.n9615 VSS.n9559 41.419
R14589 VSS.n9611 VSS.n9558 41.419
R14590 VSS.n9607 VSS.n9557 41.419
R14591 VSS.n9706 VSS.n9651 41.419
R14592 VSS.n9705 VSS.n9649 41.419
R14593 VSS.n9701 VSS.n9648 41.419
R14594 VSS.n9697 VSS.n9647 41.419
R14595 VSS.n10295 VSS.n9170 41.419
R14596 VSS.n10294 VSS.n9168 41.419
R14597 VSS.n10290 VSS.n9167 41.419
R14598 VSS.n10286 VSS.n9166 41.419
R14599 VSS.n6710 VSS.n6655 41.419
R14600 VSS.n6714 VSS.n6656 41.419
R14601 VSS.n6718 VSS.n6657 41.419
R14602 VSS.n6724 VSS.n6723 41.419
R14603 VSS.n5713 VSS.n5679 41.419
R14604 VSS.n5712 VSS.n5677 41.419
R14605 VSS.n5708 VSS.n5676 41.419
R14606 VSS.n5704 VSS.n5675 41.419
R14607 VSS.n5835 VSS.n5801 41.419
R14608 VSS.n5834 VSS.n5799 41.419
R14609 VSS.n5830 VSS.n5798 41.419
R14610 VSS.n5826 VSS.n5797 41.419
R14611 VSS.n5957 VSS.n5923 41.419
R14612 VSS.n5956 VSS.n5921 41.419
R14613 VSS.n5952 VSS.n5920 41.419
R14614 VSS.n5948 VSS.n5919 41.419
R14615 VSS.n6079 VSS.n6045 41.419
R14616 VSS.n6078 VSS.n6043 41.419
R14617 VSS.n6074 VSS.n6042 41.419
R14618 VSS.n6070 VSS.n6041 41.419
R14619 VSS.n6201 VSS.n6167 41.419
R14620 VSS.n6200 VSS.n6165 41.419
R14621 VSS.n6196 VSS.n6164 41.419
R14622 VSS.n6192 VSS.n6163 41.419
R14623 VSS.n6323 VSS.n6289 41.419
R14624 VSS.n6322 VSS.n6287 41.419
R14625 VSS.n6318 VSS.n6286 41.419
R14626 VSS.n6314 VSS.n6285 41.419
R14627 VSS.n6445 VSS.n6411 41.419
R14628 VSS.n6444 VSS.n6409 41.419
R14629 VSS.n6440 VSS.n6408 41.419
R14630 VSS.n6436 VSS.n6407 41.419
R14631 VSS.n6557 VSS.n6529 41.419
R14632 VSS.n6563 VSS.n6562 41.419
R14633 VSS.n6566 VSS.n6565 41.419
R14634 VSS.n6571 VSS.n6570 41.419
R14635 VSS.n74 VSS.n18 41.419
R14636 VSS.n73 VSS.n16 41.419
R14637 VSS.n69 VSS.n15 41.419
R14638 VSS.n65 VSS.n14 41.419
R14639 VSS.n164 VSS.n109 41.419
R14640 VSS.n163 VSS.n107 41.419
R14641 VSS.n159 VSS.n106 41.419
R14642 VSS.n155 VSS.n105 41.419
R14643 VSS.n254 VSS.n199 41.419
R14644 VSS.n253 VSS.n197 41.419
R14645 VSS.n249 VSS.n196 41.419
R14646 VSS.n245 VSS.n195 41.419
R14647 VSS.n344 VSS.n289 41.419
R14648 VSS.n343 VSS.n287 41.419
R14649 VSS.n339 VSS.n286 41.419
R14650 VSS.n335 VSS.n285 41.419
R14651 VSS.n434 VSS.n379 41.419
R14652 VSS.n433 VSS.n377 41.419
R14653 VSS.n429 VSS.n376 41.419
R14654 VSS.n425 VSS.n375 41.419
R14655 VSS.n524 VSS.n469 41.419
R14656 VSS.n523 VSS.n467 41.419
R14657 VSS.n519 VSS.n466 41.419
R14658 VSS.n515 VSS.n465 41.419
R14659 VSS.n614 VSS.n559 41.419
R14660 VSS.n613 VSS.n557 41.419
R14661 VSS.n609 VSS.n556 41.419
R14662 VSS.n605 VSS.n555 41.419
R14663 VSS.n17353 VSS.n17318 41.419
R14664 VSS.n17357 VSS.n17319 41.419
R14665 VSS.n17361 VSS.n17320 41.419
R14666 VSS.n17368 VSS.n17322 41.419
R14667 VSS.n16109 VSS.n16062 41.419
R14668 VSS.n16113 VSS.n16063 41.419
R14669 VSS.n16117 VSS.n16064 41.419
R14670 VSS.n16124 VSS.n16066 41.419
R14671 VSS.n16199 VSS.n16152 41.419
R14672 VSS.n16203 VSS.n16153 41.419
R14673 VSS.n16207 VSS.n16154 41.419
R14674 VSS.n16214 VSS.n16156 41.419
R14675 VSS.n16289 VSS.n16242 41.419
R14676 VSS.n16293 VSS.n16243 41.419
R14677 VSS.n16297 VSS.n16244 41.419
R14678 VSS.n16304 VSS.n16246 41.419
R14679 VSS.n16379 VSS.n16332 41.419
R14680 VSS.n16383 VSS.n16333 41.419
R14681 VSS.n16387 VSS.n16334 41.419
R14682 VSS.n16394 VSS.n16336 41.419
R14683 VSS.n16469 VSS.n16422 41.419
R14684 VSS.n16473 VSS.n16423 41.419
R14685 VSS.n16477 VSS.n16424 41.419
R14686 VSS.n16484 VSS.n16426 41.419
R14687 VSS.n16559 VSS.n16512 41.419
R14688 VSS.n16563 VSS.n16513 41.419
R14689 VSS.n16567 VSS.n16514 41.419
R14690 VSS.n16574 VSS.n16516 41.419
R14691 VSS.n16649 VSS.n16602 41.419
R14692 VSS.n16653 VSS.n16603 41.419
R14693 VSS.n16657 VSS.n16604 41.419
R14694 VSS.n16664 VSS.n16606 41.419
R14695 VSS.n11116 VSS.n11069 41.419
R14696 VSS.n11120 VSS.n11070 41.419
R14697 VSS.n11124 VSS.n11071 41.419
R14698 VSS.n11131 VSS.n11073 41.419
R14699 VSS.n11026 VSS.n10979 41.419
R14700 VSS.n11030 VSS.n10980 41.419
R14701 VSS.n11034 VSS.n10981 41.419
R14702 VSS.n11041 VSS.n10983 41.419
R14703 VSS.n10936 VSS.n10889 41.419
R14704 VSS.n10940 VSS.n10890 41.419
R14705 VSS.n10944 VSS.n10891 41.419
R14706 VSS.n10951 VSS.n10893 41.419
R14707 VSS.n10846 VSS.n10799 41.419
R14708 VSS.n10850 VSS.n10800 41.419
R14709 VSS.n10854 VSS.n10801 41.419
R14710 VSS.n10861 VSS.n10803 41.419
R14711 VSS.n10756 VSS.n10709 41.419
R14712 VSS.n10760 VSS.n10710 41.419
R14713 VSS.n10764 VSS.n10711 41.419
R14714 VSS.n10771 VSS.n10713 41.419
R14715 VSS.n10666 VSS.n10619 41.419
R14716 VSS.n10670 VSS.n10620 41.419
R14717 VSS.n10674 VSS.n10621 41.419
R14718 VSS.n10681 VSS.n10623 41.419
R14719 VSS.n10576 VSS.n10529 41.419
R14720 VSS.n10580 VSS.n10530 41.419
R14721 VSS.n10584 VSS.n10531 41.419
R14722 VSS.n10591 VSS.n10533 41.419
R14723 VSS.n13853 VSS.n13815 41.419
R14724 VSS.n13857 VSS.n13816 41.419
R14725 VSS.n13861 VSS.n13817 41.419
R14726 VSS.n13868 VSS.n13819 41.419
R14727 VSS.n9128 VSS.n8994 41.419
R14728 VSS.n9124 VSS.n8995 41.419
R14729 VSS.n9120 VSS.n8996 41.419
R14730 VSS.n9113 VSS.n8998 41.419
R14731 VSS.n9244 VSS.n9197 41.419
R14732 VSS.n9248 VSS.n9198 41.419
R14733 VSS.n9252 VSS.n9199 41.419
R14734 VSS.n9259 VSS.n9201 41.419
R14735 VSS.n9334 VSS.n9287 41.419
R14736 VSS.n9338 VSS.n9288 41.419
R14737 VSS.n9342 VSS.n9289 41.419
R14738 VSS.n9349 VSS.n9291 41.419
R14739 VSS.n9424 VSS.n9377 41.419
R14740 VSS.n9428 VSS.n9378 41.419
R14741 VSS.n9432 VSS.n9379 41.419
R14742 VSS.n9439 VSS.n9381 41.419
R14743 VSS.n9514 VSS.n9467 41.419
R14744 VSS.n9518 VSS.n9468 41.419
R14745 VSS.n9522 VSS.n9469 41.419
R14746 VSS.n9529 VSS.n9471 41.419
R14747 VSS.n9604 VSS.n9557 41.419
R14748 VSS.n9608 VSS.n9558 41.419
R14749 VSS.n9612 VSS.n9559 41.419
R14750 VSS.n9619 VSS.n9561 41.419
R14751 VSS.n9694 VSS.n9647 41.419
R14752 VSS.n9698 VSS.n9648 41.419
R14753 VSS.n9702 VSS.n9649 41.419
R14754 VSS.n9709 VSS.n9651 41.419
R14755 VSS.n10283 VSS.n9166 41.419
R14756 VSS.n10287 VSS.n9167 41.419
R14757 VSS.n10291 VSS.n9168 41.419
R14758 VSS.n10297 VSS.n9170 41.419
R14759 VSS.n6724 VSS.n6638 41.419
R14760 VSS.n6658 VSS.n6657 41.419
R14761 VSS.n6717 VSS.n6656 41.419
R14762 VSS.n6713 VSS.n6655 41.419
R14763 VSS.n5701 VSS.n5675 41.419
R14764 VSS.n5705 VSS.n5676 41.419
R14765 VSS.n5709 VSS.n5677 41.419
R14766 VSS.n5716 VSS.n5679 41.419
R14767 VSS.n5823 VSS.n5797 41.419
R14768 VSS.n5827 VSS.n5798 41.419
R14769 VSS.n5831 VSS.n5799 41.419
R14770 VSS.n5838 VSS.n5801 41.419
R14771 VSS.n5945 VSS.n5919 41.419
R14772 VSS.n5949 VSS.n5920 41.419
R14773 VSS.n5953 VSS.n5921 41.419
R14774 VSS.n5960 VSS.n5923 41.419
R14775 VSS.n6067 VSS.n6041 41.419
R14776 VSS.n6071 VSS.n6042 41.419
R14777 VSS.n6075 VSS.n6043 41.419
R14778 VSS.n6082 VSS.n6045 41.419
R14779 VSS.n6189 VSS.n6163 41.419
R14780 VSS.n6193 VSS.n6164 41.419
R14781 VSS.n6197 VSS.n6165 41.419
R14782 VSS.n6204 VSS.n6167 41.419
R14783 VSS.n6311 VSS.n6285 41.419
R14784 VSS.n6315 VSS.n6286 41.419
R14785 VSS.n6319 VSS.n6287 41.419
R14786 VSS.n6326 VSS.n6289 41.419
R14787 VSS.n6433 VSS.n6407 41.419
R14788 VSS.n6437 VSS.n6408 41.419
R14789 VSS.n6441 VSS.n6409 41.419
R14790 VSS.n6448 VSS.n6411 41.419
R14791 VSS.n6572 VSS.n6571 41.419
R14792 VSS.n6565 VSS.n6527 41.419
R14793 VSS.n6564 VSS.n6563 41.419
R14794 VSS.n6558 VSS.n6557 41.419
R14795 VSS.n62 VSS.n14 41.419
R14796 VSS.n66 VSS.n15 41.419
R14797 VSS.n70 VSS.n16 41.419
R14798 VSS.n77 VSS.n18 41.419
R14799 VSS.n152 VSS.n105 41.419
R14800 VSS.n156 VSS.n106 41.419
R14801 VSS.n160 VSS.n107 41.419
R14802 VSS.n167 VSS.n109 41.419
R14803 VSS.n242 VSS.n195 41.419
R14804 VSS.n246 VSS.n196 41.419
R14805 VSS.n250 VSS.n197 41.419
R14806 VSS.n257 VSS.n199 41.419
R14807 VSS.n332 VSS.n285 41.419
R14808 VSS.n336 VSS.n286 41.419
R14809 VSS.n340 VSS.n287 41.419
R14810 VSS.n347 VSS.n289 41.419
R14811 VSS.n422 VSS.n375 41.419
R14812 VSS.n426 VSS.n376 41.419
R14813 VSS.n430 VSS.n377 41.419
R14814 VSS.n437 VSS.n379 41.419
R14815 VSS.n512 VSS.n465 41.419
R14816 VSS.n516 VSS.n466 41.419
R14817 VSS.n520 VSS.n467 41.419
R14818 VSS.n527 VSS.n469 41.419
R14819 VSS.n602 VSS.n555 41.419
R14820 VSS.n606 VSS.n556 41.419
R14821 VSS.n610 VSS.n557 41.419
R14822 VSS.n617 VSS.n559 41.419
R14823 VSS.n17384 VSS.n17383 41.418
R14824 VSS.n17379 VSS.n17325 41.418
R14825 VSS.n17376 VSS.n17324 41.418
R14826 VSS.n17372 VSS.n17323 41.418
R14827 VSS.n17336 VSS.n17314 41.418
R14828 VSS.n17340 VSS.n17315 41.418
R14829 VSS.n17344 VSS.n17316 41.418
R14830 VSS.n17348 VSS.n17317 41.418
R14831 VSS.n17339 VSS.n17314 41.418
R14832 VSS.n17343 VSS.n17315 41.418
R14833 VSS.n17347 VSS.n17316 41.418
R14834 VSS.n17350 VSS.n17317 41.418
R14835 VSS.n17369 VSS.n17323 41.418
R14836 VSS.n17373 VSS.n17324 41.418
R14837 VSS.n17377 VSS.n17325 41.418
R14838 VSS.n17384 VSS.n17326 41.418
R14839 VSS.n16139 VSS.n16070 41.418
R14840 VSS.n16136 VSS.n16069 41.418
R14841 VSS.n16132 VSS.n16068 41.418
R14842 VSS.n16128 VSS.n16067 41.418
R14843 VSS.n16058 VSS.n16056 41.418
R14844 VSS.n16096 VSS.n16059 41.418
R14845 VSS.n16100 VSS.n16060 41.418
R14846 VSS.n16104 VSS.n16061 41.418
R14847 VSS.n16095 VSS.n16058 41.418
R14848 VSS.n16099 VSS.n16059 41.418
R14849 VSS.n16103 VSS.n16060 41.418
R14850 VSS.n16106 VSS.n16061 41.418
R14851 VSS.n16125 VSS.n16067 41.418
R14852 VSS.n16129 VSS.n16068 41.418
R14853 VSS.n16133 VSS.n16069 41.418
R14854 VSS.n16137 VSS.n16070 41.418
R14855 VSS.n16229 VSS.n16160 41.418
R14856 VSS.n16226 VSS.n16159 41.418
R14857 VSS.n16222 VSS.n16158 41.418
R14858 VSS.n16218 VSS.n16157 41.418
R14859 VSS.n16148 VSS.n16146 41.418
R14860 VSS.n16186 VSS.n16149 41.418
R14861 VSS.n16190 VSS.n16150 41.418
R14862 VSS.n16194 VSS.n16151 41.418
R14863 VSS.n16185 VSS.n16148 41.418
R14864 VSS.n16189 VSS.n16149 41.418
R14865 VSS.n16193 VSS.n16150 41.418
R14866 VSS.n16196 VSS.n16151 41.418
R14867 VSS.n16215 VSS.n16157 41.418
R14868 VSS.n16219 VSS.n16158 41.418
R14869 VSS.n16223 VSS.n16159 41.418
R14870 VSS.n16227 VSS.n16160 41.418
R14871 VSS.n16319 VSS.n16250 41.418
R14872 VSS.n16316 VSS.n16249 41.418
R14873 VSS.n16312 VSS.n16248 41.418
R14874 VSS.n16308 VSS.n16247 41.418
R14875 VSS.n16238 VSS.n16236 41.418
R14876 VSS.n16276 VSS.n16239 41.418
R14877 VSS.n16280 VSS.n16240 41.418
R14878 VSS.n16284 VSS.n16241 41.418
R14879 VSS.n16275 VSS.n16238 41.418
R14880 VSS.n16279 VSS.n16239 41.418
R14881 VSS.n16283 VSS.n16240 41.418
R14882 VSS.n16286 VSS.n16241 41.418
R14883 VSS.n16305 VSS.n16247 41.418
R14884 VSS.n16309 VSS.n16248 41.418
R14885 VSS.n16313 VSS.n16249 41.418
R14886 VSS.n16317 VSS.n16250 41.418
R14887 VSS.n16409 VSS.n16340 41.418
R14888 VSS.n16406 VSS.n16339 41.418
R14889 VSS.n16402 VSS.n16338 41.418
R14890 VSS.n16398 VSS.n16337 41.418
R14891 VSS.n16328 VSS.n16326 41.418
R14892 VSS.n16366 VSS.n16329 41.418
R14893 VSS.n16370 VSS.n16330 41.418
R14894 VSS.n16374 VSS.n16331 41.418
R14895 VSS.n16365 VSS.n16328 41.418
R14896 VSS.n16369 VSS.n16329 41.418
R14897 VSS.n16373 VSS.n16330 41.418
R14898 VSS.n16376 VSS.n16331 41.418
R14899 VSS.n16395 VSS.n16337 41.418
R14900 VSS.n16399 VSS.n16338 41.418
R14901 VSS.n16403 VSS.n16339 41.418
R14902 VSS.n16407 VSS.n16340 41.418
R14903 VSS.n16499 VSS.n16430 41.418
R14904 VSS.n16496 VSS.n16429 41.418
R14905 VSS.n16492 VSS.n16428 41.418
R14906 VSS.n16488 VSS.n16427 41.418
R14907 VSS.n16418 VSS.n16416 41.418
R14908 VSS.n16456 VSS.n16419 41.418
R14909 VSS.n16460 VSS.n16420 41.418
R14910 VSS.n16464 VSS.n16421 41.418
R14911 VSS.n16455 VSS.n16418 41.418
R14912 VSS.n16459 VSS.n16419 41.418
R14913 VSS.n16463 VSS.n16420 41.418
R14914 VSS.n16466 VSS.n16421 41.418
R14915 VSS.n16485 VSS.n16427 41.418
R14916 VSS.n16489 VSS.n16428 41.418
R14917 VSS.n16493 VSS.n16429 41.418
R14918 VSS.n16497 VSS.n16430 41.418
R14919 VSS.n16589 VSS.n16520 41.418
R14920 VSS.n16586 VSS.n16519 41.418
R14921 VSS.n16582 VSS.n16518 41.418
R14922 VSS.n16578 VSS.n16517 41.418
R14923 VSS.n16508 VSS.n16506 41.418
R14924 VSS.n16546 VSS.n16509 41.418
R14925 VSS.n16550 VSS.n16510 41.418
R14926 VSS.n16554 VSS.n16511 41.418
R14927 VSS.n16545 VSS.n16508 41.418
R14928 VSS.n16549 VSS.n16509 41.418
R14929 VSS.n16553 VSS.n16510 41.418
R14930 VSS.n16556 VSS.n16511 41.418
R14931 VSS.n16575 VSS.n16517 41.418
R14932 VSS.n16579 VSS.n16518 41.418
R14933 VSS.n16583 VSS.n16519 41.418
R14934 VSS.n16587 VSS.n16520 41.418
R14935 VSS.n16679 VSS.n16610 41.418
R14936 VSS.n16676 VSS.n16609 41.418
R14937 VSS.n16672 VSS.n16608 41.418
R14938 VSS.n16668 VSS.n16607 41.418
R14939 VSS.n16598 VSS.n16596 41.418
R14940 VSS.n16636 VSS.n16599 41.418
R14941 VSS.n16640 VSS.n16600 41.418
R14942 VSS.n16644 VSS.n16601 41.418
R14943 VSS.n16635 VSS.n16598 41.418
R14944 VSS.n16639 VSS.n16599 41.418
R14945 VSS.n16643 VSS.n16600 41.418
R14946 VSS.n16646 VSS.n16601 41.418
R14947 VSS.n16665 VSS.n16607 41.418
R14948 VSS.n16669 VSS.n16608 41.418
R14949 VSS.n16673 VSS.n16609 41.418
R14950 VSS.n16677 VSS.n16610 41.418
R14951 VSS.n11146 VSS.n11077 41.418
R14952 VSS.n11143 VSS.n11076 41.418
R14953 VSS.n11139 VSS.n11075 41.418
R14954 VSS.n11135 VSS.n11074 41.418
R14955 VSS.n11065 VSS.n11063 41.418
R14956 VSS.n11103 VSS.n11066 41.418
R14957 VSS.n11107 VSS.n11067 41.418
R14958 VSS.n11111 VSS.n11068 41.418
R14959 VSS.n11102 VSS.n11065 41.418
R14960 VSS.n11106 VSS.n11066 41.418
R14961 VSS.n11110 VSS.n11067 41.418
R14962 VSS.n11113 VSS.n11068 41.418
R14963 VSS.n11132 VSS.n11074 41.418
R14964 VSS.n11136 VSS.n11075 41.418
R14965 VSS.n11140 VSS.n11076 41.418
R14966 VSS.n11144 VSS.n11077 41.418
R14967 VSS.n11056 VSS.n10987 41.418
R14968 VSS.n11053 VSS.n10986 41.418
R14969 VSS.n11049 VSS.n10985 41.418
R14970 VSS.n11045 VSS.n10984 41.418
R14971 VSS.n10975 VSS.n10973 41.418
R14972 VSS.n11013 VSS.n10976 41.418
R14973 VSS.n11017 VSS.n10977 41.418
R14974 VSS.n11021 VSS.n10978 41.418
R14975 VSS.n11012 VSS.n10975 41.418
R14976 VSS.n11016 VSS.n10976 41.418
R14977 VSS.n11020 VSS.n10977 41.418
R14978 VSS.n11023 VSS.n10978 41.418
R14979 VSS.n11042 VSS.n10984 41.418
R14980 VSS.n11046 VSS.n10985 41.418
R14981 VSS.n11050 VSS.n10986 41.418
R14982 VSS.n11054 VSS.n10987 41.418
R14983 VSS.n10966 VSS.n10897 41.418
R14984 VSS.n10963 VSS.n10896 41.418
R14985 VSS.n10959 VSS.n10895 41.418
R14986 VSS.n10955 VSS.n10894 41.418
R14987 VSS.n10885 VSS.n10883 41.418
R14988 VSS.n10923 VSS.n10886 41.418
R14989 VSS.n10927 VSS.n10887 41.418
R14990 VSS.n10931 VSS.n10888 41.418
R14991 VSS.n10922 VSS.n10885 41.418
R14992 VSS.n10926 VSS.n10886 41.418
R14993 VSS.n10930 VSS.n10887 41.418
R14994 VSS.n10933 VSS.n10888 41.418
R14995 VSS.n10952 VSS.n10894 41.418
R14996 VSS.n10956 VSS.n10895 41.418
R14997 VSS.n10960 VSS.n10896 41.418
R14998 VSS.n10964 VSS.n10897 41.418
R14999 VSS.n10876 VSS.n10807 41.418
R15000 VSS.n10873 VSS.n10806 41.418
R15001 VSS.n10869 VSS.n10805 41.418
R15002 VSS.n10865 VSS.n10804 41.418
R15003 VSS.n10795 VSS.n10793 41.418
R15004 VSS.n10833 VSS.n10796 41.418
R15005 VSS.n10837 VSS.n10797 41.418
R15006 VSS.n10841 VSS.n10798 41.418
R15007 VSS.n10832 VSS.n10795 41.418
R15008 VSS.n10836 VSS.n10796 41.418
R15009 VSS.n10840 VSS.n10797 41.418
R15010 VSS.n10843 VSS.n10798 41.418
R15011 VSS.n10862 VSS.n10804 41.418
R15012 VSS.n10866 VSS.n10805 41.418
R15013 VSS.n10870 VSS.n10806 41.418
R15014 VSS.n10874 VSS.n10807 41.418
R15015 VSS.n10786 VSS.n10717 41.418
R15016 VSS.n10783 VSS.n10716 41.418
R15017 VSS.n10779 VSS.n10715 41.418
R15018 VSS.n10775 VSS.n10714 41.418
R15019 VSS.n10705 VSS.n10703 41.418
R15020 VSS.n10743 VSS.n10706 41.418
R15021 VSS.n10747 VSS.n10707 41.418
R15022 VSS.n10751 VSS.n10708 41.418
R15023 VSS.n10742 VSS.n10705 41.418
R15024 VSS.n10746 VSS.n10706 41.418
R15025 VSS.n10750 VSS.n10707 41.418
R15026 VSS.n10753 VSS.n10708 41.418
R15027 VSS.n10772 VSS.n10714 41.418
R15028 VSS.n10776 VSS.n10715 41.418
R15029 VSS.n10780 VSS.n10716 41.418
R15030 VSS.n10784 VSS.n10717 41.418
R15031 VSS.n10696 VSS.n10627 41.418
R15032 VSS.n10693 VSS.n10626 41.418
R15033 VSS.n10689 VSS.n10625 41.418
R15034 VSS.n10685 VSS.n10624 41.418
R15035 VSS.n10615 VSS.n10613 41.418
R15036 VSS.n10653 VSS.n10616 41.418
R15037 VSS.n10657 VSS.n10617 41.418
R15038 VSS.n10661 VSS.n10618 41.418
R15039 VSS.n10652 VSS.n10615 41.418
R15040 VSS.n10656 VSS.n10616 41.418
R15041 VSS.n10660 VSS.n10617 41.418
R15042 VSS.n10663 VSS.n10618 41.418
R15043 VSS.n10682 VSS.n10624 41.418
R15044 VSS.n10686 VSS.n10625 41.418
R15045 VSS.n10690 VSS.n10626 41.418
R15046 VSS.n10694 VSS.n10627 41.418
R15047 VSS.n10606 VSS.n10537 41.418
R15048 VSS.n10603 VSS.n10536 41.418
R15049 VSS.n10599 VSS.n10535 41.418
R15050 VSS.n10595 VSS.n10534 41.418
R15051 VSS.n10525 VSS.n10523 41.418
R15052 VSS.n10563 VSS.n10526 41.418
R15053 VSS.n10567 VSS.n10527 41.418
R15054 VSS.n10571 VSS.n10528 41.418
R15055 VSS.n10562 VSS.n10525 41.418
R15056 VSS.n10566 VSS.n10526 41.418
R15057 VSS.n10570 VSS.n10527 41.418
R15058 VSS.n10573 VSS.n10528 41.418
R15059 VSS.n10592 VSS.n10534 41.418
R15060 VSS.n10596 VSS.n10535 41.418
R15061 VSS.n10600 VSS.n10536 41.418
R15062 VSS.n10604 VSS.n10537 41.418
R15063 VSS.n13884 VSS.n13883 41.418
R15064 VSS.n13879 VSS.n13822 41.418
R15065 VSS.n13876 VSS.n13821 41.418
R15066 VSS.n13872 VSS.n13820 41.418
R15067 VSS.n13836 VSS.n13811 41.418
R15068 VSS.n13840 VSS.n13812 41.418
R15069 VSS.n13844 VSS.n13813 41.418
R15070 VSS.n13848 VSS.n13814 41.418
R15071 VSS.n13839 VSS.n13811 41.418
R15072 VSS.n13843 VSS.n13812 41.418
R15073 VSS.n13847 VSS.n13813 41.418
R15074 VSS.n13850 VSS.n13814 41.418
R15075 VSS.n13869 VSS.n13820 41.418
R15076 VSS.n13873 VSS.n13821 41.418
R15077 VSS.n13877 VSS.n13822 41.418
R15078 VSS.n13884 VSS.n13823 41.418
R15079 VSS.n9099 VSS.n9005 41.418
R15080 VSS.n9103 VSS.n9003 41.418
R15081 VSS.n9107 VSS.n9001 41.418
R15082 VSS.n9110 VSS.n8999 41.418
R15083 VSS.n9145 VSS.n9006 41.418
R15084 VSS.n9141 VSS.n9004 41.418
R15085 VSS.n9137 VSS.n9002 41.418
R15086 VSS.n9133 VSS.n9000 41.418
R15087 VSS.n9144 VSS.n9004 41.418
R15088 VSS.n9140 VSS.n9002 41.418
R15089 VSS.n9136 VSS.n9000 41.418
R15090 VSS.n9016 VSS.n9006 41.418
R15091 VSS.n9005 VSS.n8984 41.418
R15092 VSS.n9100 VSS.n9003 41.418
R15093 VSS.n9104 VSS.n9001 41.418
R15094 VSS.n9108 VSS.n8999 41.418
R15095 VSS.n9274 VSS.n9205 41.418
R15096 VSS.n9271 VSS.n9204 41.418
R15097 VSS.n9267 VSS.n9203 41.418
R15098 VSS.n9263 VSS.n9202 41.418
R15099 VSS.n9193 VSS.n9191 41.418
R15100 VSS.n9231 VSS.n9194 41.418
R15101 VSS.n9235 VSS.n9195 41.418
R15102 VSS.n9239 VSS.n9196 41.418
R15103 VSS.n9230 VSS.n9193 41.418
R15104 VSS.n9234 VSS.n9194 41.418
R15105 VSS.n9238 VSS.n9195 41.418
R15106 VSS.n9241 VSS.n9196 41.418
R15107 VSS.n9260 VSS.n9202 41.418
R15108 VSS.n9264 VSS.n9203 41.418
R15109 VSS.n9268 VSS.n9204 41.418
R15110 VSS.n9272 VSS.n9205 41.418
R15111 VSS.n9364 VSS.n9295 41.418
R15112 VSS.n9361 VSS.n9294 41.418
R15113 VSS.n9357 VSS.n9293 41.418
R15114 VSS.n9353 VSS.n9292 41.418
R15115 VSS.n9283 VSS.n9281 41.418
R15116 VSS.n9321 VSS.n9284 41.418
R15117 VSS.n9325 VSS.n9285 41.418
R15118 VSS.n9329 VSS.n9286 41.418
R15119 VSS.n9320 VSS.n9283 41.418
R15120 VSS.n9324 VSS.n9284 41.418
R15121 VSS.n9328 VSS.n9285 41.418
R15122 VSS.n9331 VSS.n9286 41.418
R15123 VSS.n9350 VSS.n9292 41.418
R15124 VSS.n9354 VSS.n9293 41.418
R15125 VSS.n9358 VSS.n9294 41.418
R15126 VSS.n9362 VSS.n9295 41.418
R15127 VSS.n9454 VSS.n9385 41.418
R15128 VSS.n9451 VSS.n9384 41.418
R15129 VSS.n9447 VSS.n9383 41.418
R15130 VSS.n9443 VSS.n9382 41.418
R15131 VSS.n9373 VSS.n9371 41.418
R15132 VSS.n9411 VSS.n9374 41.418
R15133 VSS.n9415 VSS.n9375 41.418
R15134 VSS.n9419 VSS.n9376 41.418
R15135 VSS.n9410 VSS.n9373 41.418
R15136 VSS.n9414 VSS.n9374 41.418
R15137 VSS.n9418 VSS.n9375 41.418
R15138 VSS.n9421 VSS.n9376 41.418
R15139 VSS.n9440 VSS.n9382 41.418
R15140 VSS.n9444 VSS.n9383 41.418
R15141 VSS.n9448 VSS.n9384 41.418
R15142 VSS.n9452 VSS.n9385 41.418
R15143 VSS.n9544 VSS.n9475 41.418
R15144 VSS.n9541 VSS.n9474 41.418
R15145 VSS.n9537 VSS.n9473 41.418
R15146 VSS.n9533 VSS.n9472 41.418
R15147 VSS.n9463 VSS.n9461 41.418
R15148 VSS.n9501 VSS.n9464 41.418
R15149 VSS.n9505 VSS.n9465 41.418
R15150 VSS.n9509 VSS.n9466 41.418
R15151 VSS.n9500 VSS.n9463 41.418
R15152 VSS.n9504 VSS.n9464 41.418
R15153 VSS.n9508 VSS.n9465 41.418
R15154 VSS.n9511 VSS.n9466 41.418
R15155 VSS.n9530 VSS.n9472 41.418
R15156 VSS.n9534 VSS.n9473 41.418
R15157 VSS.n9538 VSS.n9474 41.418
R15158 VSS.n9542 VSS.n9475 41.418
R15159 VSS.n9634 VSS.n9565 41.418
R15160 VSS.n9631 VSS.n9564 41.418
R15161 VSS.n9627 VSS.n9563 41.418
R15162 VSS.n9623 VSS.n9562 41.418
R15163 VSS.n9553 VSS.n9551 41.418
R15164 VSS.n9591 VSS.n9554 41.418
R15165 VSS.n9595 VSS.n9555 41.418
R15166 VSS.n9599 VSS.n9556 41.418
R15167 VSS.n9590 VSS.n9553 41.418
R15168 VSS.n9594 VSS.n9554 41.418
R15169 VSS.n9598 VSS.n9555 41.418
R15170 VSS.n9601 VSS.n9556 41.418
R15171 VSS.n9620 VSS.n9562 41.418
R15172 VSS.n9624 VSS.n9563 41.418
R15173 VSS.n9628 VSS.n9564 41.418
R15174 VSS.n9632 VSS.n9565 41.418
R15175 VSS.n9724 VSS.n9655 41.418
R15176 VSS.n9721 VSS.n9654 41.418
R15177 VSS.n9717 VSS.n9653 41.418
R15178 VSS.n9713 VSS.n9652 41.418
R15179 VSS.n9643 VSS.n9641 41.418
R15180 VSS.n9681 VSS.n9644 41.418
R15181 VSS.n9685 VSS.n9645 41.418
R15182 VSS.n9689 VSS.n9646 41.418
R15183 VSS.n9680 VSS.n9643 41.418
R15184 VSS.n9684 VSS.n9644 41.418
R15185 VSS.n9688 VSS.n9645 41.418
R15186 VSS.n9691 VSS.n9646 41.418
R15187 VSS.n9710 VSS.n9652 41.418
R15188 VSS.n9714 VSS.n9653 41.418
R15189 VSS.n9718 VSS.n9654 41.418
R15190 VSS.n9722 VSS.n9655 41.418
R15191 VSS.n10312 VSS.n9177 41.418
R15192 VSS.n10308 VSS.n9175 41.418
R15193 VSS.n10304 VSS.n9173 41.418
R15194 VSS.n10300 VSS.n9171 41.418
R15195 VSS.n10324 VSS.n9164 41.418
R15196 VSS.n10270 VSS.n9176 41.418
R15197 VSS.n10274 VSS.n9174 41.418
R15198 VSS.n10278 VSS.n9172 41.418
R15199 VSS.n10267 VSS.n9176 41.418
R15200 VSS.n10271 VSS.n9174 41.418
R15201 VSS.n10275 VSS.n9172 41.418
R15202 VSS.n10325 VSS.n10324 41.418
R15203 VSS.n10315 VSS.n9177 41.418
R15204 VSS.n10311 VSS.n9175 41.418
R15205 VSS.n10307 VSS.n9173 41.418
R15206 VSS.n10303 VSS.n9171 41.418
R15207 VSS.n6697 VSS.n6641 41.418
R15208 VSS.n6698 VSS.n6651 41.418
R15209 VSS.n6705 VSS.n6640 41.418
R15210 VSS.n6709 VSS.n6639 41.418
R15211 VSS.n6669 VSS.n6652 41.418
R15212 VSS.n6665 VSS.n6653 41.418
R15213 VSS.n6661 VSS.n6654 41.418
R15214 VSS.n6726 VSS.n6637 41.418
R15215 VSS.n6694 VSS.n6641 41.418
R15216 VSS.n6701 VSS.n6651 41.418
R15217 VSS.n6702 VSS.n6640 41.418
R15218 VSS.n6706 VSS.n6639 41.418
R15219 VSS.n6672 VSS.n6652 41.418
R15220 VSS.n6668 VSS.n6653 41.418
R15221 VSS.n6664 VSS.n6654 41.418
R15222 VSS.n6660 VSS.n6637 41.418
R15223 VSS.n5732 VSS.n5731 41.418
R15224 VSS.n5727 VSS.n5682 41.418
R15225 VSS.n5724 VSS.n5681 41.418
R15226 VSS.n5720 VSS.n5680 41.418
R15227 VSS.n5671 VSS.n3631 41.418
R15228 VSS.n5688 VSS.n5672 41.418
R15229 VSS.n5692 VSS.n5673 41.418
R15230 VSS.n5696 VSS.n5674 41.418
R15231 VSS.n5687 VSS.n5671 41.418
R15232 VSS.n5691 VSS.n5672 41.418
R15233 VSS.n5695 VSS.n5673 41.418
R15234 VSS.n5698 VSS.n5674 41.418
R15235 VSS.n5717 VSS.n5680 41.418
R15236 VSS.n5721 VSS.n5681 41.418
R15237 VSS.n5725 VSS.n5682 41.418
R15238 VSS.n5732 VSS.n5683 41.418
R15239 VSS.n5854 VSS.n5853 41.418
R15240 VSS.n5849 VSS.n5804 41.418
R15241 VSS.n5846 VSS.n5803 41.418
R15242 VSS.n5842 VSS.n5802 41.418
R15243 VSS.n5793 VSS.n3573 41.418
R15244 VSS.n5810 VSS.n5794 41.418
R15245 VSS.n5814 VSS.n5795 41.418
R15246 VSS.n5818 VSS.n5796 41.418
R15247 VSS.n5809 VSS.n5793 41.418
R15248 VSS.n5813 VSS.n5794 41.418
R15249 VSS.n5817 VSS.n5795 41.418
R15250 VSS.n5820 VSS.n5796 41.418
R15251 VSS.n5839 VSS.n5802 41.418
R15252 VSS.n5843 VSS.n5803 41.418
R15253 VSS.n5847 VSS.n5804 41.418
R15254 VSS.n5854 VSS.n5805 41.418
R15255 VSS.n5976 VSS.n5975 41.418
R15256 VSS.n5971 VSS.n5926 41.418
R15257 VSS.n5968 VSS.n5925 41.418
R15258 VSS.n5964 VSS.n5924 41.418
R15259 VSS.n5915 VSS.n3515 41.418
R15260 VSS.n5932 VSS.n5916 41.418
R15261 VSS.n5936 VSS.n5917 41.418
R15262 VSS.n5940 VSS.n5918 41.418
R15263 VSS.n5931 VSS.n5915 41.418
R15264 VSS.n5935 VSS.n5916 41.418
R15265 VSS.n5939 VSS.n5917 41.418
R15266 VSS.n5942 VSS.n5918 41.418
R15267 VSS.n5961 VSS.n5924 41.418
R15268 VSS.n5965 VSS.n5925 41.418
R15269 VSS.n5969 VSS.n5926 41.418
R15270 VSS.n5976 VSS.n5927 41.418
R15271 VSS.n6098 VSS.n6097 41.418
R15272 VSS.n6093 VSS.n6048 41.418
R15273 VSS.n6090 VSS.n6047 41.418
R15274 VSS.n6086 VSS.n6046 41.418
R15275 VSS.n6037 VSS.n3457 41.418
R15276 VSS.n6054 VSS.n6038 41.418
R15277 VSS.n6058 VSS.n6039 41.418
R15278 VSS.n6062 VSS.n6040 41.418
R15279 VSS.n6053 VSS.n6037 41.418
R15280 VSS.n6057 VSS.n6038 41.418
R15281 VSS.n6061 VSS.n6039 41.418
R15282 VSS.n6064 VSS.n6040 41.418
R15283 VSS.n6083 VSS.n6046 41.418
R15284 VSS.n6087 VSS.n6047 41.418
R15285 VSS.n6091 VSS.n6048 41.418
R15286 VSS.n6098 VSS.n6049 41.418
R15287 VSS.n6220 VSS.n6219 41.418
R15288 VSS.n6215 VSS.n6170 41.418
R15289 VSS.n6212 VSS.n6169 41.418
R15290 VSS.n6208 VSS.n6168 41.418
R15291 VSS.n6159 VSS.n3399 41.418
R15292 VSS.n6176 VSS.n6160 41.418
R15293 VSS.n6180 VSS.n6161 41.418
R15294 VSS.n6184 VSS.n6162 41.418
R15295 VSS.n6175 VSS.n6159 41.418
R15296 VSS.n6179 VSS.n6160 41.418
R15297 VSS.n6183 VSS.n6161 41.418
R15298 VSS.n6186 VSS.n6162 41.418
R15299 VSS.n6205 VSS.n6168 41.418
R15300 VSS.n6209 VSS.n6169 41.418
R15301 VSS.n6213 VSS.n6170 41.418
R15302 VSS.n6220 VSS.n6171 41.418
R15303 VSS.n6342 VSS.n6341 41.418
R15304 VSS.n6337 VSS.n6292 41.418
R15305 VSS.n6334 VSS.n6291 41.418
R15306 VSS.n6330 VSS.n6290 41.418
R15307 VSS.n6281 VSS.n3341 41.418
R15308 VSS.n6298 VSS.n6282 41.418
R15309 VSS.n6302 VSS.n6283 41.418
R15310 VSS.n6306 VSS.n6284 41.418
R15311 VSS.n6297 VSS.n6281 41.418
R15312 VSS.n6301 VSS.n6282 41.418
R15313 VSS.n6305 VSS.n6283 41.418
R15314 VSS.n6308 VSS.n6284 41.418
R15315 VSS.n6327 VSS.n6290 41.418
R15316 VSS.n6331 VSS.n6291 41.418
R15317 VSS.n6335 VSS.n6292 41.418
R15318 VSS.n6342 VSS.n6293 41.418
R15319 VSS.n6464 VSS.n6463 41.418
R15320 VSS.n6459 VSS.n6414 41.418
R15321 VSS.n6456 VSS.n6413 41.418
R15322 VSS.n6452 VSS.n6412 41.418
R15323 VSS.n6403 VSS.n3283 41.418
R15324 VSS.n6420 VSS.n6404 41.418
R15325 VSS.n6424 VSS.n6405 41.418
R15326 VSS.n6428 VSS.n6406 41.418
R15327 VSS.n6419 VSS.n6403 41.418
R15328 VSS.n6423 VSS.n6404 41.418
R15329 VSS.n6427 VSS.n6405 41.418
R15330 VSS.n6430 VSS.n6406 41.418
R15331 VSS.n6449 VSS.n6412 41.418
R15332 VSS.n6453 VSS.n6413 41.418
R15333 VSS.n6457 VSS.n6414 41.418
R15334 VSS.n6464 VSS.n6415 41.418
R15335 VSS.n6542 VSS.n6541 41.418
R15336 VSS.n6547 VSS.n6546 41.418
R15337 VSS.n6550 VSS.n6549 41.418
R15338 VSS.n6555 VSS.n6554 41.418
R15339 VSS.n6587 VSS.n6586 41.418
R15340 VSS.n6584 VSS.n6521 41.418
R15341 VSS.n6580 VSS.n6579 41.418
R15342 VSS.n6524 VSS.n6523 41.418
R15343 VSS.n6586 VSS.n6585 41.418
R15344 VSS.n6581 VSS.n6521 41.418
R15345 VSS.n6579 VSS.n6578 41.418
R15346 VSS.n6525 VSS.n6524 41.418
R15347 VSS.n6556 VSS.n6555 41.418
R15348 VSS.n6549 VSS.n6531 41.418
R15349 VSS.n6548 VSS.n6547 41.418
R15350 VSS.n6541 VSS.n6533 41.418
R15351 VSS.n92 VSS.n22 41.418
R15352 VSS.n89 VSS.n21 41.418
R15353 VSS.n85 VSS.n20 41.418
R15354 VSS.n81 VSS.n19 41.418
R15355 VSS.n10 VSS.n8 41.418
R15356 VSS.n49 VSS.n11 41.418
R15357 VSS.n53 VSS.n12 41.418
R15358 VSS.n57 VSS.n13 41.418
R15359 VSS.n48 VSS.n10 41.418
R15360 VSS.n52 VSS.n11 41.418
R15361 VSS.n56 VSS.n12 41.418
R15362 VSS.n59 VSS.n13 41.418
R15363 VSS.n78 VSS.n19 41.418
R15364 VSS.n82 VSS.n20 41.418
R15365 VSS.n86 VSS.n21 41.418
R15366 VSS.n90 VSS.n22 41.418
R15367 VSS.n182 VSS.n113 41.418
R15368 VSS.n179 VSS.n112 41.418
R15369 VSS.n175 VSS.n111 41.418
R15370 VSS.n171 VSS.n110 41.418
R15371 VSS.n101 VSS.n99 41.418
R15372 VSS.n139 VSS.n102 41.418
R15373 VSS.n143 VSS.n103 41.418
R15374 VSS.n147 VSS.n104 41.418
R15375 VSS.n138 VSS.n101 41.418
R15376 VSS.n142 VSS.n102 41.418
R15377 VSS.n146 VSS.n103 41.418
R15378 VSS.n149 VSS.n104 41.418
R15379 VSS.n168 VSS.n110 41.418
R15380 VSS.n172 VSS.n111 41.418
R15381 VSS.n176 VSS.n112 41.418
R15382 VSS.n180 VSS.n113 41.418
R15383 VSS.n272 VSS.n203 41.418
R15384 VSS.n269 VSS.n202 41.418
R15385 VSS.n265 VSS.n201 41.418
R15386 VSS.n261 VSS.n200 41.418
R15387 VSS.n191 VSS.n189 41.418
R15388 VSS.n229 VSS.n192 41.418
R15389 VSS.n233 VSS.n193 41.418
R15390 VSS.n237 VSS.n194 41.418
R15391 VSS.n228 VSS.n191 41.418
R15392 VSS.n232 VSS.n192 41.418
R15393 VSS.n236 VSS.n193 41.418
R15394 VSS.n239 VSS.n194 41.418
R15395 VSS.n258 VSS.n200 41.418
R15396 VSS.n262 VSS.n201 41.418
R15397 VSS.n266 VSS.n202 41.418
R15398 VSS.n270 VSS.n203 41.418
R15399 VSS.n362 VSS.n293 41.418
R15400 VSS.n359 VSS.n292 41.418
R15401 VSS.n355 VSS.n291 41.418
R15402 VSS.n351 VSS.n290 41.418
R15403 VSS.n281 VSS.n279 41.418
R15404 VSS.n319 VSS.n282 41.418
R15405 VSS.n323 VSS.n283 41.418
R15406 VSS.n327 VSS.n284 41.418
R15407 VSS.n318 VSS.n281 41.418
R15408 VSS.n322 VSS.n282 41.418
R15409 VSS.n326 VSS.n283 41.418
R15410 VSS.n329 VSS.n284 41.418
R15411 VSS.n348 VSS.n290 41.418
R15412 VSS.n352 VSS.n291 41.418
R15413 VSS.n356 VSS.n292 41.418
R15414 VSS.n360 VSS.n293 41.418
R15415 VSS.n452 VSS.n383 41.418
R15416 VSS.n449 VSS.n382 41.418
R15417 VSS.n445 VSS.n381 41.418
R15418 VSS.n441 VSS.n380 41.418
R15419 VSS.n371 VSS.n369 41.418
R15420 VSS.n409 VSS.n372 41.418
R15421 VSS.n413 VSS.n373 41.418
R15422 VSS.n417 VSS.n374 41.418
R15423 VSS.n408 VSS.n371 41.418
R15424 VSS.n412 VSS.n372 41.418
R15425 VSS.n416 VSS.n373 41.418
R15426 VSS.n419 VSS.n374 41.418
R15427 VSS.n438 VSS.n380 41.418
R15428 VSS.n442 VSS.n381 41.418
R15429 VSS.n446 VSS.n382 41.418
R15430 VSS.n450 VSS.n383 41.418
R15431 VSS.n542 VSS.n473 41.418
R15432 VSS.n539 VSS.n472 41.418
R15433 VSS.n535 VSS.n471 41.418
R15434 VSS.n531 VSS.n470 41.418
R15435 VSS.n461 VSS.n459 41.418
R15436 VSS.n499 VSS.n462 41.418
R15437 VSS.n503 VSS.n463 41.418
R15438 VSS.n507 VSS.n464 41.418
R15439 VSS.n498 VSS.n461 41.418
R15440 VSS.n502 VSS.n462 41.418
R15441 VSS.n506 VSS.n463 41.418
R15442 VSS.n509 VSS.n464 41.418
R15443 VSS.n528 VSS.n470 41.418
R15444 VSS.n532 VSS.n471 41.418
R15445 VSS.n536 VSS.n472 41.418
R15446 VSS.n540 VSS.n473 41.418
R15447 VSS.n632 VSS.n563 41.418
R15448 VSS.n629 VSS.n562 41.418
R15449 VSS.n625 VSS.n561 41.418
R15450 VSS.n621 VSS.n560 41.418
R15451 VSS.n551 VSS.n549 41.418
R15452 VSS.n589 VSS.n552 41.418
R15453 VSS.n593 VSS.n553 41.418
R15454 VSS.n597 VSS.n554 41.418
R15455 VSS.n588 VSS.n551 41.418
R15456 VSS.n592 VSS.n552 41.418
R15457 VSS.n596 VSS.n553 41.418
R15458 VSS.n599 VSS.n554 41.418
R15459 VSS.n618 VSS.n560 41.418
R15460 VSS.n622 VSS.n561 41.418
R15461 VSS.n626 VSS.n562 41.418
R15462 VSS.n630 VSS.n563 41.418
R15463 VSS.t14 VSS.n6649 40.03
R15464 VSS.t14 VSS.n6642 38.819
R15465 VSS.n6693 VSS.n6642 34.273
R15466 VSS.n3058 sky130_asc_pfet_01v8_lvt_60_1/VGND 33.334
R15467 VSS.n6677 VSS.n6649 32.457
R15468 VSS.n17705 VSS 32.416
R15469 sky130_asc_pfet_01v8_lvt_6_1/VGND sky130_asc_pfet_01v8_lvt_60_2/VGND 29.082
R15470 VSS.n17352 VSS.n17351 27.554
R15471 VSS.n16108 VSS.n16107 27.554
R15472 VSS.n16198 VSS.n16197 27.554
R15473 VSS.n16288 VSS.n16287 27.554
R15474 VSS.n16378 VSS.n16377 27.554
R15475 VSS.n16468 VSS.n16467 27.554
R15476 VSS.n16558 VSS.n16557 27.554
R15477 VSS.n16648 VSS.n16647 27.554
R15478 VSS.n11115 VSS.n11114 27.554
R15479 VSS.n11025 VSS.n11024 27.554
R15480 VSS.n10935 VSS.n10934 27.554
R15481 VSS.n10845 VSS.n10844 27.554
R15482 VSS.n10755 VSS.n10754 27.554
R15483 VSS.n10665 VSS.n10664 27.554
R15484 VSS.n10575 VSS.n10574 27.554
R15485 VSS.n13852 VSS.n13851 27.554
R15486 VSS.n9131 VSS.n9130 27.554
R15487 VSS.n9243 VSS.n9242 27.554
R15488 VSS.n9333 VSS.n9332 27.554
R15489 VSS.n9423 VSS.n9422 27.554
R15490 VSS.n9513 VSS.n9512 27.554
R15491 VSS.n9603 VSS.n9602 27.554
R15492 VSS.n9693 VSS.n9692 27.554
R15493 VSS.n10281 VSS.n10280 27.554
R15494 VSS.n5700 VSS.n5699 27.554
R15495 VSS.n5822 VSS.n5821 27.554
R15496 VSS.n5944 VSS.n5943 27.554
R15497 VSS.n6066 VSS.n6065 27.554
R15498 VSS.n6188 VSS.n6187 27.554
R15499 VSS.n6310 VSS.n6309 27.554
R15500 VSS.n6432 VSS.n6431 27.554
R15501 VSS.n6575 VSS.n6574 27.554
R15502 VSS.n61 VSS.n60 27.554
R15503 VSS.n151 VSS.n150 27.554
R15504 VSS.n241 VSS.n240 27.554
R15505 VSS.n331 VSS.n330 27.554
R15506 VSS.n421 VSS.n420 27.554
R15507 VSS.n511 VSS.n510 27.554
R15508 VSS.n601 VSS.n600 27.554
R15509 VSS.n17370 VSS.n17367 26.666
R15510 VSS.n16126 VSS.n16123 26.666
R15511 VSS.n16216 VSS.n16213 26.666
R15512 VSS.n16306 VSS.n16303 26.666
R15513 VSS.n16396 VSS.n16393 26.666
R15514 VSS.n16486 VSS.n16483 26.666
R15515 VSS.n16576 VSS.n16573 26.666
R15516 VSS.n16666 VSS.n16663 26.666
R15517 VSS.n11133 VSS.n11130 26.666
R15518 VSS.n11043 VSS.n11040 26.666
R15519 VSS.n10953 VSS.n10950 26.666
R15520 VSS.n10863 VSS.n10860 26.666
R15521 VSS.n10773 VSS.n10770 26.666
R15522 VSS.n10683 VSS.n10680 26.666
R15523 VSS.n10593 VSS.n10590 26.666
R15524 VSS.n13870 VSS.n13867 26.666
R15525 VSS.n9114 VSS.n9112 26.666
R15526 VSS.n9261 VSS.n9258 26.666
R15527 VSS.n9351 VSS.n9348 26.666
R15528 VSS.n9441 VSS.n9438 26.666
R15529 VSS.n9531 VSS.n9528 26.666
R15530 VSS.n9621 VSS.n9618 26.666
R15531 VSS.n9711 VSS.n9708 26.666
R15532 VSS.n10299 VSS.n10298 26.666
R15533 VSS.n6675 VSS.n6674 26.666
R15534 VSS.n5718 VSS.n5715 26.666
R15535 VSS.n5840 VSS.n5837 26.666
R15536 VSS.n5962 VSS.n5959 26.666
R15537 VSS.n6084 VSS.n6081 26.666
R15538 VSS.n6206 VSS.n6203 26.666
R15539 VSS.n6328 VSS.n6325 26.666
R15540 VSS.n6450 VSS.n6447 26.666
R15541 VSS.n6559 VSS.n6530 26.666
R15542 VSS.n79 VSS.n76 26.666
R15543 VSS.n169 VSS.n166 26.666
R15544 VSS.n259 VSS.n256 26.666
R15545 VSS.n349 VSS.n346 26.666
R15546 VSS.n439 VSS.n436 26.666
R15547 VSS.n529 VSS.n526 26.666
R15548 VSS.n619 VSS.n616 26.666
R15549 VSS.n17680 VSS.n17650 25.831
R15550 VSS.n10464 VSS.n10463 25.831
R15551 VSS.t30 VSS.n17320 25.542
R15552 VSS.t30 VSS.n17319 25.542
R15553 VSS.t30 VSS.n17318 25.542
R15554 VSS.t30 VSS.n17322 25.542
R15555 VSS.t54 VSS.n16064 25.542
R15556 VSS.t54 VSS.n16063 25.542
R15557 VSS.t54 VSS.n16062 25.542
R15558 VSS.t54 VSS.n16066 25.542
R15559 VSS.t50 VSS.n16154 25.542
R15560 VSS.t50 VSS.n16153 25.542
R15561 VSS.t50 VSS.n16152 25.542
R15562 VSS.t50 VSS.n16156 25.542
R15563 VSS.t42 VSS.n16244 25.542
R15564 VSS.t42 VSS.n16243 25.542
R15565 VSS.t42 VSS.n16242 25.542
R15566 VSS.t42 VSS.n16246 25.542
R15567 VSS.t68 VSS.n16334 25.542
R15568 VSS.t68 VSS.n16333 25.542
R15569 VSS.t68 VSS.n16332 25.542
R15570 VSS.t68 VSS.n16336 25.542
R15571 VSS.t74 VSS.n16424 25.542
R15572 VSS.t74 VSS.n16423 25.542
R15573 VSS.t74 VSS.n16422 25.542
R15574 VSS.t74 VSS.n16426 25.542
R15575 VSS.t90 VSS.n16514 25.542
R15576 VSS.t90 VSS.n16513 25.542
R15577 VSS.t90 VSS.n16512 25.542
R15578 VSS.t90 VSS.n16516 25.542
R15579 VSS.t28 VSS.n16604 25.542
R15580 VSS.t28 VSS.n16603 25.542
R15581 VSS.t28 VSS.n16602 25.542
R15582 VSS.t28 VSS.n16606 25.542
R15583 VSS.t58 VSS.n11071 25.542
R15584 VSS.t58 VSS.n11070 25.542
R15585 VSS.t58 VSS.n11069 25.542
R15586 VSS.t58 VSS.n11073 25.542
R15587 VSS.t32 VSS.n10981 25.542
R15588 VSS.t32 VSS.n10980 25.542
R15589 VSS.t32 VSS.n10979 25.542
R15590 VSS.t32 VSS.n10983 25.542
R15591 VSS.t92 VSS.n10891 25.542
R15592 VSS.t92 VSS.n10890 25.542
R15593 VSS.t92 VSS.n10889 25.542
R15594 VSS.t92 VSS.n10893 25.542
R15595 VSS.t88 VSS.n10801 25.542
R15596 VSS.t88 VSS.n10800 25.542
R15597 VSS.t88 VSS.n10799 25.542
R15598 VSS.t88 VSS.n10803 25.542
R15599 VSS.t72 VSS.n10711 25.542
R15600 VSS.t72 VSS.n10710 25.542
R15601 VSS.t72 VSS.n10709 25.542
R15602 VSS.t72 VSS.n10713 25.542
R15603 VSS.t78 VSS.n10621 25.542
R15604 VSS.t78 VSS.n10620 25.542
R15605 VSS.t78 VSS.n10619 25.542
R15606 VSS.t78 VSS.n10623 25.542
R15607 VSS.t82 VSS.n10531 25.542
R15608 VSS.t82 VSS.n10530 25.542
R15609 VSS.t82 VSS.n10529 25.542
R15610 VSS.t82 VSS.n10533 25.542
R15611 VSS.t62 VSS.n13817 25.542
R15612 VSS.t62 VSS.n13816 25.542
R15613 VSS.t62 VSS.n13815 25.542
R15614 VSS.t62 VSS.n13819 25.542
R15615 VSS.t20 VSS.n8996 25.542
R15616 VSS.t20 VSS.n8995 25.542
R15617 VSS.t20 VSS.n8994 25.542
R15618 VSS.t20 VSS.n8998 25.542
R15619 VSS.t34 VSS.n9199 25.542
R15620 VSS.t34 VSS.n9198 25.542
R15621 VSS.t34 VSS.n9197 25.542
R15622 VSS.t34 VSS.n9201 25.542
R15623 VSS.t26 VSS.n9289 25.542
R15624 VSS.t26 VSS.n9288 25.542
R15625 VSS.t26 VSS.n9287 25.542
R15626 VSS.t26 VSS.n9291 25.542
R15627 VSS.t52 VSS.n9379 25.542
R15628 VSS.t52 VSS.n9378 25.542
R15629 VSS.t52 VSS.n9377 25.542
R15630 VSS.t52 VSS.n9381 25.542
R15631 VSS.t56 VSS.n9469 25.542
R15632 VSS.t56 VSS.n9468 25.542
R15633 VSS.t56 VSS.n9467 25.542
R15634 VSS.t56 VSS.n9471 25.542
R15635 VSS.t80 VSS.n9559 25.542
R15636 VSS.t80 VSS.n9558 25.542
R15637 VSS.t80 VSS.n9557 25.542
R15638 VSS.t80 VSS.n9561 25.542
R15639 VSS.t18 VSS.n9649 25.542
R15640 VSS.t18 VSS.n9648 25.542
R15641 VSS.t18 VSS.n9647 25.542
R15642 VSS.t18 VSS.n9651 25.542
R15643 VSS.t38 VSS.n9168 25.542
R15644 VSS.t38 VSS.n9167 25.542
R15645 VSS.t38 VSS.n9166 25.542
R15646 VSS.t38 VSS.n9170 25.542
R15647 VSS.t14 VSS.n6655 25.542
R15648 VSS.t14 VSS.n6656 25.542
R15649 VSS.t14 VSS.n6657 25.542
R15650 VSS.t14 VSS.n6724 25.542
R15651 VSS.t46 VSS.n5677 25.542
R15652 VSS.t46 VSS.n5676 25.542
R15653 VSS.t46 VSS.n5675 25.542
R15654 VSS.t46 VSS.n5679 25.542
R15655 VSS.t70 VSS.n5799 25.542
R15656 VSS.t70 VSS.n5798 25.542
R15657 VSS.t70 VSS.n5797 25.542
R15658 VSS.t70 VSS.n5801 25.542
R15659 VSS.t66 VSS.n5921 25.542
R15660 VSS.t66 VSS.n5920 25.542
R15661 VSS.t66 VSS.n5919 25.542
R15662 VSS.t66 VSS.n5923 25.542
R15663 VSS.t64 VSS.n6043 25.542
R15664 VSS.t64 VSS.n6042 25.542
R15665 VSS.t64 VSS.n6041 25.542
R15666 VSS.t64 VSS.n6045 25.542
R15667 VSS.t84 VSS.n6165 25.542
R15668 VSS.t84 VSS.n6164 25.542
R15669 VSS.t84 VSS.n6163 25.542
R15670 VSS.t84 VSS.n6167 25.542
R15671 VSS.t86 VSS.n6287 25.542
R15672 VSS.t86 VSS.n6286 25.542
R15673 VSS.t86 VSS.n6285 25.542
R15674 VSS.t86 VSS.n6289 25.542
R15675 VSS.t24 VSS.n6409 25.542
R15676 VSS.t24 VSS.n6408 25.542
R15677 VSS.t24 VSS.n6407 25.542
R15678 VSS.t24 VSS.n6411 25.542
R15679 VSS.n6563 VSS.t44 25.542
R15680 VSS.n6565 VSS.t44 25.542
R15681 VSS.n6571 VSS.t44 25.542
R15682 VSS.n6557 VSS.t44 25.542
R15683 VSS.t60 VSS.n16 25.542
R15684 VSS.t60 VSS.n15 25.542
R15685 VSS.t60 VSS.n14 25.542
R15686 VSS.t60 VSS.n18 25.542
R15687 VSS.t48 VSS.n107 25.542
R15688 VSS.t48 VSS.n106 25.542
R15689 VSS.t48 VSS.n105 25.542
R15690 VSS.t48 VSS.n109 25.542
R15691 VSS.t76 VSS.n197 25.542
R15692 VSS.t76 VSS.n196 25.542
R15693 VSS.t76 VSS.n195 25.542
R15694 VSS.t76 VSS.n199 25.542
R15695 VSS.t22 VSS.n287 25.542
R15696 VSS.t22 VSS.n286 25.542
R15697 VSS.t22 VSS.n285 25.542
R15698 VSS.t22 VSS.n289 25.542
R15699 VSS.t16 VSS.n377 25.542
R15700 VSS.t16 VSS.n376 25.542
R15701 VSS.t16 VSS.n375 25.542
R15702 VSS.t16 VSS.n379 25.542
R15703 VSS.t36 VSS.n467 25.542
R15704 VSS.t36 VSS.n466 25.542
R15705 VSS.t36 VSS.n465 25.542
R15706 VSS.t36 VSS.n469 25.542
R15707 VSS.t40 VSS.n557 25.542
R15708 VSS.t40 VSS.n556 25.542
R15709 VSS.t40 VSS.n555 25.542
R15710 VSS.t40 VSS.n559 25.542
R15711 VSS.t30 VSS.n17314 25.542
R15712 VSS.t30 VSS.n17315 25.542
R15713 VSS.t30 VSS.n17316 25.542
R15714 VSS.t30 VSS.n17317 25.542
R15715 VSS.t30 VSS.n17323 25.542
R15716 VSS.t30 VSS.n17324 25.542
R15717 VSS.t30 VSS.n17325 25.542
R15718 VSS.t30 VSS.n17384 25.542
R15719 VSS.t54 VSS.n16058 25.542
R15720 VSS.t54 VSS.n16059 25.542
R15721 VSS.t54 VSS.n16060 25.542
R15722 VSS.t54 VSS.n16061 25.542
R15723 VSS.t54 VSS.n16067 25.542
R15724 VSS.t54 VSS.n16068 25.542
R15725 VSS.t54 VSS.n16069 25.542
R15726 VSS.t54 VSS.n16070 25.542
R15727 VSS.t50 VSS.n16148 25.542
R15728 VSS.t50 VSS.n16149 25.542
R15729 VSS.t50 VSS.n16150 25.542
R15730 VSS.t50 VSS.n16151 25.542
R15731 VSS.t50 VSS.n16157 25.542
R15732 VSS.t50 VSS.n16158 25.542
R15733 VSS.t50 VSS.n16159 25.542
R15734 VSS.t50 VSS.n16160 25.542
R15735 VSS.t42 VSS.n16238 25.542
R15736 VSS.t42 VSS.n16239 25.542
R15737 VSS.t42 VSS.n16240 25.542
R15738 VSS.t42 VSS.n16241 25.542
R15739 VSS.t42 VSS.n16247 25.542
R15740 VSS.t42 VSS.n16248 25.542
R15741 VSS.t42 VSS.n16249 25.542
R15742 VSS.t42 VSS.n16250 25.542
R15743 VSS.t68 VSS.n16328 25.542
R15744 VSS.t68 VSS.n16329 25.542
R15745 VSS.t68 VSS.n16330 25.542
R15746 VSS.t68 VSS.n16331 25.542
R15747 VSS.t68 VSS.n16337 25.542
R15748 VSS.t68 VSS.n16338 25.542
R15749 VSS.t68 VSS.n16339 25.542
R15750 VSS.t68 VSS.n16340 25.542
R15751 VSS.t74 VSS.n16418 25.542
R15752 VSS.t74 VSS.n16419 25.542
R15753 VSS.t74 VSS.n16420 25.542
R15754 VSS.t74 VSS.n16421 25.542
R15755 VSS.t74 VSS.n16427 25.542
R15756 VSS.t74 VSS.n16428 25.542
R15757 VSS.t74 VSS.n16429 25.542
R15758 VSS.t74 VSS.n16430 25.542
R15759 VSS.t90 VSS.n16508 25.542
R15760 VSS.t90 VSS.n16509 25.542
R15761 VSS.t90 VSS.n16510 25.542
R15762 VSS.t90 VSS.n16511 25.542
R15763 VSS.t90 VSS.n16517 25.542
R15764 VSS.t90 VSS.n16518 25.542
R15765 VSS.t90 VSS.n16519 25.542
R15766 VSS.t90 VSS.n16520 25.542
R15767 VSS.t28 VSS.n16598 25.542
R15768 VSS.t28 VSS.n16599 25.542
R15769 VSS.t28 VSS.n16600 25.542
R15770 VSS.t28 VSS.n16601 25.542
R15771 VSS.t28 VSS.n16607 25.542
R15772 VSS.t28 VSS.n16608 25.542
R15773 VSS.t28 VSS.n16609 25.542
R15774 VSS.t28 VSS.n16610 25.542
R15775 VSS.t58 VSS.n11065 25.542
R15776 VSS.t58 VSS.n11066 25.542
R15777 VSS.t58 VSS.n11067 25.542
R15778 VSS.t58 VSS.n11068 25.542
R15779 VSS.t58 VSS.n11074 25.542
R15780 VSS.t58 VSS.n11075 25.542
R15781 VSS.t58 VSS.n11076 25.542
R15782 VSS.t58 VSS.n11077 25.542
R15783 VSS.t32 VSS.n10975 25.542
R15784 VSS.t32 VSS.n10976 25.542
R15785 VSS.t32 VSS.n10977 25.542
R15786 VSS.t32 VSS.n10978 25.542
R15787 VSS.t32 VSS.n10984 25.542
R15788 VSS.t32 VSS.n10985 25.542
R15789 VSS.t32 VSS.n10986 25.542
R15790 VSS.t32 VSS.n10987 25.542
R15791 VSS.t92 VSS.n10885 25.542
R15792 VSS.t92 VSS.n10886 25.542
R15793 VSS.t92 VSS.n10887 25.542
R15794 VSS.t92 VSS.n10888 25.542
R15795 VSS.t92 VSS.n10894 25.542
R15796 VSS.t92 VSS.n10895 25.542
R15797 VSS.t92 VSS.n10896 25.542
R15798 VSS.t92 VSS.n10897 25.542
R15799 VSS.t88 VSS.n10795 25.542
R15800 VSS.t88 VSS.n10796 25.542
R15801 VSS.t88 VSS.n10797 25.542
R15802 VSS.t88 VSS.n10798 25.542
R15803 VSS.t88 VSS.n10804 25.542
R15804 VSS.t88 VSS.n10805 25.542
R15805 VSS.t88 VSS.n10806 25.542
R15806 VSS.t88 VSS.n10807 25.542
R15807 VSS.t72 VSS.n10705 25.542
R15808 VSS.t72 VSS.n10706 25.542
R15809 VSS.t72 VSS.n10707 25.542
R15810 VSS.t72 VSS.n10708 25.542
R15811 VSS.t72 VSS.n10714 25.542
R15812 VSS.t72 VSS.n10715 25.542
R15813 VSS.t72 VSS.n10716 25.542
R15814 VSS.t72 VSS.n10717 25.542
R15815 VSS.t78 VSS.n10615 25.542
R15816 VSS.t78 VSS.n10616 25.542
R15817 VSS.t78 VSS.n10617 25.542
R15818 VSS.t78 VSS.n10618 25.542
R15819 VSS.t78 VSS.n10624 25.542
R15820 VSS.t78 VSS.n10625 25.542
R15821 VSS.t78 VSS.n10626 25.542
R15822 VSS.t78 VSS.n10627 25.542
R15823 VSS.t82 VSS.n10525 25.542
R15824 VSS.t82 VSS.n10526 25.542
R15825 VSS.t82 VSS.n10527 25.542
R15826 VSS.t82 VSS.n10528 25.542
R15827 VSS.t82 VSS.n10534 25.542
R15828 VSS.t82 VSS.n10535 25.542
R15829 VSS.t82 VSS.n10536 25.542
R15830 VSS.t82 VSS.n10537 25.542
R15831 VSS.t62 VSS.n13811 25.542
R15832 VSS.t62 VSS.n13812 25.542
R15833 VSS.t62 VSS.n13813 25.542
R15834 VSS.t62 VSS.n13814 25.542
R15835 VSS.t62 VSS.n13820 25.542
R15836 VSS.t62 VSS.n13821 25.542
R15837 VSS.t62 VSS.n13822 25.542
R15838 VSS.t62 VSS.n13884 25.542
R15839 VSS.t20 VSS.n9006 25.542
R15840 VSS.t20 VSS.n9004 25.542
R15841 VSS.t20 VSS.n9002 25.542
R15842 VSS.t20 VSS.n9000 25.542
R15843 VSS.t20 VSS.n9005 25.542
R15844 VSS.t20 VSS.n9003 25.542
R15845 VSS.t20 VSS.n9001 25.542
R15846 VSS.t20 VSS.n8999 25.542
R15847 VSS.t34 VSS.n9193 25.542
R15848 VSS.t34 VSS.n9194 25.542
R15849 VSS.t34 VSS.n9195 25.542
R15850 VSS.t34 VSS.n9196 25.542
R15851 VSS.t34 VSS.n9202 25.542
R15852 VSS.t34 VSS.n9203 25.542
R15853 VSS.t34 VSS.n9204 25.542
R15854 VSS.t34 VSS.n9205 25.542
R15855 VSS.t26 VSS.n9283 25.542
R15856 VSS.t26 VSS.n9284 25.542
R15857 VSS.t26 VSS.n9285 25.542
R15858 VSS.t26 VSS.n9286 25.542
R15859 VSS.t26 VSS.n9292 25.542
R15860 VSS.t26 VSS.n9293 25.542
R15861 VSS.t26 VSS.n9294 25.542
R15862 VSS.t26 VSS.n9295 25.542
R15863 VSS.t52 VSS.n9373 25.542
R15864 VSS.t52 VSS.n9374 25.542
R15865 VSS.t52 VSS.n9375 25.542
R15866 VSS.t52 VSS.n9376 25.542
R15867 VSS.t52 VSS.n9382 25.542
R15868 VSS.t52 VSS.n9383 25.542
R15869 VSS.t52 VSS.n9384 25.542
R15870 VSS.t52 VSS.n9385 25.542
R15871 VSS.t56 VSS.n9463 25.542
R15872 VSS.t56 VSS.n9464 25.542
R15873 VSS.t56 VSS.n9465 25.542
R15874 VSS.t56 VSS.n9466 25.542
R15875 VSS.t56 VSS.n9472 25.542
R15876 VSS.t56 VSS.n9473 25.542
R15877 VSS.t56 VSS.n9474 25.542
R15878 VSS.t56 VSS.n9475 25.542
R15879 VSS.t80 VSS.n9553 25.542
R15880 VSS.t80 VSS.n9554 25.542
R15881 VSS.t80 VSS.n9555 25.542
R15882 VSS.t80 VSS.n9556 25.542
R15883 VSS.t80 VSS.n9562 25.542
R15884 VSS.t80 VSS.n9563 25.542
R15885 VSS.t80 VSS.n9564 25.542
R15886 VSS.t80 VSS.n9565 25.542
R15887 VSS.t18 VSS.n9643 25.542
R15888 VSS.t18 VSS.n9644 25.542
R15889 VSS.t18 VSS.n9645 25.542
R15890 VSS.t18 VSS.n9646 25.542
R15891 VSS.t18 VSS.n9652 25.542
R15892 VSS.t18 VSS.n9653 25.542
R15893 VSS.t18 VSS.n9654 25.542
R15894 VSS.t18 VSS.n9655 25.542
R15895 VSS.n10324 VSS.t38 25.542
R15896 VSS.t38 VSS.n9176 25.542
R15897 VSS.t38 VSS.n9174 25.542
R15898 VSS.t38 VSS.n9172 25.542
R15899 VSS.t38 VSS.n9177 25.542
R15900 VSS.t38 VSS.n9175 25.542
R15901 VSS.t38 VSS.n9173 25.542
R15902 VSS.t38 VSS.n9171 25.542
R15903 VSS.t14 VSS.n6641 25.542
R15904 VSS.t14 VSS.n6651 25.542
R15905 VSS.t14 VSS.n6640 25.542
R15906 VSS.t14 VSS.n6639 25.542
R15907 VSS.t14 VSS.n6652 25.542
R15908 VSS.t14 VSS.n6653 25.542
R15909 VSS.t14 VSS.n6654 25.542
R15910 VSS.t14 VSS.n6637 25.542
R15911 VSS.t46 VSS.n5671 25.542
R15912 VSS.t46 VSS.n5672 25.542
R15913 VSS.t46 VSS.n5673 25.542
R15914 VSS.t46 VSS.n5674 25.542
R15915 VSS.t46 VSS.n5680 25.542
R15916 VSS.t46 VSS.n5681 25.542
R15917 VSS.t46 VSS.n5682 25.542
R15918 VSS.t46 VSS.n5732 25.542
R15919 VSS.t70 VSS.n5793 25.542
R15920 VSS.t70 VSS.n5794 25.542
R15921 VSS.t70 VSS.n5795 25.542
R15922 VSS.t70 VSS.n5796 25.542
R15923 VSS.t70 VSS.n5802 25.542
R15924 VSS.t70 VSS.n5803 25.542
R15925 VSS.t70 VSS.n5804 25.542
R15926 VSS.t70 VSS.n5854 25.542
R15927 VSS.t66 VSS.n5915 25.542
R15928 VSS.t66 VSS.n5916 25.542
R15929 VSS.t66 VSS.n5917 25.542
R15930 VSS.t66 VSS.n5918 25.542
R15931 VSS.t66 VSS.n5924 25.542
R15932 VSS.t66 VSS.n5925 25.542
R15933 VSS.t66 VSS.n5926 25.542
R15934 VSS.t66 VSS.n5976 25.542
R15935 VSS.t64 VSS.n6037 25.542
R15936 VSS.t64 VSS.n6038 25.542
R15937 VSS.t64 VSS.n6039 25.542
R15938 VSS.t64 VSS.n6040 25.542
R15939 VSS.t64 VSS.n6046 25.542
R15940 VSS.t64 VSS.n6047 25.542
R15941 VSS.t64 VSS.n6048 25.542
R15942 VSS.t64 VSS.n6098 25.542
R15943 VSS.t84 VSS.n6159 25.542
R15944 VSS.t84 VSS.n6160 25.542
R15945 VSS.t84 VSS.n6161 25.542
R15946 VSS.t84 VSS.n6162 25.542
R15947 VSS.t84 VSS.n6168 25.542
R15948 VSS.t84 VSS.n6169 25.542
R15949 VSS.t84 VSS.n6170 25.542
R15950 VSS.t84 VSS.n6220 25.542
R15951 VSS.t86 VSS.n6281 25.542
R15952 VSS.t86 VSS.n6282 25.542
R15953 VSS.t86 VSS.n6283 25.542
R15954 VSS.t86 VSS.n6284 25.542
R15955 VSS.t86 VSS.n6290 25.542
R15956 VSS.t86 VSS.n6291 25.542
R15957 VSS.t86 VSS.n6292 25.542
R15958 VSS.t86 VSS.n6342 25.542
R15959 VSS.t24 VSS.n6403 25.542
R15960 VSS.t24 VSS.n6404 25.542
R15961 VSS.t24 VSS.n6405 25.542
R15962 VSS.t24 VSS.n6406 25.542
R15963 VSS.t24 VSS.n6412 25.542
R15964 VSS.t24 VSS.n6413 25.542
R15965 VSS.t24 VSS.n6414 25.542
R15966 VSS.t24 VSS.n6464 25.542
R15967 VSS.n6586 VSS.t44 25.542
R15968 VSS.n6521 VSS.t44 25.542
R15969 VSS.n6579 VSS.t44 25.542
R15970 VSS.n6524 VSS.t44 25.542
R15971 VSS.n6555 VSS.t44 25.542
R15972 VSS.n6549 VSS.t44 25.542
R15973 VSS.n6547 VSS.t44 25.542
R15974 VSS.n6541 VSS.t44 25.542
R15975 VSS.t60 VSS.n10 25.542
R15976 VSS.t60 VSS.n11 25.542
R15977 VSS.t60 VSS.n12 25.542
R15978 VSS.t60 VSS.n13 25.542
R15979 VSS.t60 VSS.n19 25.542
R15980 VSS.t60 VSS.n20 25.542
R15981 VSS.t60 VSS.n21 25.542
R15982 VSS.t60 VSS.n22 25.542
R15983 VSS.t48 VSS.n101 25.542
R15984 VSS.t48 VSS.n102 25.542
R15985 VSS.t48 VSS.n103 25.542
R15986 VSS.t48 VSS.n104 25.542
R15987 VSS.t48 VSS.n110 25.542
R15988 VSS.t48 VSS.n111 25.542
R15989 VSS.t48 VSS.n112 25.542
R15990 VSS.t48 VSS.n113 25.542
R15991 VSS.t76 VSS.n191 25.542
R15992 VSS.t76 VSS.n192 25.542
R15993 VSS.t76 VSS.n193 25.542
R15994 VSS.t76 VSS.n194 25.542
R15995 VSS.t76 VSS.n200 25.542
R15996 VSS.t76 VSS.n201 25.542
R15997 VSS.t76 VSS.n202 25.542
R15998 VSS.t76 VSS.n203 25.542
R15999 VSS.t22 VSS.n281 25.542
R16000 VSS.t22 VSS.n282 25.542
R16001 VSS.t22 VSS.n283 25.542
R16002 VSS.t22 VSS.n284 25.542
R16003 VSS.t22 VSS.n290 25.542
R16004 VSS.t22 VSS.n291 25.542
R16005 VSS.t22 VSS.n292 25.542
R16006 VSS.t22 VSS.n293 25.542
R16007 VSS.t16 VSS.n371 25.542
R16008 VSS.t16 VSS.n372 25.542
R16009 VSS.t16 VSS.n373 25.542
R16010 VSS.t16 VSS.n374 25.542
R16011 VSS.t16 VSS.n380 25.542
R16012 VSS.t16 VSS.n381 25.542
R16013 VSS.t16 VSS.n382 25.542
R16014 VSS.t16 VSS.n383 25.542
R16015 VSS.t36 VSS.n461 25.542
R16016 VSS.t36 VSS.n462 25.542
R16017 VSS.t36 VSS.n463 25.542
R16018 VSS.t36 VSS.n464 25.542
R16019 VSS.t36 VSS.n470 25.542
R16020 VSS.t36 VSS.n471 25.542
R16021 VSS.t36 VSS.n472 25.542
R16022 VSS.t36 VSS.n473 25.542
R16023 VSS.t40 VSS.n551 25.542
R16024 VSS.t40 VSS.n552 25.542
R16025 VSS.t40 VSS.n553 25.542
R16026 VSS.t40 VSS.n554 25.542
R16027 VSS.t40 VSS.n560 25.542
R16028 VSS.t40 VSS.n561 25.542
R16029 VSS.t40 VSS.n562 25.542
R16030 VSS.t40 VSS.n563 25.542
R16031 VSS.n6711 VSS.n6708 23.644
R16032 VSS.t14 VSS.n6650 19.67
R16033 VSS.n14719 VSS.n14366 19.504
R16034 VSS.n14715 VSS.n14372 19.504
R16035 VSS.n14703 VSS.n14380 19.504
R16036 VSS.n14696 VSS.n14388 19.504
R16037 VSS.n14692 VSS.n14392 19.504
R16038 VSS.n14680 VSS.n14399 19.504
R16039 VSS.n14674 VSS.n14407 19.504
R16040 VSS.n14670 VSS.n14411 19.504
R16041 VSS.n14658 VSS.n14418 19.504
R16042 VSS.n14651 VSS.n14426 19.504
R16043 VSS.n14647 VSS.n14430 19.504
R16044 VSS.n14635 VSS.n14437 19.504
R16045 VSS.n14876 VSS.n14296 19.504
R16046 VSS.n14888 VSS.n14294 19.504
R16047 VSS.n14896 VSS.n14287 19.504
R16048 VSS.n14907 VSS.n14281 19.504
R16049 VSS.n14911 VSS.n14275 19.504
R16050 VSS.n14923 VSS.n14273 19.504
R16051 VSS.n14930 VSS.n14266 19.504
R16052 VSS.n14941 VSS.n14260 19.504
R16053 VSS.n14945 VSS.n14254 19.504
R16054 VSS.n14957 VSS.n14252 19.504
R16055 VSS.n14965 VSS.n14245 19.504
R16056 VSS.n15329 VSS.n14240 19.504
R16057 VSS.n14627 VSS.n14478 19.504
R16058 VSS.n14623 VSS.n14485 19.504
R16059 VSS.n14611 VSS.n14492 19.504
R16060 VSS.n14604 VSS.n14500 19.504
R16061 VSS.n14600 VSS.n14504 19.504
R16062 VSS.n14588 VSS.n14511 19.504
R16063 VSS.n14582 VSS.n14519 19.504
R16064 VSS.n14578 VSS.n14523 19.504
R16065 VSS.n14566 VSS.n14530 19.504
R16066 VSS.n14559 VSS.n14538 19.504
R16067 VSS.n14555 VSS.n14542 19.504
R16068 VSS.n14871 VSS.n14303 19.504
R16069 VSS.n15228 VSS.n15087 19.504
R16070 VSS.n15224 VSS.n15094 19.504
R16071 VSS.n15212 VSS.n15101 19.504
R16072 VSS.n15205 VSS.n15109 19.504
R16073 VSS.n15201 VSS.n15113 19.504
R16074 VSS.n15189 VSS.n15120 19.504
R16075 VSS.n15183 VSS.n15128 19.504
R16076 VSS.n15179 VSS.n15132 19.504
R16077 VSS.n15167 VSS.n15139 19.504
R16078 VSS.n15160 VSS.n15147 19.504
R16079 VSS.n15156 VSS.n14141 19.504
R16080 VSS.n15442 VSS.n14142 19.504
R16081 VSS.n15320 VSS.n14978 19.504
R16082 VSS.n15316 VSS.n14982 19.504
R16083 VSS.n15304 VSS.n14989 19.504
R16084 VSS.n15297 VSS.n14997 19.504
R16085 VSS.n15293 VSS.n15001 19.504
R16086 VSS.n15281 VSS.n15008 19.504
R16087 VSS.n15275 VSS.n15016 19.504
R16088 VSS.n15271 VSS.n15020 19.504
R16089 VSS.n15259 VSS.n15027 19.504
R16090 VSS.n15252 VSS.n15035 19.504
R16091 VSS.n15248 VSS.n15039 19.504
R16092 VSS.n15236 VSS.n15046 19.504
R16093 VSS.n15887 VSS.n15563 19.504
R16094 VSS.n15883 VSS.n15569 19.504
R16095 VSS.n15871 VSS.n15576 19.504
R16096 VSS.n15864 VSS.n15584 19.504
R16097 VSS.n15860 VSS.n15588 19.504
R16098 VSS.n15848 VSS.n15595 19.504
R16099 VSS.n15842 VSS.n15603 19.504
R16100 VSS.n15838 VSS.n15607 19.504
R16101 VSS.n15826 VSS.n15614 19.504
R16102 VSS.n15819 VSS.n15622 19.504
R16103 VSS.n15815 VSS.n15626 19.504
R16104 VSS.n15803 VSS.n15633 19.504
R16105 VSS.n15459 VSS.n14131 19.504
R16106 VSS.n15470 VSS.n14125 19.504
R16107 VSS.n15474 VSS.n14119 19.504
R16108 VSS.n15486 VSS.n14117 19.504
R16109 VSS.n15494 VSS.n14110 19.504
R16110 VSS.n15505 VSS.n14104 19.504
R16111 VSS.n15509 VSS.n14098 19.504
R16112 VSS.n15520 VSS.n14096 19.504
R16113 VSS.n15528 VSS.n14089 19.504
R16114 VSS.n15539 VSS.n14083 19.504
R16115 VSS.n15543 VSS.n14077 19.504
R16116 VSS.n15555 VSS.n14075 19.504
R16117 VSS.n15795 VSS.n15674 19.504
R16118 VSS.n15791 VSS.n15681 19.504
R16119 VSS.n15779 VSS.n15688 19.504
R16120 VSS.n15772 VSS.n15696 19.504
R16121 VSS.n15768 VSS.n15700 19.504
R16122 VSS.n15756 VSS.n15707 19.504
R16123 VSS.n15750 VSS.n15715 19.504
R16124 VSS.n15746 VSS.n15719 19.504
R16125 VSS.n15734 VSS.n15726 19.504
R16126 VSS.n16020 VSS.n13999 19.504
R16127 VSS.n16016 VSS.n14003 19.504
R16128 VSS.n16004 VSS.n14010 19.504
R16129 VSS.n12798 VSS.n12721 19.504
R16130 VSS.n12806 VSS.n12714 19.504
R16131 VSS.n12817 VSS.n12708 19.504
R16132 VSS.n12821 VSS.n12702 19.504
R16133 VSS.n12833 VSS.n12700 19.504
R16134 VSS.n12841 VSS.n12693 19.504
R16135 VSS.n12851 VSS.n12687 19.504
R16136 VSS.n12855 VSS.n12681 19.504
R16137 VSS.n12867 VSS.n12679 19.504
R16138 VSS.n12875 VSS.n12671 19.504
R16139 VSS.n12672 VSS.n12666 19.504
R16140 VSS.n13059 VSS.n12663 19.504
R16141 VSS.n13155 VSS.n12580 19.504
R16142 VSS.n13163 VSS.n12573 19.504
R16143 VSS.n13174 VSS.n12567 19.504
R16144 VSS.n13178 VSS.n12561 19.504
R16145 VSS.n13190 VSS.n12559 19.504
R16146 VSS.n13198 VSS.n12552 19.504
R16147 VSS.n13208 VSS.n12546 19.504
R16148 VSS.n13212 VSS.n12540 19.504
R16149 VSS.n13224 VSS.n12538 19.504
R16150 VSS.n13232 VSS.n12530 19.504
R16151 VSS.n12531 VSS.n12525 19.504
R16152 VSS.n13308 VSS.n12522 19.504
R16153 VSS.n13054 VSS.n12893 19.504
R16154 VSS.n13042 VSS.n12897 19.504
R16155 VSS.n13035 VSS.n12906 19.504
R16156 VSS.n13031 VSS.n12910 19.504
R16157 VSS.n13019 VSS.n12917 19.504
R16158 VSS.n13012 VSS.n12925 19.504
R16159 VSS.n13008 VSS.n12929 19.504
R16160 VSS.n12997 VSS.n12936 19.504
R16161 VSS.n12990 VSS.n12944 19.504
R16162 VSS.n12986 VSS.n12948 19.504
R16163 VSS.n12974 VSS.n12955 19.504
R16164 VSS.n12967 VSS.n12964 19.504
R16165 VSS.n11676 VSS.n11671 19.504
R16166 VSS.n11684 VSS.n11664 19.504
R16167 VSS.n11695 VSS.n11658 19.504
R16168 VSS.n11699 VSS.n11652 19.504
R16169 VSS.n11711 VSS.n11650 19.504
R16170 VSS.n11719 VSS.n11643 19.504
R16171 VSS.n11729 VSS.n11637 19.504
R16172 VSS.n11733 VSS.n11631 19.504
R16173 VSS.n11745 VSS.n11629 19.504
R16174 VSS.n11753 VSS.n11622 19.504
R16175 VSS.n11764 VSS.n11615 19.504
R16176 VSS.n11769 VSS.n11768 19.504
R16177 VSS.n13303 VSS.n13250 19.504
R16178 VSS.n13291 VSS.n13254 19.504
R16179 VSS.n13284 VSS.n13263 19.504
R16180 VSS.n13280 VSS.n13267 19.504
R16181 VSS.n13454 VSS.n11433 19.504
R16182 VSS.n13450 VSS.n11437 19.504
R16183 VSS.n13438 VSS.n11444 19.504
R16184 VSS.n13432 VSS.n11452 19.504
R16185 VSS.n13428 VSS.n11456 19.504
R16186 VSS.n13416 VSS.n11463 19.504
R16187 VSS.n13409 VSS.n11471 19.504
R16188 VSS.n13405 VSS.n11475 19.504
R16189 VSS.n12395 VSS.n11912 19.504
R16190 VSS.n12391 VSS.n11916 19.504
R16191 VSS.n12379 VSS.n11923 19.504
R16192 VSS.n12372 VSS.n11931 19.504
R16193 VSS.n12368 VSS.n11935 19.504
R16194 VSS.n12356 VSS.n11942 19.504
R16195 VSS.n12350 VSS.n11950 19.504
R16196 VSS.n12346 VSS.n11954 19.504
R16197 VSS.n12334 VSS.n11961 19.504
R16198 VSS.n12327 VSS.n11969 19.504
R16199 VSS.n12323 VSS.n11973 19.504
R16200 VSS.n12311 VSS.n11980 19.504
R16201 VSS.n11810 VSS.n11601 19.504
R16202 VSS.n11822 VSS.n11599 19.504
R16203 VSS.n11830 VSS.n11592 19.504
R16204 VSS.n11841 VSS.n11586 19.504
R16205 VSS.n11845 VSS.n11580 19.504
R16206 VSS.n11857 VSS.n11578 19.504
R16207 VSS.n11864 VSS.n11571 19.504
R16208 VSS.n11875 VSS.n11565 19.504
R16209 VSS.n11879 VSS.n11559 19.504
R16210 VSS.n11891 VSS.n11557 19.504
R16211 VSS.n11899 VSS.n11550 19.504
R16212 VSS.n12404 VSS.n11545 19.504
R16213 VSS.n12303 VSS.n11988 19.504
R16214 VSS.n12299 VSS.n11995 19.504
R16215 VSS.n12287 VSS.n12002 19.504
R16216 VSS.n12280 VSS.n12010 19.504
R16217 VSS.n12276 VSS.n12014 19.504
R16218 VSS.n12264 VSS.n12021 19.504
R16219 VSS.n12258 VSS.n12029 19.504
R16220 VSS.n12254 VSS.n12033 19.504
R16221 VSS.n12242 VSS.n12040 19.504
R16222 VSS.n12235 VSS.n12048 19.504
R16223 VSS.n12231 VSS.n12052 19.504
R16224 VSS.n12219 VSS.n12059 19.504
R16225 VSS.n7833 VSS.n7674 19.504
R16226 VSS.n7829 VSS.n7679 19.504
R16227 VSS.n7817 VSS.n7687 19.504
R16228 VSS.n7810 VSS.n7695 19.504
R16229 VSS.n7806 VSS.n7699 19.504
R16230 VSS.n7794 VSS.n7706 19.504
R16231 VSS.n7788 VSS.n7714 19.504
R16232 VSS.n7784 VSS.n7718 19.504
R16233 VSS.n7772 VSS.n7725 19.504
R16234 VSS.n7765 VSS.n7733 19.504
R16235 VSS.n7761 VSS.n7737 19.504
R16236 VSS.n7750 VSS.n7749 19.504
R16237 VSS.n8181 VSS.n8020 19.504
R16238 VSS.n8173 VSS.n8022 19.504
R16239 VSS.n8169 VSS.n8033 19.504
R16240 VSS.n8157 VSS.n8041 19.504
R16241 VSS.n8150 VSS.n8049 19.504
R16242 VSS.n8146 VSS.n8053 19.504
R16243 VSS.n8134 VSS.n8060 19.504
R16244 VSS.n8128 VSS.n8068 19.504
R16245 VSS.n8124 VSS.n8072 19.504
R16246 VSS.n8112 VSS.n8079 19.504
R16247 VSS.n8105 VSS.n8087 19.504
R16248 VSS.n8101 VSS.n8090 19.504
R16249 VSS.n7921 VSS.n7595 19.504
R16250 VSS.n7933 VSS.n7593 19.504
R16251 VSS.n7941 VSS.n7586 19.504
R16252 VSS.n7952 VSS.n7580 19.504
R16253 VSS.n7956 VSS.n7574 19.504
R16254 VSS.n7968 VSS.n7572 19.504
R16255 VSS.n7975 VSS.n7565 19.504
R16256 VSS.n7986 VSS.n7559 19.504
R16257 VSS.n7990 VSS.n7553 19.504
R16258 VSS.n8002 VSS.n7551 19.504
R16259 VSS.n8010 VSS.n7544 19.504
R16260 VSS.n8190 VSS.n7538 19.504
R16261 VSS.n8539 VSS.n8378 19.504
R16262 VSS.n8531 VSS.n8380 19.504
R16263 VSS.n8527 VSS.n8391 19.504
R16264 VSS.n8515 VSS.n8399 19.504
R16265 VSS.n8508 VSS.n8407 19.504
R16266 VSS.n8504 VSS.n8411 19.504
R16267 VSS.n8492 VSS.n8418 19.504
R16268 VSS.n8486 VSS.n8426 19.504
R16269 VSS.n8482 VSS.n8430 19.504
R16270 VSS.n8470 VSS.n8437 19.504
R16271 VSS.n8463 VSS.n8445 19.504
R16272 VSS.n8459 VSS.n8448 19.504
R16273 VSS.n8279 VSS.n7455 19.504
R16274 VSS.n8291 VSS.n7453 19.504
R16275 VSS.n8299 VSS.n7446 19.504
R16276 VSS.n8310 VSS.n7440 19.504
R16277 VSS.n8314 VSS.n7434 19.504
R16278 VSS.n8326 VSS.n7432 19.504
R16279 VSS.n8333 VSS.n7425 19.504
R16280 VSS.n8344 VSS.n7419 19.504
R16281 VSS.n8348 VSS.n7413 19.504
R16282 VSS.n8360 VSS.n7411 19.504
R16283 VSS.n8368 VSS.n7404 19.504
R16284 VSS.n8548 VSS.n7398 19.504
R16285 VSS.n8761 VSS.n8736 19.504
R16286 VSS.n8753 VSS.n8738 19.504
R16287 VSS.n8926 VSS.n6905 19.504
R16288 VSS.n8922 VSS.n6909 19.504
R16289 VSS.n8910 VSS.n6916 19.504
R16290 VSS.n8903 VSS.n6924 19.504
R16291 VSS.n8899 VSS.n6928 19.504
R16292 VSS.n8888 VSS.n6935 19.504
R16293 VSS.n8881 VSS.n6943 19.504
R16294 VSS.n8877 VSS.n6947 19.504
R16295 VSS.n8865 VSS.n6954 19.504
R16296 VSS.n8858 VSS.n6962 19.504
R16297 VSS.n8637 VSS.n7315 19.504
R16298 VSS.n8649 VSS.n7313 19.504
R16299 VSS.n8657 VSS.n7306 19.504
R16300 VSS.n8668 VSS.n7300 19.504
R16301 VSS.n8672 VSS.n7294 19.504
R16302 VSS.n8684 VSS.n7292 19.504
R16303 VSS.n8691 VSS.n7285 19.504
R16304 VSS.n8702 VSS.n7279 19.504
R16305 VSS.n8706 VSS.n7273 19.504
R16306 VSS.n8718 VSS.n7271 19.504
R16307 VSS.n8726 VSS.n7264 19.504
R16308 VSS.n8770 VSS.n7258 19.504
R16309 VSS.n7075 VSS.n7066 19.504
R16310 VSS.n7086 VSS.n7060 19.504
R16311 VSS.n7090 VSS.n7054 19.504
R16312 VSS.n7102 VSS.n7052 19.504
R16313 VSS.n7110 VSS.n7045 19.504
R16314 VSS.n7121 VSS.n7039 19.504
R16315 VSS.n7125 VSS.n7033 19.504
R16316 VSS.n7136 VSS.n7031 19.504
R16317 VSS.n7144 VSS.n7024 19.504
R16318 VSS.n7155 VSS.n7018 19.504
R16319 VSS.n7159 VSS.n7012 19.504
R16320 VSS.n7172 VSS.n7009 19.504
R16321 VSS.n4251 VSS.n4174 19.504
R16322 VSS.n4259 VSS.n4167 19.504
R16323 VSS.n4270 VSS.n4161 19.504
R16324 VSS.n4274 VSS.n4155 19.504
R16325 VSS.n4286 VSS.n4153 19.504
R16326 VSS.n4294 VSS.n4146 19.504
R16327 VSS.n4304 VSS.n4140 19.504
R16328 VSS.n4308 VSS.n4134 19.504
R16329 VSS.n4320 VSS.n4132 19.504
R16330 VSS.n4328 VSS.n4124 19.504
R16331 VSS.n4125 VSS.n4119 19.504
R16332 VSS.n4512 VSS.n4116 19.504
R16333 VSS.n4608 VSS.n4033 19.504
R16334 VSS.n4616 VSS.n4026 19.504
R16335 VSS.n4627 VSS.n4020 19.504
R16336 VSS.n4631 VSS.n4014 19.504
R16337 VSS.n4643 VSS.n4012 19.504
R16338 VSS.n4651 VSS.n4005 19.504
R16339 VSS.n4661 VSS.n3999 19.504
R16340 VSS.n4665 VSS.n3993 19.504
R16341 VSS.n4677 VSS.n3991 19.504
R16342 VSS.n4685 VSS.n3983 19.504
R16343 VSS.n3984 VSS.n3978 19.504
R16344 VSS.n4869 VSS.n3975 19.504
R16345 VSS.n4507 VSS.n4346 19.504
R16346 VSS.n4495 VSS.n4350 19.504
R16347 VSS.n4488 VSS.n4359 19.504
R16348 VSS.n4484 VSS.n4363 19.504
R16349 VSS.n4472 VSS.n4370 19.504
R16350 VSS.n4465 VSS.n4378 19.504
R16351 VSS.n4461 VSS.n4382 19.504
R16352 VSS.n4450 VSS.n4389 19.504
R16353 VSS.n4443 VSS.n4397 19.504
R16354 VSS.n4439 VSS.n4401 19.504
R16355 VSS.n4427 VSS.n4408 19.504
R16356 VSS.n4420 VSS.n4417 19.504
R16357 VSS.n4965 VSS.n3892 19.504
R16358 VSS.n4973 VSS.n3885 19.504
R16359 VSS.n4984 VSS.n3879 19.504
R16360 VSS.n4988 VSS.n3873 19.504
R16361 VSS.n5000 VSS.n3871 19.504
R16362 VSS.n5008 VSS.n3864 19.504
R16363 VSS.n5018 VSS.n3858 19.504
R16364 VSS.n5022 VSS.n3852 19.504
R16365 VSS.n5034 VSS.n3850 19.504
R16366 VSS.n5042 VSS.n3842 19.504
R16367 VSS.n3843 VSS.n3837 19.504
R16368 VSS.n5226 VSS.n3834 19.504
R16369 VSS.n4864 VSS.n4703 19.504
R16370 VSS.n4852 VSS.n4707 19.504
R16371 VSS.n4845 VSS.n4716 19.504
R16372 VSS.n4841 VSS.n4720 19.504
R16373 VSS.n4829 VSS.n4727 19.504
R16374 VSS.n4822 VSS.n4735 19.504
R16375 VSS.n4818 VSS.n4739 19.504
R16376 VSS.n4807 VSS.n4746 19.504
R16377 VSS.n4800 VSS.n4754 19.504
R16378 VSS.n4796 VSS.n4758 19.504
R16379 VSS.n4784 VSS.n4765 19.504
R16380 VSS.n4777 VSS.n4774 19.504
R16381 VSS.n5322 VSS.n3751 19.504
R16382 VSS.n5330 VSS.n3744 19.504
R16383 VSS.n5341 VSS.n3738 19.504
R16384 VSS.n5345 VSS.n3732 19.504
R16385 VSS.n5357 VSS.n3730 19.504
R16386 VSS.n5365 VSS.n3723 19.504
R16387 VSS.n5375 VSS.n3717 19.504
R16388 VSS.n5379 VSS.n3711 19.504
R16389 VSS.n5391 VSS.n3709 19.504
R16390 VSS.n5399 VSS.n3701 19.504
R16391 VSS.n3702 VSS.n3696 19.504
R16392 VSS.n5572 VSS.n3693 19.504
R16393 VSS.n5221 VSS.n5060 19.504
R16394 VSS.n5209 VSS.n5064 19.504
R16395 VSS.n5202 VSS.n5073 19.504
R16396 VSS.n5198 VSS.n5077 19.504
R16397 VSS.n5186 VSS.n5084 19.504
R16398 VSS.n5179 VSS.n5092 19.504
R16399 VSS.n5175 VSS.n5096 19.504
R16400 VSS.n5164 VSS.n5103 19.504
R16401 VSS.n5157 VSS.n5111 19.504
R16402 VSS.n5153 VSS.n5115 19.504
R16403 VSS.n5141 VSS.n5122 19.504
R16404 VSS.n5134 VSS.n5131 19.504
R16405 VSS.n5567 VSS.n5417 19.504
R16406 VSS.n5555 VSS.n5421 19.504
R16407 VSS.n5548 VSS.n5430 19.504
R16408 VSS.n5544 VSS.n5434 19.504
R16409 VSS.n5532 VSS.n5441 19.504
R16410 VSS.n5525 VSS.n5449 19.504
R16411 VSS.n5521 VSS.n5453 19.504
R16412 VSS.n5510 VSS.n5460 19.504
R16413 VSS.n5503 VSS.n5468 19.504
R16414 VSS.n5499 VSS.n5472 19.504
R16415 VSS.n5487 VSS.n5479 19.504
R16416 VSS.n5660 VSS.n3639 19.504
R16417 VSS.n1960 VSS.n1607 19.504
R16418 VSS.n1956 VSS.n1613 19.504
R16419 VSS.n1944 VSS.n1621 19.504
R16420 VSS.n1937 VSS.n1629 19.504
R16421 VSS.n1933 VSS.n1633 19.504
R16422 VSS.n1921 VSS.n1640 19.504
R16423 VSS.n1915 VSS.n1648 19.504
R16424 VSS.n1911 VSS.n1652 19.504
R16425 VSS.n1899 VSS.n1659 19.504
R16426 VSS.n1892 VSS.n1667 19.504
R16427 VSS.n1888 VSS.n1671 19.504
R16428 VSS.n1876 VSS.n1678 19.504
R16429 VSS.n2117 VSS.n1537 19.504
R16430 VSS.n2129 VSS.n1535 19.504
R16431 VSS.n2137 VSS.n1528 19.504
R16432 VSS.n2148 VSS.n1522 19.504
R16433 VSS.n2152 VSS.n1516 19.504
R16434 VSS.n2164 VSS.n1514 19.504
R16435 VSS.n2171 VSS.n1507 19.504
R16436 VSS.n2182 VSS.n1501 19.504
R16437 VSS.n2186 VSS.n1495 19.504
R16438 VSS.n2198 VSS.n1493 19.504
R16439 VSS.n2206 VSS.n1486 19.504
R16440 VSS.n2570 VSS.n1481 19.504
R16441 VSS.n1868 VSS.n1719 19.504
R16442 VSS.n1864 VSS.n1726 19.504
R16443 VSS.n1852 VSS.n1733 19.504
R16444 VSS.n1845 VSS.n1741 19.504
R16445 VSS.n1841 VSS.n1745 19.504
R16446 VSS.n1829 VSS.n1752 19.504
R16447 VSS.n1823 VSS.n1760 19.504
R16448 VSS.n1819 VSS.n1764 19.504
R16449 VSS.n1807 VSS.n1771 19.504
R16450 VSS.n1800 VSS.n1779 19.504
R16451 VSS.n1796 VSS.n1783 19.504
R16452 VSS.n2112 VSS.n1544 19.504
R16453 VSS.n2469 VSS.n2328 19.504
R16454 VSS.n2465 VSS.n2335 19.504
R16455 VSS.n2453 VSS.n2342 19.504
R16456 VSS.n2446 VSS.n2350 19.504
R16457 VSS.n2442 VSS.n2354 19.504
R16458 VSS.n2430 VSS.n2361 19.504
R16459 VSS.n2424 VSS.n2369 19.504
R16460 VSS.n2420 VSS.n2373 19.504
R16461 VSS.n2408 VSS.n2380 19.504
R16462 VSS.n2401 VSS.n2388 19.504
R16463 VSS.n2397 VSS.n1382 19.504
R16464 VSS.n2683 VSS.n1383 19.504
R16465 VSS.n2561 VSS.n2219 19.504
R16466 VSS.n2557 VSS.n2223 19.504
R16467 VSS.n2545 VSS.n2230 19.504
R16468 VSS.n2538 VSS.n2238 19.504
R16469 VSS.n2534 VSS.n2242 19.504
R16470 VSS.n2522 VSS.n2249 19.504
R16471 VSS.n2516 VSS.n2257 19.504
R16472 VSS.n2512 VSS.n2261 19.504
R16473 VSS.n2500 VSS.n2268 19.504
R16474 VSS.n2493 VSS.n2276 19.504
R16475 VSS.n2489 VSS.n2280 19.504
R16476 VSS.n2477 VSS.n2287 19.504
R16477 VSS.n2700 VSS.n1372 19.504
R16478 VSS.n2711 VSS.n1366 19.504
R16479 VSS.n2715 VSS.n1360 19.504
R16480 VSS.n2727 VSS.n1358 19.504
R16481 VSS.n2735 VSS.n1351 19.504
R16482 VSS.n2746 VSS.n1345 19.504
R16483 VSS.n2750 VSS.n1339 19.504
R16484 VSS.n2761 VSS.n1337 19.504
R16485 VSS.n2769 VSS.n1330 19.504
R16486 VSS.n2780 VSS.n1324 19.504
R16487 VSS.n2784 VSS.n1318 19.504
R16488 VSS.n2796 VSS.n1316 19.504
R16489 VSS.n2961 VSS.n2804 19.504
R16490 VSS.n2957 VSS.n2810 19.504
R16491 VSS.n2945 VSS.n2817 19.504
R16492 VSS.n2938 VSS.n2825 19.504
R16493 VSS.n2934 VSS.n2829 19.504
R16494 VSS.n2922 VSS.n2836 19.504
R16495 VSS.n2916 VSS.n2844 19.504
R16496 VSS.n2912 VSS.n2848 19.504
R16497 VSS.n2900 VSS.n2855 19.504
R16498 VSS.n2893 VSS.n2863 19.504
R16499 VSS.n2889 VSS.n2867 19.504
R16500 VSS.n2878 VSS.n1270 19.504
R16501 VSS.n17686 VSS.n17685 19.393
R16502 VSS.n10444 VSS.n10429 19.392
R16503 VSS.n10469 VSS.n10424 19.392
R16504 VSS.n17672 VSS.n17651 19.392
R16505 VSS.n17692 VSS.n17691 19.349
R16506 VSS.n10449 VSS.n10430 19.349
R16507 VSS.n10474 VSS.n10422 19.349
R16508 VSS.n17670 VSS.n17653 19.349
R16509 VSS.n17696 VSS.n17695 19.301
R16510 VSS.t20 VSS.n8997 19.3
R16511 VSS.t38 VSS.n9169 19.3
R16512 VSS.n10454 VSS.n10431 19.3
R16513 VSS.n10479 VSS.n10420 19.3
R16514 VSS.n17665 VSS.n17655 19.3
R16515 VSS.n10461 VSS.n10460 19.247
R16516 VSS.n10484 VSS.n10418 19.247
R16517 VSS.n17660 VSS.n17657 19.247
R16518 VSS.n17702 VSS.n17701 19.247
R16519 VSS.n14472 VSS.n14439 18.614
R16520 VSS.n14863 VSS.n14304 18.614
R16521 VSS.n15333 VSS.n14237 18.614
R16522 VSS.n15081 VSS.n15048 18.614
R16523 VSS.n15441 VSS.n15440 18.614
R16524 VSS.n15893 VSS.n14070 18.614
R16525 VSS.n15668 VSS.n15635 18.614
R16526 VSS.n12664 VSS.n12657 18.614
R16527 VSS.n13147 VSS.n12582 18.614
R16528 VSS.n12523 VSS.n12516 18.614
R16529 VSS.n13396 VSS.n11483 18.614
R16530 VSS.n11805 VSS.n11608 18.614
R16531 VSS.n12408 VSS.n11542 18.614
R16532 VSS.n12103 VSS.n11982 18.614
R16533 VSS.n7916 VSS.n7602 18.614
R16534 VSS.n7539 VSS.n7535 18.614
R16535 VSS.n8274 VSS.n7462 18.614
R16536 VSS.n7399 VSS.n7395 18.614
R16537 VSS.n8632 VSS.n7322 18.614
R16538 VSS.n7259 VSS.n7255 18.614
R16539 VSS.n8854 VSS.n6963 18.614
R16540 VSS.n4117 VSS.n4110 18.614
R16541 VSS.n4600 VSS.n4035 18.614
R16542 VSS.n3976 VSS.n3969 18.614
R16543 VSS.n4957 VSS.n3894 18.614
R16544 VSS.n3835 VSS.n3828 18.614
R16545 VSS.n5314 VSS.n3753 18.614
R16546 VSS.n3694 VSS.n3687 18.614
R16547 VSS.n1713 VSS.n1680 18.614
R16548 VSS.n2104 VSS.n1545 18.614
R16549 VSS.n2574 VSS.n1478 18.614
R16550 VSS.n2322 VSS.n2289 18.614
R16551 VSS.n2682 VSS.n2681 18.614
R16552 VSS.n2967 VSS.n1311 18.614
R16553 VSS.n14752 VSS.n14350 17.453
R16554 VSS.n12766 VSS.n12765 17.453
R16555 VSS.n7866 VSS.n7865 17.453
R16556 VSS.n6855 VSS.n6744 17.453
R16557 VSS.n4219 VSS.n4218 17.453
R16558 VSS.n1993 VSS.n1591 17.453
R16559 VSS.n6692 VSS.n6691 17.422
R16560 VSS.n15974 VSS.n15973 17.065
R16561 VSS.n12189 VSS.n12188 17.065
R16562 VSS.n7203 VSS.n7202 17.065
R16563 VSS.n5631 VSS.n3657 17.065
R16564 VSS.n3020 VSS.n1283 17.065
R16565 VSS.n17386 VSS.n17385 16.666
R16566 VSS.n16047 VSS.n16034 16.666
R16567 VSS.n17454 VSS.n16037 16.666
R16568 VSS.n17445 VSS.n16033 16.666
R16569 VSS.n17439 VSS.n16038 16.666
R16570 VSS.n17433 VSS.n16032 16.666
R16571 VSS.n17427 VSS.n16039 16.666
R16572 VSS.n17421 VSS.n16031 16.666
R16573 VSS.n17461 VSS.n16029 16.666
R16574 VSS.n17224 VSS.n16090 16.666
R16575 VSS.n17298 VSS.n16076 16.666
R16576 VSS.n17289 VSS.n16073 16.666
R16577 VSS.n17283 VSS.n16077 16.666
R16578 VSS.n17277 VSS.n16072 16.666
R16579 VSS.n17271 VSS.n16078 16.666
R16580 VSS.n17265 VSS.n16071 16.666
R16581 VSS.n17306 VSS.n16080 16.666
R16582 VSS.n17134 VSS.n16180 16.666
R16583 VSS.n17208 VSS.n16166 16.666
R16584 VSS.n17199 VSS.n16163 16.666
R16585 VSS.n17193 VSS.n16167 16.666
R16586 VSS.n17187 VSS.n16162 16.666
R16587 VSS.n17181 VSS.n16168 16.666
R16588 VSS.n17175 VSS.n16161 16.666
R16589 VSS.n17216 VSS.n16170 16.666
R16590 VSS.n17044 VSS.n16270 16.666
R16591 VSS.n17118 VSS.n16256 16.666
R16592 VSS.n17109 VSS.n16253 16.666
R16593 VSS.n17103 VSS.n16257 16.666
R16594 VSS.n17097 VSS.n16252 16.666
R16595 VSS.n17091 VSS.n16258 16.666
R16596 VSS.n17085 VSS.n16251 16.666
R16597 VSS.n17126 VSS.n16260 16.666
R16598 VSS.n16954 VSS.n16360 16.666
R16599 VSS.n17028 VSS.n16346 16.666
R16600 VSS.n17019 VSS.n16343 16.666
R16601 VSS.n17013 VSS.n16347 16.666
R16602 VSS.n17007 VSS.n16342 16.666
R16603 VSS.n17001 VSS.n16348 16.666
R16604 VSS.n16995 VSS.n16341 16.666
R16605 VSS.n17036 VSS.n16350 16.666
R16606 VSS.n16864 VSS.n16450 16.666
R16607 VSS.n16938 VSS.n16436 16.666
R16608 VSS.n16929 VSS.n16433 16.666
R16609 VSS.n16923 VSS.n16437 16.666
R16610 VSS.n16917 VSS.n16432 16.666
R16611 VSS.n16911 VSS.n16438 16.666
R16612 VSS.n16905 VSS.n16431 16.666
R16613 VSS.n16946 VSS.n16440 16.666
R16614 VSS.n16774 VSS.n16540 16.666
R16615 VSS.n16848 VSS.n16526 16.666
R16616 VSS.n16839 VSS.n16523 16.666
R16617 VSS.n16833 VSS.n16527 16.666
R16618 VSS.n16827 VSS.n16522 16.666
R16619 VSS.n16821 VSS.n16528 16.666
R16620 VSS.n16815 VSS.n16521 16.666
R16621 VSS.n16856 VSS.n16530 16.666
R16622 VSS.n16684 VSS.n16630 16.666
R16623 VSS.n16758 VSS.n16616 16.666
R16624 VSS.n16749 VSS.n16613 16.666
R16625 VSS.n16743 VSS.n16617 16.666
R16626 VSS.n16737 VSS.n16612 16.666
R16627 VSS.n16731 VSS.n16618 16.666
R16628 VSS.n16725 VSS.n16611 16.666
R16629 VSS.n16766 VSS.n16620 16.666
R16630 VSS.n11097 VSS.n11083 16.666
R16631 VSS.n11226 VSS.n11080 16.666
R16632 VSS.n11217 VSS.n11084 16.666
R16633 VSS.n11211 VSS.n11079 16.666
R16634 VSS.n11205 VSS.n11085 16.666
R16635 VSS.n11199 VSS.n11078 16.666
R16636 VSS.n11233 VSS.n11087 16.666
R16637 VSS.n11188 VSS.n11082 16.666
R16638 VSS.n11180 VSS.n11062 16.666
R16639 VSS.n11007 VSS.n10993 16.666
R16640 VSS.n11316 VSS.n10990 16.666
R16641 VSS.n11307 VSS.n10994 16.666
R16642 VSS.n11301 VSS.n10989 16.666
R16643 VSS.n11295 VSS.n10995 16.666
R16644 VSS.n11289 VSS.n10988 16.666
R16645 VSS.n11323 VSS.n10997 16.666
R16646 VSS.n11278 VSS.n10992 16.666
R16647 VSS.n11270 VSS.n10972 16.666
R16648 VSS.n10917 VSS.n10903 16.666
R16649 VSS.n11406 VSS.n10900 16.666
R16650 VSS.n11397 VSS.n10904 16.666
R16651 VSS.n11391 VSS.n10899 16.666
R16652 VSS.n11385 VSS.n10905 16.666
R16653 VSS.n11379 VSS.n10898 16.666
R16654 VSS.n11413 VSS.n10907 16.666
R16655 VSS.n11368 VSS.n10902 16.666
R16656 VSS.n11360 VSS.n10882 16.666
R16657 VSS.n10827 VSS.n10813 16.666
R16658 VSS.n13526 VSS.n10810 16.666
R16659 VSS.n13517 VSS.n10814 16.666
R16660 VSS.n13510 VSS.n10809 16.666
R16661 VSS.n13504 VSS.n10815 16.666
R16662 VSS.n13498 VSS.n10808 16.666
R16663 VSS.n13533 VSS.n10817 16.666
R16664 VSS.n13487 VSS.n10812 16.666
R16665 VSS.n13479 VSS.n10792 16.666
R16666 VSS.n10737 VSS.n10723 16.666
R16667 VSS.n13616 VSS.n10720 16.666
R16668 VSS.n13607 VSS.n10724 16.666
R16669 VSS.n13601 VSS.n10719 16.666
R16670 VSS.n13595 VSS.n10725 16.666
R16671 VSS.n13589 VSS.n10718 16.666
R16672 VSS.n13623 VSS.n10727 16.666
R16673 VSS.n13578 VSS.n10722 16.666
R16674 VSS.n13570 VSS.n10702 16.666
R16675 VSS.n10647 VSS.n10633 16.666
R16676 VSS.n13706 VSS.n10630 16.666
R16677 VSS.n13697 VSS.n10634 16.666
R16678 VSS.n13691 VSS.n10629 16.666
R16679 VSS.n13685 VSS.n10635 16.666
R16680 VSS.n13679 VSS.n10628 16.666
R16681 VSS.n13713 VSS.n10637 16.666
R16682 VSS.n13668 VSS.n10632 16.666
R16683 VSS.n13660 VSS.n10612 16.666
R16684 VSS.n10557 VSS.n10543 16.666
R16685 VSS.n13796 VSS.n10540 16.666
R16686 VSS.n13787 VSS.n10544 16.666
R16687 VSS.n13781 VSS.n10539 16.666
R16688 VSS.n13775 VSS.n10545 16.666
R16689 VSS.n13769 VSS.n10538 16.666
R16690 VSS.n13803 VSS.n10547 16.666
R16691 VSS.n13758 VSS.n10542 16.666
R16692 VSS.n13750 VSS.n10522 16.666
R16693 VSS.n13886 VSS.n13885 16.666
R16694 VSS.n10514 VSS.n10503 16.666
R16695 VSS.n13946 VSS.n10505 16.666
R16696 VSS.n13937 VSS.n10502 16.666
R16697 VSS.n13931 VSS.n10506 16.666
R16698 VSS.n13925 VSS.n10501 16.666
R16699 VSS.n13919 VSS.n10507 16.666
R16700 VSS.n10500 VSS.n10499 16.666
R16701 VSS.n13954 VSS.n13953 16.666
R16702 VSS.n9034 VSS.n8985 16.666
R16703 VSS.n9042 VSS.n8989 16.666
R16704 VSS.n9050 VSS.n8988 16.666
R16705 VSS.n9058 VSS.n8990 16.666
R16706 VSS.n9066 VSS.n8987 16.666
R16707 VSS.n9074 VSS.n8991 16.666
R16708 VSS.n9082 VSS.n8986 16.666
R16709 VSS.n9090 VSS.n8992 16.666
R16710 VSS.n10179 VSS.n9225 16.666
R16711 VSS.n10253 VSS.n9211 16.666
R16712 VSS.n10244 VSS.n9208 16.666
R16713 VSS.n10238 VSS.n9212 16.666
R16714 VSS.n10232 VSS.n9207 16.666
R16715 VSS.n10226 VSS.n9213 16.666
R16716 VSS.n10220 VSS.n9206 16.666
R16717 VSS.n10261 VSS.n9215 16.666
R16718 VSS.n10089 VSS.n9315 16.666
R16719 VSS.n10163 VSS.n9301 16.666
R16720 VSS.n10154 VSS.n9298 16.666
R16721 VSS.n10148 VSS.n9302 16.666
R16722 VSS.n10142 VSS.n9297 16.666
R16723 VSS.n10136 VSS.n9303 16.666
R16724 VSS.n10130 VSS.n9296 16.666
R16725 VSS.n10171 VSS.n9305 16.666
R16726 VSS.n9999 VSS.n9405 16.666
R16727 VSS.n10073 VSS.n9391 16.666
R16728 VSS.n10064 VSS.n9388 16.666
R16729 VSS.n10058 VSS.n9392 16.666
R16730 VSS.n10052 VSS.n9387 16.666
R16731 VSS.n10046 VSS.n9393 16.666
R16732 VSS.n10040 VSS.n9386 16.666
R16733 VSS.n10081 VSS.n9395 16.666
R16734 VSS.n9909 VSS.n9495 16.666
R16735 VSS.n9983 VSS.n9481 16.666
R16736 VSS.n9974 VSS.n9478 16.666
R16737 VSS.n9968 VSS.n9482 16.666
R16738 VSS.n9962 VSS.n9477 16.666
R16739 VSS.n9956 VSS.n9483 16.666
R16740 VSS.n9950 VSS.n9476 16.666
R16741 VSS.n9991 VSS.n9485 16.666
R16742 VSS.n9819 VSS.n9585 16.666
R16743 VSS.n9893 VSS.n9571 16.666
R16744 VSS.n9884 VSS.n9568 16.666
R16745 VSS.n9878 VSS.n9572 16.666
R16746 VSS.n9872 VSS.n9567 16.666
R16747 VSS.n9866 VSS.n9573 16.666
R16748 VSS.n9860 VSS.n9566 16.666
R16749 VSS.n9901 VSS.n9575 16.666
R16750 VSS.n9729 VSS.n9675 16.666
R16751 VSS.n9803 VSS.n9661 16.666
R16752 VSS.n9794 VSS.n9658 16.666
R16753 VSS.n9788 VSS.n9662 16.666
R16754 VSS.n9782 VSS.n9657 16.666
R16755 VSS.n9776 VSS.n9663 16.666
R16756 VSS.n9770 VSS.n9656 16.666
R16757 VSS.n9811 VSS.n9665 16.666
R16758 VSS.n10323 VSS.n9180 16.666
R16759 VSS.n10368 VSS.n8934 16.666
R16760 VSS.n10362 VSS.n8936 16.666
R16761 VSS.n10356 VSS.n8941 16.666
R16762 VSS.n10350 VSS.n8947 16.666
R16763 VSS.n10344 VSS.n8953 16.666
R16764 VSS.n10338 VSS.n8958 16.666
R16765 VSS.n10332 VSS.n8965 16.666
R16766 VSS.n5783 VSS.n3581 16.666
R16767 VSS.n5777 VSS.n3583 16.666
R16768 VSS.n5771 VSS.n3588 16.666
R16769 VSS.n5765 VSS.n3594 16.666
R16770 VSS.n5759 VSS.n3600 16.666
R16771 VSS.n5753 VSS.n3606 16.666
R16772 VSS.n5747 VSS.n3611 16.666
R16773 VSS.n5741 VSS.n3618 16.666
R16774 VSS.n5905 VSS.n3523 16.666
R16775 VSS.n5899 VSS.n3525 16.666
R16776 VSS.n5893 VSS.n3530 16.666
R16777 VSS.n5887 VSS.n3536 16.666
R16778 VSS.n5881 VSS.n3542 16.666
R16779 VSS.n5875 VSS.n3548 16.666
R16780 VSS.n5869 VSS.n3553 16.666
R16781 VSS.n5863 VSS.n3560 16.666
R16782 VSS.n6027 VSS.n3465 16.666
R16783 VSS.n6021 VSS.n3467 16.666
R16784 VSS.n6015 VSS.n3472 16.666
R16785 VSS.n6009 VSS.n3478 16.666
R16786 VSS.n6003 VSS.n3484 16.666
R16787 VSS.n5997 VSS.n3490 16.666
R16788 VSS.n5991 VSS.n3495 16.666
R16789 VSS.n5985 VSS.n3502 16.666
R16790 VSS.n6149 VSS.n3407 16.666
R16791 VSS.n6143 VSS.n3409 16.666
R16792 VSS.n6137 VSS.n3414 16.666
R16793 VSS.n6131 VSS.n3420 16.666
R16794 VSS.n6125 VSS.n3426 16.666
R16795 VSS.n6119 VSS.n3432 16.666
R16796 VSS.n6113 VSS.n3437 16.666
R16797 VSS.n6107 VSS.n3444 16.666
R16798 VSS.n6271 VSS.n3349 16.666
R16799 VSS.n6265 VSS.n3351 16.666
R16800 VSS.n6259 VSS.n3356 16.666
R16801 VSS.n6253 VSS.n3362 16.666
R16802 VSS.n6247 VSS.n3368 16.666
R16803 VSS.n6241 VSS.n3374 16.666
R16804 VSS.n6235 VSS.n3379 16.666
R16805 VSS.n6229 VSS.n3386 16.666
R16806 VSS.n6393 VSS.n3291 16.666
R16807 VSS.n6387 VSS.n3293 16.666
R16808 VSS.n6381 VSS.n3298 16.666
R16809 VSS.n6375 VSS.n3304 16.666
R16810 VSS.n6369 VSS.n3310 16.666
R16811 VSS.n6363 VSS.n3316 16.666
R16812 VSS.n6357 VSS.n3321 16.666
R16813 VSS.n6351 VSS.n3328 16.666
R16814 VSS.n6515 VSS.n3233 16.666
R16815 VSS.n6509 VSS.n3235 16.666
R16816 VSS.n6503 VSS.n3240 16.666
R16817 VSS.n6497 VSS.n3246 16.666
R16818 VSS.n6491 VSS.n3252 16.666
R16819 VSS.n6485 VSS.n3258 16.666
R16820 VSS.n6479 VSS.n3263 16.666
R16821 VSS.n6473 VSS.n3270 16.666
R16822 VSS.n6535 VSS.n6534 16.666
R16823 VSS.n6599 VSS.n3141 16.666
R16824 VSS.n3182 VSS.n3144 16.666
R16825 VSS.n3190 VSS.n3146 16.666
R16826 VSS.n3198 VSS.n3143 16.666
R16827 VSS.n3206 VSS.n3147 16.666
R16828 VSS.n3214 VSS.n3142 16.666
R16829 VSS.n3222 VSS.n3148 16.666
R16830 VSS.n1177 VSS.n42 16.666
R16831 VSS.n1246 VSS.n28 16.666
R16832 VSS.n1237 VSS.n25 16.666
R16833 VSS.n1231 VSS.n29 16.666
R16834 VSS.n1225 VSS.n24 16.666
R16835 VSS.n1219 VSS.n30 16.666
R16836 VSS.n1213 VSS.n23 16.666
R16837 VSS.n1253 VSS.n32 16.666
R16838 VSS.n1087 VSS.n133 16.666
R16839 VSS.n1161 VSS.n119 16.666
R16840 VSS.n1152 VSS.n116 16.666
R16841 VSS.n1146 VSS.n120 16.666
R16842 VSS.n1140 VSS.n115 16.666
R16843 VSS.n1134 VSS.n121 16.666
R16844 VSS.n1128 VSS.n114 16.666
R16845 VSS.n1169 VSS.n123 16.666
R16846 VSS.n997 VSS.n223 16.666
R16847 VSS.n1071 VSS.n209 16.666
R16848 VSS.n1062 VSS.n206 16.666
R16849 VSS.n1056 VSS.n210 16.666
R16850 VSS.n1050 VSS.n205 16.666
R16851 VSS.n1044 VSS.n211 16.666
R16852 VSS.n1038 VSS.n204 16.666
R16853 VSS.n1079 VSS.n213 16.666
R16854 VSS.n907 VSS.n313 16.666
R16855 VSS.n981 VSS.n299 16.666
R16856 VSS.n972 VSS.n296 16.666
R16857 VSS.n966 VSS.n300 16.666
R16858 VSS.n960 VSS.n295 16.666
R16859 VSS.n954 VSS.n301 16.666
R16860 VSS.n948 VSS.n294 16.666
R16861 VSS.n989 VSS.n303 16.666
R16862 VSS.n817 VSS.n403 16.666
R16863 VSS.n891 VSS.n389 16.666
R16864 VSS.n882 VSS.n386 16.666
R16865 VSS.n876 VSS.n390 16.666
R16866 VSS.n870 VSS.n385 16.666
R16867 VSS.n864 VSS.n391 16.666
R16868 VSS.n858 VSS.n384 16.666
R16869 VSS.n899 VSS.n393 16.666
R16870 VSS.n727 VSS.n493 16.666
R16871 VSS.n801 VSS.n479 16.666
R16872 VSS.n792 VSS.n476 16.666
R16873 VSS.n786 VSS.n480 16.666
R16874 VSS.n780 VSS.n475 16.666
R16875 VSS.n774 VSS.n481 16.666
R16876 VSS.n768 VSS.n474 16.666
R16877 VSS.n809 VSS.n483 16.666
R16878 VSS.n637 VSS.n583 16.666
R16879 VSS.n711 VSS.n569 16.666
R16880 VSS.n702 VSS.n566 16.666
R16881 VSS.n696 VSS.n570 16.666
R16882 VSS.n690 VSS.n565 16.666
R16883 VSS.n684 VSS.n571 16.666
R16884 VSS.n678 VSS.n564 16.666
R16885 VSS.n719 VSS.n573 16.666
R16886 sky130_asc_pnp_05v5_W3p40L3p40_7_0/Collector VSS.n1267 16.505
R16887 VSS.n17337 VSS.n17335 16
R16888 VSS.n17338 VSS.n17337 16
R16889 VSS.n17341 VSS.n17338 16
R16890 VSS.n17342 VSS.n17341 16
R16891 VSS.n17345 VSS.n17342 16
R16892 VSS.n17346 VSS.n17345 16
R16893 VSS.n17349 VSS.n17346 16
R16894 VSS.n17351 VSS.n17349 16
R16895 VSS.n17367 VSS.n17366 16
R16896 VSS.n17366 VSS.n17363 16
R16897 VSS.n17363 VSS.n17362 16
R16898 VSS.n17362 VSS.n17359 16
R16899 VSS.n17359 VSS.n17358 16
R16900 VSS.n17358 VSS.n17355 16
R16901 VSS.n17355 VSS.n17354 16
R16902 VSS.n17354 VSS.n17352 16
R16903 VSS.n17382 VSS.n17330 16
R16904 VSS.n17382 VSS.n17381 16
R16905 VSS.n17381 VSS.n17380 16
R16906 VSS.n17380 VSS.n17378 16
R16907 VSS.n17378 VSS.n17375 16
R16908 VSS.n17375 VSS.n17374 16
R16909 VSS.n17374 VSS.n17371 16
R16910 VSS.n17371 VSS.n17370 16
R16911 VSS.n17308 VSS.n16054 16
R16912 VSS.n16094 VSS.n16054 16
R16913 VSS.n16097 VSS.n16094 16
R16914 VSS.n16098 VSS.n16097 16
R16915 VSS.n16101 VSS.n16098 16
R16916 VSS.n16102 VSS.n16101 16
R16917 VSS.n16105 VSS.n16102 16
R16918 VSS.n16107 VSS.n16105 16
R16919 VSS.n16123 VSS.n16122 16
R16920 VSS.n16122 VSS.n16119 16
R16921 VSS.n16119 VSS.n16118 16
R16922 VSS.n16118 VSS.n16115 16
R16923 VSS.n16115 VSS.n16114 16
R16924 VSS.n16114 VSS.n16111 16
R16925 VSS.n16111 VSS.n16110 16
R16926 VSS.n16110 VSS.n16108 16
R16927 VSS.n16141 VSS.n16140 16
R16928 VSS.n16140 VSS.n16138 16
R16929 VSS.n16138 VSS.n16135 16
R16930 VSS.n16135 VSS.n16134 16
R16931 VSS.n16134 VSS.n16131 16
R16932 VSS.n16131 VSS.n16130 16
R16933 VSS.n16130 VSS.n16127 16
R16934 VSS.n16127 VSS.n16126 16
R16935 VSS.n17218 VSS.n16144 16
R16936 VSS.n16184 VSS.n16144 16
R16937 VSS.n16187 VSS.n16184 16
R16938 VSS.n16188 VSS.n16187 16
R16939 VSS.n16191 VSS.n16188 16
R16940 VSS.n16192 VSS.n16191 16
R16941 VSS.n16195 VSS.n16192 16
R16942 VSS.n16197 VSS.n16195 16
R16943 VSS.n16213 VSS.n16212 16
R16944 VSS.n16212 VSS.n16209 16
R16945 VSS.n16209 VSS.n16208 16
R16946 VSS.n16208 VSS.n16205 16
R16947 VSS.n16205 VSS.n16204 16
R16948 VSS.n16204 VSS.n16201 16
R16949 VSS.n16201 VSS.n16200 16
R16950 VSS.n16200 VSS.n16198 16
R16951 VSS.n16231 VSS.n16230 16
R16952 VSS.n16230 VSS.n16228 16
R16953 VSS.n16228 VSS.n16225 16
R16954 VSS.n16225 VSS.n16224 16
R16955 VSS.n16224 VSS.n16221 16
R16956 VSS.n16221 VSS.n16220 16
R16957 VSS.n16220 VSS.n16217 16
R16958 VSS.n16217 VSS.n16216 16
R16959 VSS.n17128 VSS.n16234 16
R16960 VSS.n16274 VSS.n16234 16
R16961 VSS.n16277 VSS.n16274 16
R16962 VSS.n16278 VSS.n16277 16
R16963 VSS.n16281 VSS.n16278 16
R16964 VSS.n16282 VSS.n16281 16
R16965 VSS.n16285 VSS.n16282 16
R16966 VSS.n16287 VSS.n16285 16
R16967 VSS.n16303 VSS.n16302 16
R16968 VSS.n16302 VSS.n16299 16
R16969 VSS.n16299 VSS.n16298 16
R16970 VSS.n16298 VSS.n16295 16
R16971 VSS.n16295 VSS.n16294 16
R16972 VSS.n16294 VSS.n16291 16
R16973 VSS.n16291 VSS.n16290 16
R16974 VSS.n16290 VSS.n16288 16
R16975 VSS.n16321 VSS.n16320 16
R16976 VSS.n16320 VSS.n16318 16
R16977 VSS.n16318 VSS.n16315 16
R16978 VSS.n16315 VSS.n16314 16
R16979 VSS.n16314 VSS.n16311 16
R16980 VSS.n16311 VSS.n16310 16
R16981 VSS.n16310 VSS.n16307 16
R16982 VSS.n16307 VSS.n16306 16
R16983 VSS.n17038 VSS.n16324 16
R16984 VSS.n16364 VSS.n16324 16
R16985 VSS.n16367 VSS.n16364 16
R16986 VSS.n16368 VSS.n16367 16
R16987 VSS.n16371 VSS.n16368 16
R16988 VSS.n16372 VSS.n16371 16
R16989 VSS.n16375 VSS.n16372 16
R16990 VSS.n16377 VSS.n16375 16
R16991 VSS.n16393 VSS.n16392 16
R16992 VSS.n16392 VSS.n16389 16
R16993 VSS.n16389 VSS.n16388 16
R16994 VSS.n16388 VSS.n16385 16
R16995 VSS.n16385 VSS.n16384 16
R16996 VSS.n16384 VSS.n16381 16
R16997 VSS.n16381 VSS.n16380 16
R16998 VSS.n16380 VSS.n16378 16
R16999 VSS.n16411 VSS.n16410 16
R17000 VSS.n16410 VSS.n16408 16
R17001 VSS.n16408 VSS.n16405 16
R17002 VSS.n16405 VSS.n16404 16
R17003 VSS.n16404 VSS.n16401 16
R17004 VSS.n16401 VSS.n16400 16
R17005 VSS.n16400 VSS.n16397 16
R17006 VSS.n16397 VSS.n16396 16
R17007 VSS.n16948 VSS.n16414 16
R17008 VSS.n16454 VSS.n16414 16
R17009 VSS.n16457 VSS.n16454 16
R17010 VSS.n16458 VSS.n16457 16
R17011 VSS.n16461 VSS.n16458 16
R17012 VSS.n16462 VSS.n16461 16
R17013 VSS.n16465 VSS.n16462 16
R17014 VSS.n16467 VSS.n16465 16
R17015 VSS.n16483 VSS.n16482 16
R17016 VSS.n16482 VSS.n16479 16
R17017 VSS.n16479 VSS.n16478 16
R17018 VSS.n16478 VSS.n16475 16
R17019 VSS.n16475 VSS.n16474 16
R17020 VSS.n16474 VSS.n16471 16
R17021 VSS.n16471 VSS.n16470 16
R17022 VSS.n16470 VSS.n16468 16
R17023 VSS.n16501 VSS.n16500 16
R17024 VSS.n16500 VSS.n16498 16
R17025 VSS.n16498 VSS.n16495 16
R17026 VSS.n16495 VSS.n16494 16
R17027 VSS.n16494 VSS.n16491 16
R17028 VSS.n16491 VSS.n16490 16
R17029 VSS.n16490 VSS.n16487 16
R17030 VSS.n16487 VSS.n16486 16
R17031 VSS.n16858 VSS.n16504 16
R17032 VSS.n16544 VSS.n16504 16
R17033 VSS.n16547 VSS.n16544 16
R17034 VSS.n16548 VSS.n16547 16
R17035 VSS.n16551 VSS.n16548 16
R17036 VSS.n16552 VSS.n16551 16
R17037 VSS.n16555 VSS.n16552 16
R17038 VSS.n16557 VSS.n16555 16
R17039 VSS.n16573 VSS.n16572 16
R17040 VSS.n16572 VSS.n16569 16
R17041 VSS.n16569 VSS.n16568 16
R17042 VSS.n16568 VSS.n16565 16
R17043 VSS.n16565 VSS.n16564 16
R17044 VSS.n16564 VSS.n16561 16
R17045 VSS.n16561 VSS.n16560 16
R17046 VSS.n16560 VSS.n16558 16
R17047 VSS.n16591 VSS.n16590 16
R17048 VSS.n16590 VSS.n16588 16
R17049 VSS.n16588 VSS.n16585 16
R17050 VSS.n16585 VSS.n16584 16
R17051 VSS.n16584 VSS.n16581 16
R17052 VSS.n16581 VSS.n16580 16
R17053 VSS.n16580 VSS.n16577 16
R17054 VSS.n16577 VSS.n16576 16
R17055 VSS.n16768 VSS.n16594 16
R17056 VSS.n16634 VSS.n16594 16
R17057 VSS.n16637 VSS.n16634 16
R17058 VSS.n16638 VSS.n16637 16
R17059 VSS.n16641 VSS.n16638 16
R17060 VSS.n16642 VSS.n16641 16
R17061 VSS.n16645 VSS.n16642 16
R17062 VSS.n16647 VSS.n16645 16
R17063 VSS.n16663 VSS.n16662 16
R17064 VSS.n16662 VSS.n16659 16
R17065 VSS.n16659 VSS.n16658 16
R17066 VSS.n16658 VSS.n16655 16
R17067 VSS.n16655 VSS.n16654 16
R17068 VSS.n16654 VSS.n16651 16
R17069 VSS.n16651 VSS.n16650 16
R17070 VSS.n16650 VSS.n16648 16
R17071 VSS.n16681 VSS.n16680 16
R17072 VSS.n16680 VSS.n16678 16
R17073 VSS.n16678 VSS.n16675 16
R17074 VSS.n16675 VSS.n16674 16
R17075 VSS.n16674 VSS.n16671 16
R17076 VSS.n16671 VSS.n16670 16
R17077 VSS.n16670 VSS.n16667 16
R17078 VSS.n16667 VSS.n16666 16
R17079 VSS.n11235 VSS.n11061 16
R17080 VSS.n11101 VSS.n11061 16
R17081 VSS.n11104 VSS.n11101 16
R17082 VSS.n11105 VSS.n11104 16
R17083 VSS.n11108 VSS.n11105 16
R17084 VSS.n11109 VSS.n11108 16
R17085 VSS.n11112 VSS.n11109 16
R17086 VSS.n11114 VSS.n11112 16
R17087 VSS.n11130 VSS.n11129 16
R17088 VSS.n11129 VSS.n11126 16
R17089 VSS.n11126 VSS.n11125 16
R17090 VSS.n11125 VSS.n11122 16
R17091 VSS.n11122 VSS.n11121 16
R17092 VSS.n11121 VSS.n11118 16
R17093 VSS.n11118 VSS.n11117 16
R17094 VSS.n11117 VSS.n11115 16
R17095 VSS.n11148 VSS.n11147 16
R17096 VSS.n11147 VSS.n11145 16
R17097 VSS.n11145 VSS.n11142 16
R17098 VSS.n11142 VSS.n11141 16
R17099 VSS.n11141 VSS.n11138 16
R17100 VSS.n11138 VSS.n11137 16
R17101 VSS.n11137 VSS.n11134 16
R17102 VSS.n11134 VSS.n11133 16
R17103 VSS.n11325 VSS.n10971 16
R17104 VSS.n11011 VSS.n10971 16
R17105 VSS.n11014 VSS.n11011 16
R17106 VSS.n11015 VSS.n11014 16
R17107 VSS.n11018 VSS.n11015 16
R17108 VSS.n11019 VSS.n11018 16
R17109 VSS.n11022 VSS.n11019 16
R17110 VSS.n11024 VSS.n11022 16
R17111 VSS.n11040 VSS.n11039 16
R17112 VSS.n11039 VSS.n11036 16
R17113 VSS.n11036 VSS.n11035 16
R17114 VSS.n11035 VSS.n11032 16
R17115 VSS.n11032 VSS.n11031 16
R17116 VSS.n11031 VSS.n11028 16
R17117 VSS.n11028 VSS.n11027 16
R17118 VSS.n11027 VSS.n11025 16
R17119 VSS.n11058 VSS.n11057 16
R17120 VSS.n11057 VSS.n11055 16
R17121 VSS.n11055 VSS.n11052 16
R17122 VSS.n11052 VSS.n11051 16
R17123 VSS.n11051 VSS.n11048 16
R17124 VSS.n11048 VSS.n11047 16
R17125 VSS.n11047 VSS.n11044 16
R17126 VSS.n11044 VSS.n11043 16
R17127 VSS.n11415 VSS.n10881 16
R17128 VSS.n10921 VSS.n10881 16
R17129 VSS.n10924 VSS.n10921 16
R17130 VSS.n10925 VSS.n10924 16
R17131 VSS.n10928 VSS.n10925 16
R17132 VSS.n10929 VSS.n10928 16
R17133 VSS.n10932 VSS.n10929 16
R17134 VSS.n10934 VSS.n10932 16
R17135 VSS.n10950 VSS.n10949 16
R17136 VSS.n10949 VSS.n10946 16
R17137 VSS.n10946 VSS.n10945 16
R17138 VSS.n10945 VSS.n10942 16
R17139 VSS.n10942 VSS.n10941 16
R17140 VSS.n10941 VSS.n10938 16
R17141 VSS.n10938 VSS.n10937 16
R17142 VSS.n10937 VSS.n10935 16
R17143 VSS.n10968 VSS.n10967 16
R17144 VSS.n10967 VSS.n10965 16
R17145 VSS.n10965 VSS.n10962 16
R17146 VSS.n10962 VSS.n10961 16
R17147 VSS.n10961 VSS.n10958 16
R17148 VSS.n10958 VSS.n10957 16
R17149 VSS.n10957 VSS.n10954 16
R17150 VSS.n10954 VSS.n10953 16
R17151 VSS.n13535 VSS.n10791 16
R17152 VSS.n10831 VSS.n10791 16
R17153 VSS.n10834 VSS.n10831 16
R17154 VSS.n10835 VSS.n10834 16
R17155 VSS.n10838 VSS.n10835 16
R17156 VSS.n10839 VSS.n10838 16
R17157 VSS.n10842 VSS.n10839 16
R17158 VSS.n10844 VSS.n10842 16
R17159 VSS.n10860 VSS.n10859 16
R17160 VSS.n10859 VSS.n10856 16
R17161 VSS.n10856 VSS.n10855 16
R17162 VSS.n10855 VSS.n10852 16
R17163 VSS.n10852 VSS.n10851 16
R17164 VSS.n10851 VSS.n10848 16
R17165 VSS.n10848 VSS.n10847 16
R17166 VSS.n10847 VSS.n10845 16
R17167 VSS.n10878 VSS.n10877 16
R17168 VSS.n10877 VSS.n10875 16
R17169 VSS.n10875 VSS.n10872 16
R17170 VSS.n10872 VSS.n10871 16
R17171 VSS.n10871 VSS.n10868 16
R17172 VSS.n10868 VSS.n10867 16
R17173 VSS.n10867 VSS.n10864 16
R17174 VSS.n10864 VSS.n10863 16
R17175 VSS.n13625 VSS.n10701 16
R17176 VSS.n10741 VSS.n10701 16
R17177 VSS.n10744 VSS.n10741 16
R17178 VSS.n10745 VSS.n10744 16
R17179 VSS.n10748 VSS.n10745 16
R17180 VSS.n10749 VSS.n10748 16
R17181 VSS.n10752 VSS.n10749 16
R17182 VSS.n10754 VSS.n10752 16
R17183 VSS.n10770 VSS.n10769 16
R17184 VSS.n10769 VSS.n10766 16
R17185 VSS.n10766 VSS.n10765 16
R17186 VSS.n10765 VSS.n10762 16
R17187 VSS.n10762 VSS.n10761 16
R17188 VSS.n10761 VSS.n10758 16
R17189 VSS.n10758 VSS.n10757 16
R17190 VSS.n10757 VSS.n10755 16
R17191 VSS.n10788 VSS.n10787 16
R17192 VSS.n10787 VSS.n10785 16
R17193 VSS.n10785 VSS.n10782 16
R17194 VSS.n10782 VSS.n10781 16
R17195 VSS.n10781 VSS.n10778 16
R17196 VSS.n10778 VSS.n10777 16
R17197 VSS.n10777 VSS.n10774 16
R17198 VSS.n10774 VSS.n10773 16
R17199 VSS.n13715 VSS.n10611 16
R17200 VSS.n10651 VSS.n10611 16
R17201 VSS.n10654 VSS.n10651 16
R17202 VSS.n10655 VSS.n10654 16
R17203 VSS.n10658 VSS.n10655 16
R17204 VSS.n10659 VSS.n10658 16
R17205 VSS.n10662 VSS.n10659 16
R17206 VSS.n10664 VSS.n10662 16
R17207 VSS.n10680 VSS.n10679 16
R17208 VSS.n10679 VSS.n10676 16
R17209 VSS.n10676 VSS.n10675 16
R17210 VSS.n10675 VSS.n10672 16
R17211 VSS.n10672 VSS.n10671 16
R17212 VSS.n10671 VSS.n10668 16
R17213 VSS.n10668 VSS.n10667 16
R17214 VSS.n10667 VSS.n10665 16
R17215 VSS.n10698 VSS.n10697 16
R17216 VSS.n10697 VSS.n10695 16
R17217 VSS.n10695 VSS.n10692 16
R17218 VSS.n10692 VSS.n10691 16
R17219 VSS.n10691 VSS.n10688 16
R17220 VSS.n10688 VSS.n10687 16
R17221 VSS.n10687 VSS.n10684 16
R17222 VSS.n10684 VSS.n10683 16
R17223 VSS.n13805 VSS.n10521 16
R17224 VSS.n10561 VSS.n10521 16
R17225 VSS.n10564 VSS.n10561 16
R17226 VSS.n10565 VSS.n10564 16
R17227 VSS.n10568 VSS.n10565 16
R17228 VSS.n10569 VSS.n10568 16
R17229 VSS.n10572 VSS.n10569 16
R17230 VSS.n10574 VSS.n10572 16
R17231 VSS.n10590 VSS.n10589 16
R17232 VSS.n10589 VSS.n10586 16
R17233 VSS.n10586 VSS.n10585 16
R17234 VSS.n10585 VSS.n10582 16
R17235 VSS.n10582 VSS.n10581 16
R17236 VSS.n10581 VSS.n10578 16
R17237 VSS.n10578 VSS.n10577 16
R17238 VSS.n10577 VSS.n10575 16
R17239 VSS.n10608 VSS.n10607 16
R17240 VSS.n10607 VSS.n10605 16
R17241 VSS.n10605 VSS.n10602 16
R17242 VSS.n10602 VSS.n10601 16
R17243 VSS.n10601 VSS.n10598 16
R17244 VSS.n10598 VSS.n10597 16
R17245 VSS.n10597 VSS.n10594 16
R17246 VSS.n10594 VSS.n10593 16
R17247 VSS.n13837 VSS.n13835 16
R17248 VSS.n13838 VSS.n13837 16
R17249 VSS.n13841 VSS.n13838 16
R17250 VSS.n13842 VSS.n13841 16
R17251 VSS.n13845 VSS.n13842 16
R17252 VSS.n13846 VSS.n13845 16
R17253 VSS.n13849 VSS.n13846 16
R17254 VSS.n13851 VSS.n13849 16
R17255 VSS.n13867 VSS.n13866 16
R17256 VSS.n13866 VSS.n13863 16
R17257 VSS.n13863 VSS.n13862 16
R17258 VSS.n13862 VSS.n13859 16
R17259 VSS.n13859 VSS.n13858 16
R17260 VSS.n13858 VSS.n13855 16
R17261 VSS.n13855 VSS.n13854 16
R17262 VSS.n13854 VSS.n13852 16
R17263 VSS.n13882 VSS.n13827 16
R17264 VSS.n13882 VSS.n13881 16
R17265 VSS.n13881 VSS.n13880 16
R17266 VSS.n13880 VSS.n13878 16
R17267 VSS.n13878 VSS.n13875 16
R17268 VSS.n13875 VSS.n13874 16
R17269 VSS.n13874 VSS.n13871 16
R17270 VSS.n13871 VSS.n13870 16
R17271 VSS.n9147 VSS.n9146 16
R17272 VSS.n9146 VSS.n9143 16
R17273 VSS.n9143 VSS.n9142 16
R17274 VSS.n9142 VSS.n9139 16
R17275 VSS.n9139 VSS.n9138 16
R17276 VSS.n9138 VSS.n9135 16
R17277 VSS.n9135 VSS.n9134 16
R17278 VSS.n9134 VSS.n9131 16
R17279 VSS.n9115 VSS.n9114 16
R17280 VSS.n9118 VSS.n9115 16
R17281 VSS.n9119 VSS.n9118 16
R17282 VSS.n9122 VSS.n9119 16
R17283 VSS.n9123 VSS.n9122 16
R17284 VSS.n9126 VSS.n9123 16
R17285 VSS.n9127 VSS.n9126 16
R17286 VSS.n9130 VSS.n9127 16
R17287 VSS.n9098 VSS.n8982 16
R17288 VSS.n9101 VSS.n9098 16
R17289 VSS.n9102 VSS.n9101 16
R17290 VSS.n9105 VSS.n9102 16
R17291 VSS.n9106 VSS.n9105 16
R17292 VSS.n9109 VSS.n9106 16
R17293 VSS.n9111 VSS.n9109 16
R17294 VSS.n9112 VSS.n9111 16
R17295 VSS.n10263 VSS.n9189 16
R17296 VSS.n9229 VSS.n9189 16
R17297 VSS.n9232 VSS.n9229 16
R17298 VSS.n9233 VSS.n9232 16
R17299 VSS.n9236 VSS.n9233 16
R17300 VSS.n9237 VSS.n9236 16
R17301 VSS.n9240 VSS.n9237 16
R17302 VSS.n9242 VSS.n9240 16
R17303 VSS.n9258 VSS.n9257 16
R17304 VSS.n9257 VSS.n9254 16
R17305 VSS.n9254 VSS.n9253 16
R17306 VSS.n9253 VSS.n9250 16
R17307 VSS.n9250 VSS.n9249 16
R17308 VSS.n9249 VSS.n9246 16
R17309 VSS.n9246 VSS.n9245 16
R17310 VSS.n9245 VSS.n9243 16
R17311 VSS.n9276 VSS.n9275 16
R17312 VSS.n9275 VSS.n9273 16
R17313 VSS.n9273 VSS.n9270 16
R17314 VSS.n9270 VSS.n9269 16
R17315 VSS.n9269 VSS.n9266 16
R17316 VSS.n9266 VSS.n9265 16
R17317 VSS.n9265 VSS.n9262 16
R17318 VSS.n9262 VSS.n9261 16
R17319 VSS.n10173 VSS.n9279 16
R17320 VSS.n9319 VSS.n9279 16
R17321 VSS.n9322 VSS.n9319 16
R17322 VSS.n9323 VSS.n9322 16
R17323 VSS.n9326 VSS.n9323 16
R17324 VSS.n9327 VSS.n9326 16
R17325 VSS.n9330 VSS.n9327 16
R17326 VSS.n9332 VSS.n9330 16
R17327 VSS.n9348 VSS.n9347 16
R17328 VSS.n9347 VSS.n9344 16
R17329 VSS.n9344 VSS.n9343 16
R17330 VSS.n9343 VSS.n9340 16
R17331 VSS.n9340 VSS.n9339 16
R17332 VSS.n9339 VSS.n9336 16
R17333 VSS.n9336 VSS.n9335 16
R17334 VSS.n9335 VSS.n9333 16
R17335 VSS.n9366 VSS.n9365 16
R17336 VSS.n9365 VSS.n9363 16
R17337 VSS.n9363 VSS.n9360 16
R17338 VSS.n9360 VSS.n9359 16
R17339 VSS.n9359 VSS.n9356 16
R17340 VSS.n9356 VSS.n9355 16
R17341 VSS.n9355 VSS.n9352 16
R17342 VSS.n9352 VSS.n9351 16
R17343 VSS.n10083 VSS.n9369 16
R17344 VSS.n9409 VSS.n9369 16
R17345 VSS.n9412 VSS.n9409 16
R17346 VSS.n9413 VSS.n9412 16
R17347 VSS.n9416 VSS.n9413 16
R17348 VSS.n9417 VSS.n9416 16
R17349 VSS.n9420 VSS.n9417 16
R17350 VSS.n9422 VSS.n9420 16
R17351 VSS.n9438 VSS.n9437 16
R17352 VSS.n9437 VSS.n9434 16
R17353 VSS.n9434 VSS.n9433 16
R17354 VSS.n9433 VSS.n9430 16
R17355 VSS.n9430 VSS.n9429 16
R17356 VSS.n9429 VSS.n9426 16
R17357 VSS.n9426 VSS.n9425 16
R17358 VSS.n9425 VSS.n9423 16
R17359 VSS.n9456 VSS.n9455 16
R17360 VSS.n9455 VSS.n9453 16
R17361 VSS.n9453 VSS.n9450 16
R17362 VSS.n9450 VSS.n9449 16
R17363 VSS.n9449 VSS.n9446 16
R17364 VSS.n9446 VSS.n9445 16
R17365 VSS.n9445 VSS.n9442 16
R17366 VSS.n9442 VSS.n9441 16
R17367 VSS.n9993 VSS.n9459 16
R17368 VSS.n9499 VSS.n9459 16
R17369 VSS.n9502 VSS.n9499 16
R17370 VSS.n9503 VSS.n9502 16
R17371 VSS.n9506 VSS.n9503 16
R17372 VSS.n9507 VSS.n9506 16
R17373 VSS.n9510 VSS.n9507 16
R17374 VSS.n9512 VSS.n9510 16
R17375 VSS.n9528 VSS.n9527 16
R17376 VSS.n9527 VSS.n9524 16
R17377 VSS.n9524 VSS.n9523 16
R17378 VSS.n9523 VSS.n9520 16
R17379 VSS.n9520 VSS.n9519 16
R17380 VSS.n9519 VSS.n9516 16
R17381 VSS.n9516 VSS.n9515 16
R17382 VSS.n9515 VSS.n9513 16
R17383 VSS.n9546 VSS.n9545 16
R17384 VSS.n9545 VSS.n9543 16
R17385 VSS.n9543 VSS.n9540 16
R17386 VSS.n9540 VSS.n9539 16
R17387 VSS.n9539 VSS.n9536 16
R17388 VSS.n9536 VSS.n9535 16
R17389 VSS.n9535 VSS.n9532 16
R17390 VSS.n9532 VSS.n9531 16
R17391 VSS.n9903 VSS.n9549 16
R17392 VSS.n9589 VSS.n9549 16
R17393 VSS.n9592 VSS.n9589 16
R17394 VSS.n9593 VSS.n9592 16
R17395 VSS.n9596 VSS.n9593 16
R17396 VSS.n9597 VSS.n9596 16
R17397 VSS.n9600 VSS.n9597 16
R17398 VSS.n9602 VSS.n9600 16
R17399 VSS.n9618 VSS.n9617 16
R17400 VSS.n9617 VSS.n9614 16
R17401 VSS.n9614 VSS.n9613 16
R17402 VSS.n9613 VSS.n9610 16
R17403 VSS.n9610 VSS.n9609 16
R17404 VSS.n9609 VSS.n9606 16
R17405 VSS.n9606 VSS.n9605 16
R17406 VSS.n9605 VSS.n9603 16
R17407 VSS.n9636 VSS.n9635 16
R17408 VSS.n9635 VSS.n9633 16
R17409 VSS.n9633 VSS.n9630 16
R17410 VSS.n9630 VSS.n9629 16
R17411 VSS.n9629 VSS.n9626 16
R17412 VSS.n9626 VSS.n9625 16
R17413 VSS.n9625 VSS.n9622 16
R17414 VSS.n9622 VSS.n9621 16
R17415 VSS.n9813 VSS.n9639 16
R17416 VSS.n9679 VSS.n9639 16
R17417 VSS.n9682 VSS.n9679 16
R17418 VSS.n9683 VSS.n9682 16
R17419 VSS.n9686 VSS.n9683 16
R17420 VSS.n9687 VSS.n9686 16
R17421 VSS.n9690 VSS.n9687 16
R17422 VSS.n9692 VSS.n9690 16
R17423 VSS.n9708 VSS.n9707 16
R17424 VSS.n9707 VSS.n9704 16
R17425 VSS.n9704 VSS.n9703 16
R17426 VSS.n9703 VSS.n9700 16
R17427 VSS.n9700 VSS.n9699 16
R17428 VSS.n9699 VSS.n9696 16
R17429 VSS.n9696 VSS.n9695 16
R17430 VSS.n9695 VSS.n9693 16
R17431 VSS.n9726 VSS.n9725 16
R17432 VSS.n9725 VSS.n9723 16
R17433 VSS.n9723 VSS.n9720 16
R17434 VSS.n9720 VSS.n9719 16
R17435 VSS.n9719 VSS.n9716 16
R17436 VSS.n9716 VSS.n9715 16
R17437 VSS.n9715 VSS.n9712 16
R17438 VSS.n9712 VSS.n9711 16
R17439 VSS.n10266 VSS.n9163 16
R17440 VSS.n10268 VSS.n10266 16
R17441 VSS.n10269 VSS.n10268 16
R17442 VSS.n10272 VSS.n10269 16
R17443 VSS.n10273 VSS.n10272 16
R17444 VSS.n10276 VSS.n10273 16
R17445 VSS.n10277 VSS.n10276 16
R17446 VSS.n10280 VSS.n10277 16
R17447 VSS.n10298 VSS.n10296 16
R17448 VSS.n10296 VSS.n10293 16
R17449 VSS.n10293 VSS.n10292 16
R17450 VSS.n10292 VSS.n10289 16
R17451 VSS.n10289 VSS.n10288 16
R17452 VSS.n10288 VSS.n10285 16
R17453 VSS.n10285 VSS.n10284 16
R17454 VSS.n10284 VSS.n10281 16
R17455 VSS.n10316 VSS.n10313 16
R17456 VSS.n10313 VSS.n10310 16
R17457 VSS.n10310 VSS.n10309 16
R17458 VSS.n10309 VSS.n10306 16
R17459 VSS.n10306 VSS.n10305 16
R17460 VSS.n10305 VSS.n10302 16
R17461 VSS.n10302 VSS.n10301 16
R17462 VSS.n10301 VSS.n10299 16
R17463 VSS.n6691 VSS.n6690 16
R17464 VSS.n6690 VSS.n6688 16
R17465 VSS.n6688 VSS.n6686 16
R17466 VSS.n6686 VSS.n6684 16
R17467 VSS.n6684 VSS.n6682 16
R17468 VSS.n6682 VSS.n6680 16
R17469 VSS.n6680 VSS.n6678 16
R17470 VSS.n6678 VSS.n6675 16
R17471 VSS.n6695 VSS.n6692 16
R17472 VSS.n6696 VSS.n6695 16
R17473 VSS.n6699 VSS.n6696 16
R17474 VSS.n6703 VSS.n6700 16
R17475 VSS.n6707 VSS.n6704 16
R17476 VSS.n6708 VSS.n6707 16
R17477 VSS.n6712 VSS.n6711 16
R17478 VSS.n6715 VSS.n6712 16
R17479 VSS.n6716 VSS.n6715 16
R17480 VSS.n6719 VSS.n6716 16
R17481 VSS.n6720 VSS.n6719 16
R17482 VSS.n6722 VSS.n6720 16
R17483 VSS.n6722 VSS.n6721 16
R17484 VSS.n6721 VSS.n6635 16
R17485 VSS.n6674 VSS.n6671 16
R17486 VSS.n6671 VSS.n6670 16
R17487 VSS.n6670 VSS.n6667 16
R17488 VSS.n6667 VSS.n6666 16
R17489 VSS.n6666 VSS.n6663 16
R17490 VSS.n6663 VSS.n6662 16
R17491 VSS.n6662 VSS.n6636 16
R17492 VSS.n6727 VSS.n6636 16
R17493 VSS.n5685 VSS.n5667 16
R17494 VSS.n5686 VSS.n5685 16
R17495 VSS.n5689 VSS.n5686 16
R17496 VSS.n5690 VSS.n5689 16
R17497 VSS.n5693 VSS.n5690 16
R17498 VSS.n5694 VSS.n5693 16
R17499 VSS.n5697 VSS.n5694 16
R17500 VSS.n5699 VSS.n5697 16
R17501 VSS.n5715 VSS.n5714 16
R17502 VSS.n5714 VSS.n5711 16
R17503 VSS.n5711 VSS.n5710 16
R17504 VSS.n5710 VSS.n5707 16
R17505 VSS.n5707 VSS.n5706 16
R17506 VSS.n5706 VSS.n5703 16
R17507 VSS.n5703 VSS.n5702 16
R17508 VSS.n5702 VSS.n5700 16
R17509 VSS.n5730 VSS.n5684 16
R17510 VSS.n5730 VSS.n5729 16
R17511 VSS.n5729 VSS.n5728 16
R17512 VSS.n5728 VSS.n5726 16
R17513 VSS.n5726 VSS.n5723 16
R17514 VSS.n5723 VSS.n5722 16
R17515 VSS.n5722 VSS.n5719 16
R17516 VSS.n5719 VSS.n5718 16
R17517 VSS.n5807 VSS.n5789 16
R17518 VSS.n5808 VSS.n5807 16
R17519 VSS.n5811 VSS.n5808 16
R17520 VSS.n5812 VSS.n5811 16
R17521 VSS.n5815 VSS.n5812 16
R17522 VSS.n5816 VSS.n5815 16
R17523 VSS.n5819 VSS.n5816 16
R17524 VSS.n5821 VSS.n5819 16
R17525 VSS.n5837 VSS.n5836 16
R17526 VSS.n5836 VSS.n5833 16
R17527 VSS.n5833 VSS.n5832 16
R17528 VSS.n5832 VSS.n5829 16
R17529 VSS.n5829 VSS.n5828 16
R17530 VSS.n5828 VSS.n5825 16
R17531 VSS.n5825 VSS.n5824 16
R17532 VSS.n5824 VSS.n5822 16
R17533 VSS.n5852 VSS.n5806 16
R17534 VSS.n5852 VSS.n5851 16
R17535 VSS.n5851 VSS.n5850 16
R17536 VSS.n5850 VSS.n5848 16
R17537 VSS.n5848 VSS.n5845 16
R17538 VSS.n5845 VSS.n5844 16
R17539 VSS.n5844 VSS.n5841 16
R17540 VSS.n5841 VSS.n5840 16
R17541 VSS.n5929 VSS.n5911 16
R17542 VSS.n5930 VSS.n5929 16
R17543 VSS.n5933 VSS.n5930 16
R17544 VSS.n5934 VSS.n5933 16
R17545 VSS.n5937 VSS.n5934 16
R17546 VSS.n5938 VSS.n5937 16
R17547 VSS.n5941 VSS.n5938 16
R17548 VSS.n5943 VSS.n5941 16
R17549 VSS.n5959 VSS.n5958 16
R17550 VSS.n5958 VSS.n5955 16
R17551 VSS.n5955 VSS.n5954 16
R17552 VSS.n5954 VSS.n5951 16
R17553 VSS.n5951 VSS.n5950 16
R17554 VSS.n5950 VSS.n5947 16
R17555 VSS.n5947 VSS.n5946 16
R17556 VSS.n5946 VSS.n5944 16
R17557 VSS.n5974 VSS.n5928 16
R17558 VSS.n5974 VSS.n5973 16
R17559 VSS.n5973 VSS.n5972 16
R17560 VSS.n5972 VSS.n5970 16
R17561 VSS.n5970 VSS.n5967 16
R17562 VSS.n5967 VSS.n5966 16
R17563 VSS.n5966 VSS.n5963 16
R17564 VSS.n5963 VSS.n5962 16
R17565 VSS.n6051 VSS.n6033 16
R17566 VSS.n6052 VSS.n6051 16
R17567 VSS.n6055 VSS.n6052 16
R17568 VSS.n6056 VSS.n6055 16
R17569 VSS.n6059 VSS.n6056 16
R17570 VSS.n6060 VSS.n6059 16
R17571 VSS.n6063 VSS.n6060 16
R17572 VSS.n6065 VSS.n6063 16
R17573 VSS.n6081 VSS.n6080 16
R17574 VSS.n6080 VSS.n6077 16
R17575 VSS.n6077 VSS.n6076 16
R17576 VSS.n6076 VSS.n6073 16
R17577 VSS.n6073 VSS.n6072 16
R17578 VSS.n6072 VSS.n6069 16
R17579 VSS.n6069 VSS.n6068 16
R17580 VSS.n6068 VSS.n6066 16
R17581 VSS.n6096 VSS.n6050 16
R17582 VSS.n6096 VSS.n6095 16
R17583 VSS.n6095 VSS.n6094 16
R17584 VSS.n6094 VSS.n6092 16
R17585 VSS.n6092 VSS.n6089 16
R17586 VSS.n6089 VSS.n6088 16
R17587 VSS.n6088 VSS.n6085 16
R17588 VSS.n6085 VSS.n6084 16
R17589 VSS.n6173 VSS.n6155 16
R17590 VSS.n6174 VSS.n6173 16
R17591 VSS.n6177 VSS.n6174 16
R17592 VSS.n6178 VSS.n6177 16
R17593 VSS.n6181 VSS.n6178 16
R17594 VSS.n6182 VSS.n6181 16
R17595 VSS.n6185 VSS.n6182 16
R17596 VSS.n6187 VSS.n6185 16
R17597 VSS.n6203 VSS.n6202 16
R17598 VSS.n6202 VSS.n6199 16
R17599 VSS.n6199 VSS.n6198 16
R17600 VSS.n6198 VSS.n6195 16
R17601 VSS.n6195 VSS.n6194 16
R17602 VSS.n6194 VSS.n6191 16
R17603 VSS.n6191 VSS.n6190 16
R17604 VSS.n6190 VSS.n6188 16
R17605 VSS.n6218 VSS.n6172 16
R17606 VSS.n6218 VSS.n6217 16
R17607 VSS.n6217 VSS.n6216 16
R17608 VSS.n6216 VSS.n6214 16
R17609 VSS.n6214 VSS.n6211 16
R17610 VSS.n6211 VSS.n6210 16
R17611 VSS.n6210 VSS.n6207 16
R17612 VSS.n6207 VSS.n6206 16
R17613 VSS.n6295 VSS.n6277 16
R17614 VSS.n6296 VSS.n6295 16
R17615 VSS.n6299 VSS.n6296 16
R17616 VSS.n6300 VSS.n6299 16
R17617 VSS.n6303 VSS.n6300 16
R17618 VSS.n6304 VSS.n6303 16
R17619 VSS.n6307 VSS.n6304 16
R17620 VSS.n6309 VSS.n6307 16
R17621 VSS.n6325 VSS.n6324 16
R17622 VSS.n6324 VSS.n6321 16
R17623 VSS.n6321 VSS.n6320 16
R17624 VSS.n6320 VSS.n6317 16
R17625 VSS.n6317 VSS.n6316 16
R17626 VSS.n6316 VSS.n6313 16
R17627 VSS.n6313 VSS.n6312 16
R17628 VSS.n6312 VSS.n6310 16
R17629 VSS.n6340 VSS.n6294 16
R17630 VSS.n6340 VSS.n6339 16
R17631 VSS.n6339 VSS.n6338 16
R17632 VSS.n6338 VSS.n6336 16
R17633 VSS.n6336 VSS.n6333 16
R17634 VSS.n6333 VSS.n6332 16
R17635 VSS.n6332 VSS.n6329 16
R17636 VSS.n6329 VSS.n6328 16
R17637 VSS.n6417 VSS.n6399 16
R17638 VSS.n6418 VSS.n6417 16
R17639 VSS.n6421 VSS.n6418 16
R17640 VSS.n6422 VSS.n6421 16
R17641 VSS.n6425 VSS.n6422 16
R17642 VSS.n6426 VSS.n6425 16
R17643 VSS.n6429 VSS.n6426 16
R17644 VSS.n6431 VSS.n6429 16
R17645 VSS.n6447 VSS.n6446 16
R17646 VSS.n6446 VSS.n6443 16
R17647 VSS.n6443 VSS.n6442 16
R17648 VSS.n6442 VSS.n6439 16
R17649 VSS.n6439 VSS.n6438 16
R17650 VSS.n6438 VSS.n6435 16
R17651 VSS.n6435 VSS.n6434 16
R17652 VSS.n6434 VSS.n6432 16
R17653 VSS.n6462 VSS.n6416 16
R17654 VSS.n6462 VSS.n6461 16
R17655 VSS.n6461 VSS.n6460 16
R17656 VSS.n6460 VSS.n6458 16
R17657 VSS.n6458 VSS.n6455 16
R17658 VSS.n6455 VSS.n6454 16
R17659 VSS.n6454 VSS.n6451 16
R17660 VSS.n6451 VSS.n6450 16
R17661 VSS.n6589 VSS.n6588 16
R17662 VSS.n6588 VSS.n6520 16
R17663 VSS.n6583 VSS.n6520 16
R17664 VSS.n6583 VSS.n6582 16
R17665 VSS.n6582 VSS.n6522 16
R17666 VSS.n6577 VSS.n6522 16
R17667 VSS.n6577 VSS.n6576 16
R17668 VSS.n6576 VSS.n6575 16
R17669 VSS.n6560 VSS.n6559 16
R17670 VSS.n6561 VSS.n6560 16
R17671 VSS.n6561 VSS.n6528 16
R17672 VSS.n6567 VSS.n6528 16
R17673 VSS.n6568 VSS.n6567 16
R17674 VSS.n6569 VSS.n6568 16
R17675 VSS.n6569 VSS.n6526 16
R17676 VSS.n6574 VSS.n6526 16
R17677 VSS.n6543 VSS.n6539 16
R17678 VSS.n6544 VSS.n6543 16
R17679 VSS.n6545 VSS.n6544 16
R17680 VSS.n6545 VSS.n6532 16
R17681 VSS.n6551 VSS.n6532 16
R17682 VSS.n6552 VSS.n6551 16
R17683 VSS.n6553 VSS.n6552 16
R17684 VSS.n6553 VSS.n6530 16
R17685 VSS.n46 VSS.n3 16
R17686 VSS.n47 VSS.n46 16
R17687 VSS.n50 VSS.n47 16
R17688 VSS.n51 VSS.n50 16
R17689 VSS.n54 VSS.n51 16
R17690 VSS.n55 VSS.n54 16
R17691 VSS.n58 VSS.n55 16
R17692 VSS.n60 VSS.n58 16
R17693 VSS.n76 VSS.n75 16
R17694 VSS.n75 VSS.n72 16
R17695 VSS.n72 VSS.n71 16
R17696 VSS.n71 VSS.n68 16
R17697 VSS.n68 VSS.n67 16
R17698 VSS.n67 VSS.n64 16
R17699 VSS.n64 VSS.n63 16
R17700 VSS.n63 VSS.n61 16
R17701 VSS.n94 VSS.n93 16
R17702 VSS.n93 VSS.n91 16
R17703 VSS.n91 VSS.n88 16
R17704 VSS.n88 VSS.n87 16
R17705 VSS.n87 VSS.n84 16
R17706 VSS.n84 VSS.n83 16
R17707 VSS.n83 VSS.n80 16
R17708 VSS.n80 VSS.n79 16
R17709 VSS.n1171 VSS.n97 16
R17710 VSS.n137 VSS.n97 16
R17711 VSS.n140 VSS.n137 16
R17712 VSS.n141 VSS.n140 16
R17713 VSS.n144 VSS.n141 16
R17714 VSS.n145 VSS.n144 16
R17715 VSS.n148 VSS.n145 16
R17716 VSS.n150 VSS.n148 16
R17717 VSS.n166 VSS.n165 16
R17718 VSS.n165 VSS.n162 16
R17719 VSS.n162 VSS.n161 16
R17720 VSS.n161 VSS.n158 16
R17721 VSS.n158 VSS.n157 16
R17722 VSS.n157 VSS.n154 16
R17723 VSS.n154 VSS.n153 16
R17724 VSS.n153 VSS.n151 16
R17725 VSS.n184 VSS.n183 16
R17726 VSS.n183 VSS.n181 16
R17727 VSS.n181 VSS.n178 16
R17728 VSS.n178 VSS.n177 16
R17729 VSS.n177 VSS.n174 16
R17730 VSS.n174 VSS.n173 16
R17731 VSS.n173 VSS.n170 16
R17732 VSS.n170 VSS.n169 16
R17733 VSS.n1081 VSS.n187 16
R17734 VSS.n227 VSS.n187 16
R17735 VSS.n230 VSS.n227 16
R17736 VSS.n231 VSS.n230 16
R17737 VSS.n234 VSS.n231 16
R17738 VSS.n235 VSS.n234 16
R17739 VSS.n238 VSS.n235 16
R17740 VSS.n240 VSS.n238 16
R17741 VSS.n256 VSS.n255 16
R17742 VSS.n255 VSS.n252 16
R17743 VSS.n252 VSS.n251 16
R17744 VSS.n251 VSS.n248 16
R17745 VSS.n248 VSS.n247 16
R17746 VSS.n247 VSS.n244 16
R17747 VSS.n244 VSS.n243 16
R17748 VSS.n243 VSS.n241 16
R17749 VSS.n274 VSS.n273 16
R17750 VSS.n273 VSS.n271 16
R17751 VSS.n271 VSS.n268 16
R17752 VSS.n268 VSS.n267 16
R17753 VSS.n267 VSS.n264 16
R17754 VSS.n264 VSS.n263 16
R17755 VSS.n263 VSS.n260 16
R17756 VSS.n260 VSS.n259 16
R17757 VSS.n991 VSS.n277 16
R17758 VSS.n317 VSS.n277 16
R17759 VSS.n320 VSS.n317 16
R17760 VSS.n321 VSS.n320 16
R17761 VSS.n324 VSS.n321 16
R17762 VSS.n325 VSS.n324 16
R17763 VSS.n328 VSS.n325 16
R17764 VSS.n330 VSS.n328 16
R17765 VSS.n346 VSS.n345 16
R17766 VSS.n345 VSS.n342 16
R17767 VSS.n342 VSS.n341 16
R17768 VSS.n341 VSS.n338 16
R17769 VSS.n338 VSS.n337 16
R17770 VSS.n337 VSS.n334 16
R17771 VSS.n334 VSS.n333 16
R17772 VSS.n333 VSS.n331 16
R17773 VSS.n364 VSS.n363 16
R17774 VSS.n363 VSS.n361 16
R17775 VSS.n361 VSS.n358 16
R17776 VSS.n358 VSS.n357 16
R17777 VSS.n357 VSS.n354 16
R17778 VSS.n354 VSS.n353 16
R17779 VSS.n353 VSS.n350 16
R17780 VSS.n350 VSS.n349 16
R17781 VSS.n901 VSS.n367 16
R17782 VSS.n407 VSS.n367 16
R17783 VSS.n410 VSS.n407 16
R17784 VSS.n411 VSS.n410 16
R17785 VSS.n414 VSS.n411 16
R17786 VSS.n415 VSS.n414 16
R17787 VSS.n418 VSS.n415 16
R17788 VSS.n420 VSS.n418 16
R17789 VSS.n436 VSS.n435 16
R17790 VSS.n435 VSS.n432 16
R17791 VSS.n432 VSS.n431 16
R17792 VSS.n431 VSS.n428 16
R17793 VSS.n428 VSS.n427 16
R17794 VSS.n427 VSS.n424 16
R17795 VSS.n424 VSS.n423 16
R17796 VSS.n423 VSS.n421 16
R17797 VSS.n454 VSS.n453 16
R17798 VSS.n453 VSS.n451 16
R17799 VSS.n451 VSS.n448 16
R17800 VSS.n448 VSS.n447 16
R17801 VSS.n447 VSS.n444 16
R17802 VSS.n444 VSS.n443 16
R17803 VSS.n443 VSS.n440 16
R17804 VSS.n440 VSS.n439 16
R17805 VSS.n811 VSS.n457 16
R17806 VSS.n497 VSS.n457 16
R17807 VSS.n500 VSS.n497 16
R17808 VSS.n501 VSS.n500 16
R17809 VSS.n504 VSS.n501 16
R17810 VSS.n505 VSS.n504 16
R17811 VSS.n508 VSS.n505 16
R17812 VSS.n510 VSS.n508 16
R17813 VSS.n526 VSS.n525 16
R17814 VSS.n525 VSS.n522 16
R17815 VSS.n522 VSS.n521 16
R17816 VSS.n521 VSS.n518 16
R17817 VSS.n518 VSS.n517 16
R17818 VSS.n517 VSS.n514 16
R17819 VSS.n514 VSS.n513 16
R17820 VSS.n513 VSS.n511 16
R17821 VSS.n544 VSS.n543 16
R17822 VSS.n543 VSS.n541 16
R17823 VSS.n541 VSS.n538 16
R17824 VSS.n538 VSS.n537 16
R17825 VSS.n537 VSS.n534 16
R17826 VSS.n534 VSS.n533 16
R17827 VSS.n533 VSS.n530 16
R17828 VSS.n530 VSS.n529 16
R17829 VSS.n721 VSS.n547 16
R17830 VSS.n587 VSS.n547 16
R17831 VSS.n590 VSS.n587 16
R17832 VSS.n591 VSS.n590 16
R17833 VSS.n594 VSS.n591 16
R17834 VSS.n595 VSS.n594 16
R17835 VSS.n598 VSS.n595 16
R17836 VSS.n600 VSS.n598 16
R17837 VSS.n616 VSS.n615 16
R17838 VSS.n615 VSS.n612 16
R17839 VSS.n612 VSS.n611 16
R17840 VSS.n611 VSS.n608 16
R17841 VSS.n608 VSS.n607 16
R17842 VSS.n607 VSS.n604 16
R17843 VSS.n604 VSS.n603 16
R17844 VSS.n603 VSS.n601 16
R17845 VSS.n634 VSS.n633 16
R17846 VSS.n633 VSS.n631 16
R17847 VSS.n631 VSS.n628 16
R17848 VSS.n628 VSS.n627 16
R17849 VSS.n627 VSS.n624 16
R17850 VSS.n624 VSS.n623 16
R17851 VSS.n623 VSS.n620 16
R17852 VSS.n620 VSS.n619 16
R17853 VSS.n17334 VSS.n17331 14.755
R17854 VSS.n17309 VSS.n16053 14.755
R17855 VSS.n17219 VSS.n16143 14.755
R17856 VSS.n17129 VSS.n16233 14.755
R17857 VSS.n17039 VSS.n16323 14.755
R17858 VSS.n16949 VSS.n16413 14.755
R17859 VSS.n16859 VSS.n16503 14.755
R17860 VSS.n16769 VSS.n16593 14.755
R17861 VSS.n11236 VSS.n11060 14.755
R17862 VSS.n11326 VSS.n10970 14.755
R17863 VSS.n11416 VSS.n10880 14.755
R17864 VSS.n13536 VSS.n10790 14.755
R17865 VSS.n13626 VSS.n10700 14.755
R17866 VSS.n13716 VSS.n10610 14.755
R17867 VSS.n13806 VSS.n10520 14.755
R17868 VSS.n13834 VSS.n13828 14.755
R17869 VSS.n9149 VSS.n9148 14.755
R17870 VSS.n10264 VSS.n9188 14.755
R17871 VSS.n10174 VSS.n9278 14.755
R17872 VSS.n10084 VSS.n9368 14.755
R17873 VSS.n9994 VSS.n9458 14.755
R17874 VSS.n9904 VSS.n9548 14.755
R17875 VSS.n9814 VSS.n9638 14.755
R17876 VSS.n9162 VSS.n8978 14.755
R17877 VSS.n5666 VSS.n3632 14.755
R17878 VSS.n5788 VSS.n3574 14.755
R17879 VSS.n5910 VSS.n3516 14.755
R17880 VSS.n6032 VSS.n3458 14.755
R17881 VSS.n6154 VSS.n3400 14.755
R17882 VSS.n6276 VSS.n3342 14.755
R17883 VSS.n6398 VSS.n3284 14.755
R17884 VSS.n6591 VSS.n6590 14.755
R17885 VSS.n1172 VSS.n96 14.755
R17886 VSS.n1082 VSS.n186 14.755
R17887 VSS.n992 VSS.n276 14.755
R17888 VSS.n902 VSS.n366 14.755
R17889 VSS.n812 VSS.n456 14.755
R17890 VSS.n722 VSS.n546 14.755
R17891 VSS.n17304 VSS.n16075 14.615
R17892 VSS.n17214 VSS.n16165 14.615
R17893 VSS.n17124 VSS.n16255 14.615
R17894 VSS.n17034 VSS.n16345 14.615
R17895 VSS.n16944 VSS.n16435 14.615
R17896 VSS.n16854 VSS.n16525 14.615
R17897 VSS.n16764 VSS.n16615 14.615
R17898 VSS.n10259 VSS.n9210 14.615
R17899 VSS.n10169 VSS.n9300 14.615
R17900 VSS.n10079 VSS.n9390 14.615
R17901 VSS.n9989 VSS.n9480 14.615
R17902 VSS.n9899 VSS.n9570 14.615
R17903 VSS.n9809 VSS.n9660 14.615
R17904 VSS.n8977 VSS.n8971 14.615
R17905 VSS.n3630 VSS.n3624 14.615
R17906 VSS.n3572 VSS.n3566 14.615
R17907 VSS.n3514 VSS.n3508 14.615
R17908 VSS.n3456 VSS.n3450 14.615
R17909 VSS.n3398 VSS.n3392 14.615
R17910 VSS.n3340 VSS.n3334 14.615
R17911 VSS.n3282 VSS.n3276 14.615
R17912 VSS.n6597 VSS.n3157 14.615
R17913 VSS.n27 VSS.n7 14.615
R17914 VSS.n1167 VSS.n118 14.615
R17915 VSS.n1077 VSS.n208 14.615
R17916 VSS.n987 VSS.n298 14.615
R17917 VSS.n897 VSS.n388 14.615
R17918 VSS.n807 VSS.n478 14.615
R17919 VSS.n717 VSS.n568 14.615
R17920 VSS.n6728 VSS.n6727 13.866
R17921 VSS.n6700 sky130_asc_pnp_05v5_W3p40L3p40_1_0/Base 13.688
R17922 VSS.n6728 VSS.n6635 13.688
R17923 VSS.n14723 VSS.n14366 13.653
R17924 VSS.n14715 VSS.n14370 13.653
R17925 VSS.n14707 VSS.n14380 13.653
R17926 VSS.n14388 VSS.n14382 13.653
R17927 VSS.n14692 VSS.n14389 13.653
R17928 VSS.n14684 VSS.n14399 13.653
R17929 VSS.n14407 VSS.n14401 13.653
R17930 VSS.n14670 VSS.n14408 13.653
R17931 VSS.n14662 VSS.n14418 13.653
R17932 VSS.n14426 VSS.n14420 13.653
R17933 VSS.n14647 VSS.n14427 13.653
R17934 VSS.n14639 VSS.n14437 13.653
R17935 VSS.n14876 VSS.n14300 13.653
R17936 VSS.n14884 VSS.n14294 13.653
R17937 VSS.n14896 VSS.n14289 13.653
R17938 VSS.n14900 VSS.n14281 13.653
R17939 VSS.n14911 VSS.n14279 13.653
R17940 VSS.n14919 VSS.n14273 13.653
R17941 VSS.n14930 VSS.n14268 13.653
R17942 VSS.n14934 VSS.n14260 13.653
R17943 VSS.n14945 VSS.n14258 13.653
R17944 VSS.n14953 VSS.n14252 13.653
R17945 VSS.n14965 VSS.n14247 13.653
R17946 VSS.n14969 VSS.n14240 13.653
R17947 VSS.n14481 VSS.n14478 13.653
R17948 VSS.n14623 VSS.n14479 13.653
R17949 VSS.n14615 VSS.n14492 13.653
R17950 VSS.n14500 VSS.n14494 13.653
R17951 VSS.n14600 VSS.n14501 13.653
R17952 VSS.n14592 VSS.n14511 13.653
R17953 VSS.n14519 VSS.n14513 13.653
R17954 VSS.n14578 VSS.n14520 13.653
R17955 VSS.n14570 VSS.n14530 13.653
R17956 VSS.n14538 VSS.n14532 13.653
R17957 VSS.n14555 VSS.n14539 13.653
R17958 VSS.n14545 VSS.n14303 13.653
R17959 VSS.n15090 VSS.n15087 13.653
R17960 VSS.n15224 VSS.n15088 13.653
R17961 VSS.n15216 VSS.n15101 13.653
R17962 VSS.n15109 VSS.n15103 13.653
R17963 VSS.n15201 VSS.n15110 13.653
R17964 VSS.n15193 VSS.n15120 13.653
R17965 VSS.n15128 VSS.n15122 13.653
R17966 VSS.n15179 VSS.n15129 13.653
R17967 VSS.n15171 VSS.n15139 13.653
R17968 VSS.n15147 VSS.n15141 13.653
R17969 VSS.n15156 VSS.n15148 13.653
R17970 VSS.n15446 VSS.n14142 13.653
R17971 VSS.n14978 VSS.n14977 13.653
R17972 VSS.n15316 VSS.n14979 13.653
R17973 VSS.n15308 VSS.n14989 13.653
R17974 VSS.n14997 VSS.n14991 13.653
R17975 VSS.n15293 VSS.n14998 13.653
R17976 VSS.n15285 VSS.n15008 13.653
R17977 VSS.n15016 VSS.n15010 13.653
R17978 VSS.n15271 VSS.n15017 13.653
R17979 VSS.n15263 VSS.n15027 13.653
R17980 VSS.n15035 VSS.n15029 13.653
R17981 VSS.n15248 VSS.n15036 13.653
R17982 VSS.n15240 VSS.n15046 13.653
R17983 VSS.n15565 VSS.n15563 13.653
R17984 VSS.n15883 VSS.n15564 13.653
R17985 VSS.n15875 VSS.n15576 13.653
R17986 VSS.n15584 VSS.n15578 13.653
R17987 VSS.n15860 VSS.n15585 13.653
R17988 VSS.n15852 VSS.n15595 13.653
R17989 VSS.n15603 VSS.n15597 13.653
R17990 VSS.n15838 VSS.n15604 13.653
R17991 VSS.n15830 VSS.n15614 13.653
R17992 VSS.n15622 VSS.n15616 13.653
R17993 VSS.n15815 VSS.n15623 13.653
R17994 VSS.n15807 VSS.n15633 13.653
R17995 VSS.n15459 VSS.n14133 13.653
R17996 VSS.n15463 VSS.n14125 13.653
R17997 VSS.n15474 VSS.n14123 13.653
R17998 VSS.n15482 VSS.n14117 13.653
R17999 VSS.n15494 VSS.n14112 13.653
R18000 VSS.n15498 VSS.n14104 13.653
R18001 VSS.n15509 VSS.n14102 13.653
R18002 VSS.n15516 VSS.n14096 13.653
R18003 VSS.n15528 VSS.n14091 13.653
R18004 VSS.n15532 VSS.n14083 13.653
R18005 VSS.n15543 VSS.n14081 13.653
R18006 VSS.n15551 VSS.n14075 13.653
R18007 VSS.n15677 VSS.n15674 13.653
R18008 VSS.n15791 VSS.n15675 13.653
R18009 VSS.n15783 VSS.n15688 13.653
R18010 VSS.n15696 VSS.n15690 13.653
R18011 VSS.n15768 VSS.n15697 13.653
R18012 VSS.n15760 VSS.n15707 13.653
R18013 VSS.n15715 VSS.n15709 13.653
R18014 VSS.n15746 VSS.n15716 13.653
R18015 VSS.n15738 VSS.n15726 13.653
R18016 VSS.n15728 VSS.n13999 13.653
R18017 VSS.n16016 VSS.n14000 13.653
R18018 VSS.n16008 VSS.n14010 13.653
R18019 VSS.n12794 VSS.n12721 13.653
R18020 VSS.n12806 VSS.n12716 13.653
R18021 VSS.n12810 VSS.n12708 13.653
R18022 VSS.n12821 VSS.n12706 13.653
R18023 VSS.n12829 VSS.n12700 13.653
R18024 VSS.n12841 VSS.n12695 13.653
R18025 VSS.n12845 VSS.n12687 13.653
R18026 VSS.n12855 VSS.n12685 13.653
R18027 VSS.n12863 VSS.n12679 13.653
R18028 VSS.n12875 VSS.n12674 13.653
R18029 VSS.n12880 VSS.n12672 13.653
R18030 VSS.n12889 VSS.n12663 13.653
R18031 VSS.n13151 VSS.n12580 13.653
R18032 VSS.n13163 VSS.n12575 13.653
R18033 VSS.n13167 VSS.n12567 13.653
R18034 VSS.n13178 VSS.n12565 13.653
R18035 VSS.n13186 VSS.n12559 13.653
R18036 VSS.n13198 VSS.n12554 13.653
R18037 VSS.n13202 VSS.n12546 13.653
R18038 VSS.n13212 VSS.n12544 13.653
R18039 VSS.n13220 VSS.n12538 13.653
R18040 VSS.n13232 VSS.n12533 13.653
R18041 VSS.n13237 VSS.n12531 13.653
R18042 VSS.n13246 VSS.n12522 13.653
R18043 VSS.n13055 VSS.n13054 13.653
R18044 VSS.n13046 VSS.n12897 13.653
R18045 VSS.n12906 VSS.n12900 13.653
R18046 VSS.n13031 VSS.n12907 13.653
R18047 VSS.n13023 VSS.n12917 13.653
R18048 VSS.n12925 VSS.n12919 13.653
R18049 VSS.n13008 VSS.n12926 13.653
R18050 VSS.n13001 VSS.n12936 13.653
R18051 VSS.n12944 VSS.n12938 13.653
R18052 VSS.n12986 VSS.n12945 13.653
R18053 VSS.n12978 VSS.n12955 13.653
R18054 VSS.n12964 VSS.n12957 13.653
R18055 VSS.n11672 VSS.n11671 13.653
R18056 VSS.n11684 VSS.n11666 13.653
R18057 VSS.n11688 VSS.n11658 13.653
R18058 VSS.n11699 VSS.n11656 13.653
R18059 VSS.n11707 VSS.n11650 13.653
R18060 VSS.n11719 VSS.n11645 13.653
R18061 VSS.n11723 VSS.n11637 13.653
R18062 VSS.n11733 VSS.n11635 13.653
R18063 VSS.n11741 VSS.n11629 13.653
R18064 VSS.n11753 VSS.n11624 13.653
R18065 VSS.n11757 VSS.n11615 13.653
R18066 VSS.n11768 VSS.n11613 13.653
R18067 VSS.n13304 VSS.n13303 13.653
R18068 VSS.n13295 VSS.n13254 13.653
R18069 VSS.n13263 VSS.n13257 13.653
R18070 VSS.n13280 VSS.n13264 13.653
R18071 VSS.n13270 VSS.n11433 13.653
R18072 VSS.n13450 VSS.n11434 13.653
R18073 VSS.n13442 VSS.n11444 13.653
R18074 VSS.n11452 VSS.n11446 13.653
R18075 VSS.n13428 VSS.n11453 13.653
R18076 VSS.n13420 VSS.n11463 13.653
R18077 VSS.n11471 VSS.n11465 13.653
R18078 VSS.n13405 VSS.n11472 13.653
R18079 VSS.n11912 VSS.n11911 13.653
R18080 VSS.n12391 VSS.n11913 13.653
R18081 VSS.n12383 VSS.n11923 13.653
R18082 VSS.n11931 VSS.n11925 13.653
R18083 VSS.n12368 VSS.n11932 13.653
R18084 VSS.n12360 VSS.n11942 13.653
R18085 VSS.n11950 VSS.n11944 13.653
R18086 VSS.n12346 VSS.n11951 13.653
R18087 VSS.n12338 VSS.n11961 13.653
R18088 VSS.n11969 VSS.n11963 13.653
R18089 VSS.n12323 VSS.n11970 13.653
R18090 VSS.n12315 VSS.n11980 13.653
R18091 VSS.n11810 VSS.n11605 13.653
R18092 VSS.n11818 VSS.n11599 13.653
R18093 VSS.n11830 VSS.n11594 13.653
R18094 VSS.n11834 VSS.n11586 13.653
R18095 VSS.n11845 VSS.n11584 13.653
R18096 VSS.n11853 VSS.n11578 13.653
R18097 VSS.n11864 VSS.n11573 13.653
R18098 VSS.n11868 VSS.n11565 13.653
R18099 VSS.n11879 VSS.n11563 13.653
R18100 VSS.n11887 VSS.n11557 13.653
R18101 VSS.n11899 VSS.n11552 13.653
R18102 VSS.n11903 VSS.n11545 13.653
R18103 VSS.n11991 VSS.n11988 13.653
R18104 VSS.n12299 VSS.n11989 13.653
R18105 VSS.n12291 VSS.n12002 13.653
R18106 VSS.n12010 VSS.n12004 13.653
R18107 VSS.n12276 VSS.n12011 13.653
R18108 VSS.n12268 VSS.n12021 13.653
R18109 VSS.n12029 VSS.n12023 13.653
R18110 VSS.n12254 VSS.n12030 13.653
R18111 VSS.n12246 VSS.n12040 13.653
R18112 VSS.n12048 VSS.n12042 13.653
R18113 VSS.n12231 VSS.n12049 13.653
R18114 VSS.n12223 VSS.n12059 13.653
R18115 VSS.n7837 VSS.n7674 13.653
R18116 VSS.n7829 VSS.n7677 13.653
R18117 VSS.n7821 VSS.n7687 13.653
R18118 VSS.n7695 VSS.n7689 13.653
R18119 VSS.n7806 VSS.n7696 13.653
R18120 VSS.n7798 VSS.n7706 13.653
R18121 VSS.n7714 VSS.n7708 13.653
R18122 VSS.n7784 VSS.n7715 13.653
R18123 VSS.n7776 VSS.n7725 13.653
R18124 VSS.n7733 VSS.n7727 13.653
R18125 VSS.n7761 VSS.n7734 13.653
R18126 VSS.n7753 VSS.n7750 13.653
R18127 VSS.n8182 VSS.n8181 13.653
R18128 VSS.n8177 VSS.n8022 13.653
R18129 VSS.n8169 VSS.n8031 13.653
R18130 VSS.n8161 VSS.n8041 13.653
R18131 VSS.n8049 VSS.n8043 13.653
R18132 VSS.n8146 VSS.n8050 13.653
R18133 VSS.n8138 VSS.n8060 13.653
R18134 VSS.n8068 VSS.n8062 13.653
R18135 VSS.n8124 VSS.n8069 13.653
R18136 VSS.n8116 VSS.n8079 13.653
R18137 VSS.n8087 VSS.n8081 13.653
R18138 VSS.n8101 VSS.n8088 13.653
R18139 VSS.n7921 VSS.n7599 13.653
R18140 VSS.n7929 VSS.n7593 13.653
R18141 VSS.n7941 VSS.n7588 13.653
R18142 VSS.n7945 VSS.n7580 13.653
R18143 VSS.n7956 VSS.n7578 13.653
R18144 VSS.n7964 VSS.n7572 13.653
R18145 VSS.n7975 VSS.n7567 13.653
R18146 VSS.n7979 VSS.n7559 13.653
R18147 VSS.n7990 VSS.n7557 13.653
R18148 VSS.n7998 VSS.n7551 13.653
R18149 VSS.n8010 VSS.n7546 13.653
R18150 VSS.n8014 VSS.n7538 13.653
R18151 VSS.n8540 VSS.n8539 13.653
R18152 VSS.n8535 VSS.n8380 13.653
R18153 VSS.n8527 VSS.n8389 13.653
R18154 VSS.n8519 VSS.n8399 13.653
R18155 VSS.n8407 VSS.n8401 13.653
R18156 VSS.n8504 VSS.n8408 13.653
R18157 VSS.n8496 VSS.n8418 13.653
R18158 VSS.n8426 VSS.n8420 13.653
R18159 VSS.n8482 VSS.n8427 13.653
R18160 VSS.n8474 VSS.n8437 13.653
R18161 VSS.n8445 VSS.n8439 13.653
R18162 VSS.n8459 VSS.n8446 13.653
R18163 VSS.n8279 VSS.n7459 13.653
R18164 VSS.n8287 VSS.n7453 13.653
R18165 VSS.n8299 VSS.n7448 13.653
R18166 VSS.n8303 VSS.n7440 13.653
R18167 VSS.n8314 VSS.n7438 13.653
R18168 VSS.n8322 VSS.n7432 13.653
R18169 VSS.n8333 VSS.n7427 13.653
R18170 VSS.n8337 VSS.n7419 13.653
R18171 VSS.n8348 VSS.n7417 13.653
R18172 VSS.n8356 VSS.n7411 13.653
R18173 VSS.n8368 VSS.n7406 13.653
R18174 VSS.n8372 VSS.n7398 13.653
R18175 VSS.n8762 VSS.n8761 13.653
R18176 VSS.n8757 VSS.n8738 13.653
R18177 VSS.n8750 VSS.n6905 13.653
R18178 VSS.n8922 VSS.n6906 13.653
R18179 VSS.n8914 VSS.n6916 13.653
R18180 VSS.n6924 VSS.n6918 13.653
R18181 VSS.n8899 VSS.n6925 13.653
R18182 VSS.n8892 VSS.n6935 13.653
R18183 VSS.n6943 VSS.n6937 13.653
R18184 VSS.n8877 VSS.n6944 13.653
R18185 VSS.n8869 VSS.n6954 13.653
R18186 VSS.n6962 VSS.n6956 13.653
R18187 VSS.n8637 VSS.n7319 13.653
R18188 VSS.n8645 VSS.n7313 13.653
R18189 VSS.n8657 VSS.n7308 13.653
R18190 VSS.n8661 VSS.n7300 13.653
R18191 VSS.n8672 VSS.n7298 13.653
R18192 VSS.n8680 VSS.n7292 13.653
R18193 VSS.n8691 VSS.n7287 13.653
R18194 VSS.n8695 VSS.n7279 13.653
R18195 VSS.n8706 VSS.n7277 13.653
R18196 VSS.n8714 VSS.n7271 13.653
R18197 VSS.n8726 VSS.n7266 13.653
R18198 VSS.n8730 VSS.n7258 13.653
R18199 VSS.n7075 VSS.n7067 13.653
R18200 VSS.n7079 VSS.n7060 13.653
R18201 VSS.n7090 VSS.n7058 13.653
R18202 VSS.n7098 VSS.n7052 13.653
R18203 VSS.n7110 VSS.n7047 13.653
R18204 VSS.n7114 VSS.n7039 13.653
R18205 VSS.n7125 VSS.n7037 13.653
R18206 VSS.n7132 VSS.n7031 13.653
R18207 VSS.n7144 VSS.n7026 13.653
R18208 VSS.n7148 VSS.n7018 13.653
R18209 VSS.n7159 VSS.n7016 13.653
R18210 VSS.n7167 VSS.n7009 13.653
R18211 VSS.n4247 VSS.n4174 13.653
R18212 VSS.n4259 VSS.n4169 13.653
R18213 VSS.n4263 VSS.n4161 13.653
R18214 VSS.n4274 VSS.n4159 13.653
R18215 VSS.n4282 VSS.n4153 13.653
R18216 VSS.n4294 VSS.n4148 13.653
R18217 VSS.n4298 VSS.n4140 13.653
R18218 VSS.n4308 VSS.n4138 13.653
R18219 VSS.n4316 VSS.n4132 13.653
R18220 VSS.n4328 VSS.n4127 13.653
R18221 VSS.n4333 VSS.n4125 13.653
R18222 VSS.n4342 VSS.n4116 13.653
R18223 VSS.n4604 VSS.n4033 13.653
R18224 VSS.n4616 VSS.n4028 13.653
R18225 VSS.n4620 VSS.n4020 13.653
R18226 VSS.n4631 VSS.n4018 13.653
R18227 VSS.n4639 VSS.n4012 13.653
R18228 VSS.n4651 VSS.n4007 13.653
R18229 VSS.n4655 VSS.n3999 13.653
R18230 VSS.n4665 VSS.n3997 13.653
R18231 VSS.n4673 VSS.n3991 13.653
R18232 VSS.n4685 VSS.n3986 13.653
R18233 VSS.n4690 VSS.n3984 13.653
R18234 VSS.n4699 VSS.n3975 13.653
R18235 VSS.n4508 VSS.n4507 13.653
R18236 VSS.n4499 VSS.n4350 13.653
R18237 VSS.n4359 VSS.n4353 13.653
R18238 VSS.n4484 VSS.n4360 13.653
R18239 VSS.n4476 VSS.n4370 13.653
R18240 VSS.n4378 VSS.n4372 13.653
R18241 VSS.n4461 VSS.n4379 13.653
R18242 VSS.n4454 VSS.n4389 13.653
R18243 VSS.n4397 VSS.n4391 13.653
R18244 VSS.n4439 VSS.n4398 13.653
R18245 VSS.n4431 VSS.n4408 13.653
R18246 VSS.n4417 VSS.n4410 13.653
R18247 VSS.n4961 VSS.n3892 13.653
R18248 VSS.n4973 VSS.n3887 13.653
R18249 VSS.n4977 VSS.n3879 13.653
R18250 VSS.n4988 VSS.n3877 13.653
R18251 VSS.n4996 VSS.n3871 13.653
R18252 VSS.n5008 VSS.n3866 13.653
R18253 VSS.n5012 VSS.n3858 13.653
R18254 VSS.n5022 VSS.n3856 13.653
R18255 VSS.n5030 VSS.n3850 13.653
R18256 VSS.n5042 VSS.n3845 13.653
R18257 VSS.n5047 VSS.n3843 13.653
R18258 VSS.n5056 VSS.n3834 13.653
R18259 VSS.n4865 VSS.n4864 13.653
R18260 VSS.n4856 VSS.n4707 13.653
R18261 VSS.n4716 VSS.n4710 13.653
R18262 VSS.n4841 VSS.n4717 13.653
R18263 VSS.n4833 VSS.n4727 13.653
R18264 VSS.n4735 VSS.n4729 13.653
R18265 VSS.n4818 VSS.n4736 13.653
R18266 VSS.n4811 VSS.n4746 13.653
R18267 VSS.n4754 VSS.n4748 13.653
R18268 VSS.n4796 VSS.n4755 13.653
R18269 VSS.n4788 VSS.n4765 13.653
R18270 VSS.n4774 VSS.n4767 13.653
R18271 VSS.n5318 VSS.n3751 13.653
R18272 VSS.n5330 VSS.n3746 13.653
R18273 VSS.n5334 VSS.n3738 13.653
R18274 VSS.n5345 VSS.n3736 13.653
R18275 VSS.n5353 VSS.n3730 13.653
R18276 VSS.n5365 VSS.n3725 13.653
R18277 VSS.n5369 VSS.n3717 13.653
R18278 VSS.n5379 VSS.n3715 13.653
R18279 VSS.n5387 VSS.n3709 13.653
R18280 VSS.n5399 VSS.n3704 13.653
R18281 VSS.n5404 VSS.n3702 13.653
R18282 VSS.n5413 VSS.n3693 13.653
R18283 VSS.n5222 VSS.n5221 13.653
R18284 VSS.n5213 VSS.n5064 13.653
R18285 VSS.n5073 VSS.n5067 13.653
R18286 VSS.n5198 VSS.n5074 13.653
R18287 VSS.n5190 VSS.n5084 13.653
R18288 VSS.n5092 VSS.n5086 13.653
R18289 VSS.n5175 VSS.n5093 13.653
R18290 VSS.n5168 VSS.n5103 13.653
R18291 VSS.n5111 VSS.n5105 13.653
R18292 VSS.n5153 VSS.n5112 13.653
R18293 VSS.n5145 VSS.n5122 13.653
R18294 VSS.n5131 VSS.n5124 13.653
R18295 VSS.n5568 VSS.n5567 13.653
R18296 VSS.n5559 VSS.n5421 13.653
R18297 VSS.n5430 VSS.n5424 13.653
R18298 VSS.n5544 VSS.n5431 13.653
R18299 VSS.n5536 VSS.n5441 13.653
R18300 VSS.n5449 VSS.n5443 13.653
R18301 VSS.n5521 VSS.n5450 13.653
R18302 VSS.n5514 VSS.n5460 13.653
R18303 VSS.n5468 VSS.n5462 13.653
R18304 VSS.n5499 VSS.n5469 13.653
R18305 VSS.n5491 VSS.n5479 13.653
R18306 VSS.n5481 VSS.n3639 13.653
R18307 VSS.n1964 VSS.n1607 13.653
R18308 VSS.n1956 VSS.n1611 13.653
R18309 VSS.n1948 VSS.n1621 13.653
R18310 VSS.n1629 VSS.n1623 13.653
R18311 VSS.n1933 VSS.n1630 13.653
R18312 VSS.n1925 VSS.n1640 13.653
R18313 VSS.n1648 VSS.n1642 13.653
R18314 VSS.n1911 VSS.n1649 13.653
R18315 VSS.n1903 VSS.n1659 13.653
R18316 VSS.n1667 VSS.n1661 13.653
R18317 VSS.n1888 VSS.n1668 13.653
R18318 VSS.n1880 VSS.n1678 13.653
R18319 VSS.n2117 VSS.n1541 13.653
R18320 VSS.n2125 VSS.n1535 13.653
R18321 VSS.n2137 VSS.n1530 13.653
R18322 VSS.n2141 VSS.n1522 13.653
R18323 VSS.n2152 VSS.n1520 13.653
R18324 VSS.n2160 VSS.n1514 13.653
R18325 VSS.n2171 VSS.n1509 13.653
R18326 VSS.n2175 VSS.n1501 13.653
R18327 VSS.n2186 VSS.n1499 13.653
R18328 VSS.n2194 VSS.n1493 13.653
R18329 VSS.n2206 VSS.n1488 13.653
R18330 VSS.n2210 VSS.n1481 13.653
R18331 VSS.n1722 VSS.n1719 13.653
R18332 VSS.n1864 VSS.n1720 13.653
R18333 VSS.n1856 VSS.n1733 13.653
R18334 VSS.n1741 VSS.n1735 13.653
R18335 VSS.n1841 VSS.n1742 13.653
R18336 VSS.n1833 VSS.n1752 13.653
R18337 VSS.n1760 VSS.n1754 13.653
R18338 VSS.n1819 VSS.n1761 13.653
R18339 VSS.n1811 VSS.n1771 13.653
R18340 VSS.n1779 VSS.n1773 13.653
R18341 VSS.n1796 VSS.n1780 13.653
R18342 VSS.n1786 VSS.n1544 13.653
R18343 VSS.n2331 VSS.n2328 13.653
R18344 VSS.n2465 VSS.n2329 13.653
R18345 VSS.n2457 VSS.n2342 13.653
R18346 VSS.n2350 VSS.n2344 13.653
R18347 VSS.n2442 VSS.n2351 13.653
R18348 VSS.n2434 VSS.n2361 13.653
R18349 VSS.n2369 VSS.n2363 13.653
R18350 VSS.n2420 VSS.n2370 13.653
R18351 VSS.n2412 VSS.n2380 13.653
R18352 VSS.n2388 VSS.n2382 13.653
R18353 VSS.n2397 VSS.n2389 13.653
R18354 VSS.n2687 VSS.n1383 13.653
R18355 VSS.n2219 VSS.n2218 13.653
R18356 VSS.n2557 VSS.n2220 13.653
R18357 VSS.n2549 VSS.n2230 13.653
R18358 VSS.n2238 VSS.n2232 13.653
R18359 VSS.n2534 VSS.n2239 13.653
R18360 VSS.n2526 VSS.n2249 13.653
R18361 VSS.n2257 VSS.n2251 13.653
R18362 VSS.n2512 VSS.n2258 13.653
R18363 VSS.n2504 VSS.n2268 13.653
R18364 VSS.n2276 VSS.n2270 13.653
R18365 VSS.n2489 VSS.n2277 13.653
R18366 VSS.n2481 VSS.n2287 13.653
R18367 VSS.n2700 VSS.n1374 13.653
R18368 VSS.n2704 VSS.n1366 13.653
R18369 VSS.n2715 VSS.n1364 13.653
R18370 VSS.n2723 VSS.n1358 13.653
R18371 VSS.n2735 VSS.n1353 13.653
R18372 VSS.n2739 VSS.n1345 13.653
R18373 VSS.n2750 VSS.n1343 13.653
R18374 VSS.n2757 VSS.n1337 13.653
R18375 VSS.n2769 VSS.n1332 13.653
R18376 VSS.n2773 VSS.n1324 13.653
R18377 VSS.n2784 VSS.n1322 13.653
R18378 VSS.n2792 VSS.n1316 13.653
R18379 VSS.n2806 VSS.n2804 13.653
R18380 VSS.n2957 VSS.n2805 13.653
R18381 VSS.n2949 VSS.n2817 13.653
R18382 VSS.n2825 VSS.n2819 13.653
R18383 VSS.n2934 VSS.n2826 13.653
R18384 VSS.n2926 VSS.n2836 13.653
R18385 VSS.n2844 VSS.n2838 13.653
R18386 VSS.n2912 VSS.n2845 13.653
R18387 VSS.n2904 VSS.n2855 13.653
R18388 VSS.n2863 VSS.n2857 13.653
R18389 VSS.n2889 VSS.n2864 13.653
R18390 VSS.n2881 VSS.n2878 13.653
R18391 VSS.n1261 VSS.n4 13.511
R18392 VSS.n6825 VSS.n6756 13.058
R18393 VSS.n9155 VSS.n9015 13.014
R18394 VSS.n6704 sky130_asc_pnp_05v5_W3p40L3p40_1_0/xm1/Base 12.977
R18395 VSS.n6801 VSS.n6769 12.412
R18396 sky130_asc_res_xhigh_po_2p85_1_0/VGND sky130_asc_pnp_05v5_W3p40L3p40_8_2/VGND 11.947
R18397 VSS.n17392 VSS.n16034 11.666
R18398 VSS.n17458 VSS.n16037 11.666
R18399 VSS.n17448 VSS.n16033 11.666
R18400 VSS.n17402 VSS.n16038 11.666
R18401 VSS.n17405 VSS.n16032 11.666
R18402 VSS.n17409 VSS.n16039 11.666
R18403 VSS.n17413 VSS.n16031 11.666
R18404 VSS.n17416 VSS.n16029 11.666
R18405 VSS.n17224 VSS.n16082 11.666
R18406 VSS.n17302 VSS.n16076 11.666
R18407 VSS.n17292 VSS.n16073 11.666
R18408 VSS.n17233 VSS.n16077 11.666
R18409 VSS.n17236 VSS.n16072 11.666
R18410 VSS.n17240 VSS.n16078 11.666
R18411 VSS.n17244 VSS.n16071 11.666
R18412 VSS.n17306 VSS.n16079 11.666
R18413 VSS.n17250 VSS.n16075 11.666
R18414 VSS.n17134 VSS.n16172 11.666
R18415 VSS.n17212 VSS.n16166 11.666
R18416 VSS.n17202 VSS.n16163 11.666
R18417 VSS.n17143 VSS.n16167 11.666
R18418 VSS.n17146 VSS.n16162 11.666
R18419 VSS.n17150 VSS.n16168 11.666
R18420 VSS.n17154 VSS.n16161 11.666
R18421 VSS.n17216 VSS.n16169 11.666
R18422 VSS.n17160 VSS.n16165 11.666
R18423 VSS.n17044 VSS.n16262 11.666
R18424 VSS.n17122 VSS.n16256 11.666
R18425 VSS.n17112 VSS.n16253 11.666
R18426 VSS.n17053 VSS.n16257 11.666
R18427 VSS.n17056 VSS.n16252 11.666
R18428 VSS.n17060 VSS.n16258 11.666
R18429 VSS.n17064 VSS.n16251 11.666
R18430 VSS.n17126 VSS.n16259 11.666
R18431 VSS.n17070 VSS.n16255 11.666
R18432 VSS.n16954 VSS.n16352 11.666
R18433 VSS.n17032 VSS.n16346 11.666
R18434 VSS.n17022 VSS.n16343 11.666
R18435 VSS.n16963 VSS.n16347 11.666
R18436 VSS.n16966 VSS.n16342 11.666
R18437 VSS.n16970 VSS.n16348 11.666
R18438 VSS.n16974 VSS.n16341 11.666
R18439 VSS.n17036 VSS.n16349 11.666
R18440 VSS.n16980 VSS.n16345 11.666
R18441 VSS.n16864 VSS.n16442 11.666
R18442 VSS.n16942 VSS.n16436 11.666
R18443 VSS.n16932 VSS.n16433 11.666
R18444 VSS.n16873 VSS.n16437 11.666
R18445 VSS.n16876 VSS.n16432 11.666
R18446 VSS.n16880 VSS.n16438 11.666
R18447 VSS.n16884 VSS.n16431 11.666
R18448 VSS.n16946 VSS.n16439 11.666
R18449 VSS.n16890 VSS.n16435 11.666
R18450 VSS.n16774 VSS.n16532 11.666
R18451 VSS.n16852 VSS.n16526 11.666
R18452 VSS.n16842 VSS.n16523 11.666
R18453 VSS.n16783 VSS.n16527 11.666
R18454 VSS.n16786 VSS.n16522 11.666
R18455 VSS.n16790 VSS.n16528 11.666
R18456 VSS.n16794 VSS.n16521 11.666
R18457 VSS.n16856 VSS.n16529 11.666
R18458 VSS.n16800 VSS.n16525 11.666
R18459 VSS.n16684 VSS.n16622 11.666
R18460 VSS.n16762 VSS.n16616 11.666
R18461 VSS.n16752 VSS.n16613 11.666
R18462 VSS.n16693 VSS.n16617 11.666
R18463 VSS.n16696 VSS.n16612 11.666
R18464 VSS.n16700 VSS.n16618 11.666
R18465 VSS.n16704 VSS.n16611 11.666
R18466 VSS.n16766 VSS.n16619 11.666
R18467 VSS.n16710 VSS.n16615 11.666
R18468 VSS.n11230 VSS.n11080 11.666
R18469 VSS.n11220 VSS.n11084 11.666
R18470 VSS.n11160 VSS.n11079 11.666
R18471 VSS.n11163 VSS.n11085 11.666
R18472 VSS.n11167 VSS.n11078 11.666
R18473 VSS.n11233 VSS.n11086 11.666
R18474 VSS.n11173 VSS.n11082 11.666
R18475 VSS.n11180 VSS.n11179 11.666
R18476 VSS.n11320 VSS.n10990 11.666
R18477 VSS.n11310 VSS.n10994 11.666
R18478 VSS.n11250 VSS.n10989 11.666
R18479 VSS.n11253 VSS.n10995 11.666
R18480 VSS.n11257 VSS.n10988 11.666
R18481 VSS.n11323 VSS.n10996 11.666
R18482 VSS.n11263 VSS.n10992 11.666
R18483 VSS.n11270 VSS.n11269 11.666
R18484 VSS.n11410 VSS.n10900 11.666
R18485 VSS.n11400 VSS.n10904 11.666
R18486 VSS.n11340 VSS.n10899 11.666
R18487 VSS.n11343 VSS.n10905 11.666
R18488 VSS.n11347 VSS.n10898 11.666
R18489 VSS.n11413 VSS.n10906 11.666
R18490 VSS.n11353 VSS.n10902 11.666
R18491 VSS.n11360 VSS.n11359 11.666
R18492 VSS.n13530 VSS.n10810 11.666
R18493 VSS.n13520 VSS.n10814 11.666
R18494 VSS.n13459 VSS.n10809 11.666
R18495 VSS.n13462 VSS.n10815 11.666
R18496 VSS.n13466 VSS.n10808 11.666
R18497 VSS.n13533 VSS.n10816 11.666
R18498 VSS.n13472 VSS.n10812 11.666
R18499 VSS.n13479 VSS.n13478 11.666
R18500 VSS.n13620 VSS.n10720 11.666
R18501 VSS.n13610 VSS.n10724 11.666
R18502 VSS.n13550 VSS.n10719 11.666
R18503 VSS.n13553 VSS.n10725 11.666
R18504 VSS.n13557 VSS.n10718 11.666
R18505 VSS.n13623 VSS.n10726 11.666
R18506 VSS.n13563 VSS.n10722 11.666
R18507 VSS.n13570 VSS.n13569 11.666
R18508 VSS.n13710 VSS.n10630 11.666
R18509 VSS.n13700 VSS.n10634 11.666
R18510 VSS.n13640 VSS.n10629 11.666
R18511 VSS.n13643 VSS.n10635 11.666
R18512 VSS.n13647 VSS.n10628 11.666
R18513 VSS.n13713 VSS.n10636 11.666
R18514 VSS.n13653 VSS.n10632 11.666
R18515 VSS.n13660 VSS.n13659 11.666
R18516 VSS.n13800 VSS.n10540 11.666
R18517 VSS.n13790 VSS.n10544 11.666
R18518 VSS.n13730 VSS.n10539 11.666
R18519 VSS.n13733 VSS.n10545 11.666
R18520 VSS.n13737 VSS.n10538 11.666
R18521 VSS.n13803 VSS.n10546 11.666
R18522 VSS.n13743 VSS.n10542 11.666
R18523 VSS.n13750 VSS.n13749 11.666
R18524 VSS.n13892 VSS.n10503 11.666
R18525 VSS.n13950 VSS.n10505 11.666
R18526 VSS.n13940 VSS.n10502 11.666
R18527 VSS.n13902 VSS.n10506 11.666
R18528 VSS.n13905 VSS.n10501 11.666
R18529 VSS.n13909 VSS.n10507 11.666
R18530 VSS.n13914 VSS.n10500 11.666
R18531 VSS.n13955 VSS.n13954 11.666
R18532 VSS.n9037 VSS.n8989 11.666
R18533 VSS.n9045 VSS.n8988 11.666
R18534 VSS.n9053 VSS.n8990 11.666
R18535 VSS.n9061 VSS.n8987 11.666
R18536 VSS.n9069 VSS.n8991 11.666
R18537 VSS.n9077 VSS.n8986 11.666
R18538 VSS.n9085 VSS.n8992 11.666
R18539 VSS.n9093 VSS.n9015 11.666
R18540 VSS.n10179 VSS.n9217 11.666
R18541 VSS.n10257 VSS.n9211 11.666
R18542 VSS.n10247 VSS.n9208 11.666
R18543 VSS.n10188 VSS.n9212 11.666
R18544 VSS.n10191 VSS.n9207 11.666
R18545 VSS.n10195 VSS.n9213 11.666
R18546 VSS.n10199 VSS.n9206 11.666
R18547 VSS.n10261 VSS.n9214 11.666
R18548 VSS.n10205 VSS.n9210 11.666
R18549 VSS.n10089 VSS.n9307 11.666
R18550 VSS.n10167 VSS.n9301 11.666
R18551 VSS.n10157 VSS.n9298 11.666
R18552 VSS.n10098 VSS.n9302 11.666
R18553 VSS.n10101 VSS.n9297 11.666
R18554 VSS.n10105 VSS.n9303 11.666
R18555 VSS.n10109 VSS.n9296 11.666
R18556 VSS.n10171 VSS.n9304 11.666
R18557 VSS.n10115 VSS.n9300 11.666
R18558 VSS.n9999 VSS.n9397 11.666
R18559 VSS.n10077 VSS.n9391 11.666
R18560 VSS.n10067 VSS.n9388 11.666
R18561 VSS.n10008 VSS.n9392 11.666
R18562 VSS.n10011 VSS.n9387 11.666
R18563 VSS.n10015 VSS.n9393 11.666
R18564 VSS.n10019 VSS.n9386 11.666
R18565 VSS.n10081 VSS.n9394 11.666
R18566 VSS.n10025 VSS.n9390 11.666
R18567 VSS.n9909 VSS.n9487 11.666
R18568 VSS.n9987 VSS.n9481 11.666
R18569 VSS.n9977 VSS.n9478 11.666
R18570 VSS.n9918 VSS.n9482 11.666
R18571 VSS.n9921 VSS.n9477 11.666
R18572 VSS.n9925 VSS.n9483 11.666
R18573 VSS.n9929 VSS.n9476 11.666
R18574 VSS.n9991 VSS.n9484 11.666
R18575 VSS.n9935 VSS.n9480 11.666
R18576 VSS.n9819 VSS.n9577 11.666
R18577 VSS.n9897 VSS.n9571 11.666
R18578 VSS.n9887 VSS.n9568 11.666
R18579 VSS.n9828 VSS.n9572 11.666
R18580 VSS.n9831 VSS.n9567 11.666
R18581 VSS.n9835 VSS.n9573 11.666
R18582 VSS.n9839 VSS.n9566 11.666
R18583 VSS.n9901 VSS.n9574 11.666
R18584 VSS.n9845 VSS.n9570 11.666
R18585 VSS.n9729 VSS.n9667 11.666
R18586 VSS.n9807 VSS.n9661 11.666
R18587 VSS.n9797 VSS.n9658 11.666
R18588 VSS.n9738 VSS.n9662 11.666
R18589 VSS.n9741 VSS.n9657 11.666
R18590 VSS.n9745 VSS.n9663 11.666
R18591 VSS.n9749 VSS.n9656 11.666
R18592 VSS.n9811 VSS.n9664 11.666
R18593 VSS.n9755 VSS.n9660 11.666
R18594 VSS.n9183 VSS.n8934 11.666
R18595 VSS.n10366 VSS.n8936 11.666
R18596 VSS.n10360 VSS.n8941 11.666
R18597 VSS.n10354 VSS.n8947 11.666
R18598 VSS.n10348 VSS.n8953 11.666
R18599 VSS.n10342 VSS.n8958 11.666
R18600 VSS.n10336 VSS.n8965 11.666
R18601 VSS.n10330 VSS.n8971 11.666
R18602 VSS.n5669 VSS.n3581 11.666
R18603 VSS.n5781 VSS.n3583 11.666
R18604 VSS.n5775 VSS.n3588 11.666
R18605 VSS.n5769 VSS.n3594 11.666
R18606 VSS.n5763 VSS.n3600 11.666
R18607 VSS.n5757 VSS.n3606 11.666
R18608 VSS.n5751 VSS.n3611 11.666
R18609 VSS.n5745 VSS.n3618 11.666
R18610 VSS.n5739 VSS.n3624 11.666
R18611 VSS.n5791 VSS.n3523 11.666
R18612 VSS.n5903 VSS.n3525 11.666
R18613 VSS.n5897 VSS.n3530 11.666
R18614 VSS.n5891 VSS.n3536 11.666
R18615 VSS.n5885 VSS.n3542 11.666
R18616 VSS.n5879 VSS.n3548 11.666
R18617 VSS.n5873 VSS.n3553 11.666
R18618 VSS.n5867 VSS.n3560 11.666
R18619 VSS.n5861 VSS.n3566 11.666
R18620 VSS.n5913 VSS.n3465 11.666
R18621 VSS.n6025 VSS.n3467 11.666
R18622 VSS.n6019 VSS.n3472 11.666
R18623 VSS.n6013 VSS.n3478 11.666
R18624 VSS.n6007 VSS.n3484 11.666
R18625 VSS.n6001 VSS.n3490 11.666
R18626 VSS.n5995 VSS.n3495 11.666
R18627 VSS.n5989 VSS.n3502 11.666
R18628 VSS.n5983 VSS.n3508 11.666
R18629 VSS.n6035 VSS.n3407 11.666
R18630 VSS.n6147 VSS.n3409 11.666
R18631 VSS.n6141 VSS.n3414 11.666
R18632 VSS.n6135 VSS.n3420 11.666
R18633 VSS.n6129 VSS.n3426 11.666
R18634 VSS.n6123 VSS.n3432 11.666
R18635 VSS.n6117 VSS.n3437 11.666
R18636 VSS.n6111 VSS.n3444 11.666
R18637 VSS.n6105 VSS.n3450 11.666
R18638 VSS.n6157 VSS.n3349 11.666
R18639 VSS.n6269 VSS.n3351 11.666
R18640 VSS.n6263 VSS.n3356 11.666
R18641 VSS.n6257 VSS.n3362 11.666
R18642 VSS.n6251 VSS.n3368 11.666
R18643 VSS.n6245 VSS.n3374 11.666
R18644 VSS.n6239 VSS.n3379 11.666
R18645 VSS.n6233 VSS.n3386 11.666
R18646 VSS.n6227 VSS.n3392 11.666
R18647 VSS.n6279 VSS.n3291 11.666
R18648 VSS.n6391 VSS.n3293 11.666
R18649 VSS.n6385 VSS.n3298 11.666
R18650 VSS.n6379 VSS.n3304 11.666
R18651 VSS.n6373 VSS.n3310 11.666
R18652 VSS.n6367 VSS.n3316 11.666
R18653 VSS.n6361 VSS.n3321 11.666
R18654 VSS.n6355 VSS.n3328 11.666
R18655 VSS.n6349 VSS.n3334 11.666
R18656 VSS.n6401 VSS.n3233 11.666
R18657 VSS.n6513 VSS.n3235 11.666
R18658 VSS.n6507 VSS.n3240 11.666
R18659 VSS.n6501 VSS.n3246 11.666
R18660 VSS.n6495 VSS.n3252 11.666
R18661 VSS.n6489 VSS.n3258 11.666
R18662 VSS.n6483 VSS.n3263 11.666
R18663 VSS.n6477 VSS.n3270 11.666
R18664 VSS.n6471 VSS.n3276 11.666
R18665 VSS.n6535 VSS.n3149 11.666
R18666 VSS.n6600 VSS.n6599 11.666
R18667 VSS.n3177 VSS.n3144 11.666
R18668 VSS.n3185 VSS.n3146 11.666
R18669 VSS.n3193 VSS.n3143 11.666
R18670 VSS.n3201 VSS.n3147 11.666
R18671 VSS.n3209 VSS.n3142 11.666
R18672 VSS.n3217 VSS.n3148 11.666
R18673 VSS.n3225 VSS.n3157 11.666
R18674 VSS.n1177 VSS.n34 11.666
R18675 VSS.n1250 VSS.n28 11.666
R18676 VSS.n1240 VSS.n25 11.666
R18677 VSS.n1186 VSS.n29 11.666
R18678 VSS.n1189 VSS.n24 11.666
R18679 VSS.n1193 VSS.n30 11.666
R18680 VSS.n1197 VSS.n23 11.666
R18681 VSS.n1253 VSS.n31 11.666
R18682 VSS.n1203 VSS.n27 11.666
R18683 VSS.n1087 VSS.n125 11.666
R18684 VSS.n1165 VSS.n119 11.666
R18685 VSS.n1155 VSS.n116 11.666
R18686 VSS.n1096 VSS.n120 11.666
R18687 VSS.n1099 VSS.n115 11.666
R18688 VSS.n1103 VSS.n121 11.666
R18689 VSS.n1107 VSS.n114 11.666
R18690 VSS.n1169 VSS.n122 11.666
R18691 VSS.n1113 VSS.n118 11.666
R18692 VSS.n997 VSS.n215 11.666
R18693 VSS.n1075 VSS.n209 11.666
R18694 VSS.n1065 VSS.n206 11.666
R18695 VSS.n1006 VSS.n210 11.666
R18696 VSS.n1009 VSS.n205 11.666
R18697 VSS.n1013 VSS.n211 11.666
R18698 VSS.n1017 VSS.n204 11.666
R18699 VSS.n1079 VSS.n212 11.666
R18700 VSS.n1023 VSS.n208 11.666
R18701 VSS.n907 VSS.n305 11.666
R18702 VSS.n985 VSS.n299 11.666
R18703 VSS.n975 VSS.n296 11.666
R18704 VSS.n916 VSS.n300 11.666
R18705 VSS.n919 VSS.n295 11.666
R18706 VSS.n923 VSS.n301 11.666
R18707 VSS.n927 VSS.n294 11.666
R18708 VSS.n989 VSS.n302 11.666
R18709 VSS.n933 VSS.n298 11.666
R18710 VSS.n817 VSS.n395 11.666
R18711 VSS.n895 VSS.n389 11.666
R18712 VSS.n885 VSS.n386 11.666
R18713 VSS.n826 VSS.n390 11.666
R18714 VSS.n829 VSS.n385 11.666
R18715 VSS.n833 VSS.n391 11.666
R18716 VSS.n837 VSS.n384 11.666
R18717 VSS.n899 VSS.n392 11.666
R18718 VSS.n843 VSS.n388 11.666
R18719 VSS.n727 VSS.n485 11.666
R18720 VSS.n805 VSS.n479 11.666
R18721 VSS.n795 VSS.n476 11.666
R18722 VSS.n736 VSS.n480 11.666
R18723 VSS.n739 VSS.n475 11.666
R18724 VSS.n743 VSS.n481 11.666
R18725 VSS.n747 VSS.n474 11.666
R18726 VSS.n809 VSS.n482 11.666
R18727 VSS.n753 VSS.n478 11.666
R18728 VSS.n637 VSS.n575 11.666
R18729 VSS.n715 VSS.n569 11.666
R18730 VSS.n705 VSS.n566 11.666
R18731 VSS.n646 VSS.n570 11.666
R18732 VSS.n649 VSS.n565 11.666
R18733 VSS.n653 VSS.n571 11.666
R18734 VSS.n657 VSS.n564 11.666
R18735 VSS.n719 VSS.n572 11.666
R18736 VSS.n663 VSS.n568 11.666
R18737 VSS.n14729 VSS.n14728 11.636
R18738 VSS.n14730 VSS.n14729 11.636
R18739 VSS.n14730 VSS.n14358 11.636
R18740 VSS.n14736 VSS.n14358 11.636
R18741 VSS.n14737 VSS.n14736 11.636
R18742 VSS.n14738 VSS.n14737 11.636
R18743 VSS.n14738 VSS.n14354 11.636
R18744 VSS.n14744 VSS.n14354 11.636
R18745 VSS.n14745 VSS.n14744 11.636
R18746 VSS.n14746 VSS.n14745 11.636
R18747 VSS.n14746 VSS.n14350 11.636
R18748 VSS.n15997 VSS.n14015 11.636
R18749 VSS.n15991 VSS.n14015 11.636
R18750 VSS.n15991 VSS.n15990 11.636
R18751 VSS.n15990 VSS.n15989 11.636
R18752 VSS.n15989 VSS.n14019 11.636
R18753 VSS.n15983 VSS.n14019 11.636
R18754 VSS.n15983 VSS.n15982 11.636
R18755 VSS.n15982 VSS.n15981 11.636
R18756 VSS.n15981 VSS.n14023 11.636
R18757 VSS.n15975 VSS.n14023 11.636
R18758 VSS.n15975 VSS.n15974 11.636
R18759 VSS.n15951 VSS.n15950 11.636
R18760 VSS.n15951 VSS.n14035 11.636
R18761 VSS.n15957 VSS.n14035 11.636
R18762 VSS.n15958 VSS.n15957 11.636
R18763 VSS.n15959 VSS.n15958 11.636
R18764 VSS.n15959 VSS.n14031 11.636
R18765 VSS.n15965 VSS.n14031 11.636
R18766 VSS.n15966 VSS.n15965 11.636
R18767 VSS.n15967 VSS.n15966 11.636
R18768 VSS.n15967 VSS.n14027 11.636
R18769 VSS.n15973 VSS.n14027 11.636
R18770 VSS.n15923 VSS.n15922 11.636
R18771 VSS.n15924 VSS.n15923 11.636
R18772 VSS.n15924 VSS.n14050 11.636
R18773 VSS.n15930 VSS.n14050 11.636
R18774 VSS.n15931 VSS.n15930 11.636
R18775 VSS.n15932 VSS.n15931 11.636
R18776 VSS.n15932 VSS.n14046 11.636
R18777 VSS.n15939 VSS.n14046 11.636
R18778 VSS.n15940 VSS.n15939 11.636
R18779 VSS.n15941 VSS.n15940 11.636
R18780 VSS.n15941 VSS.n14039 11.636
R18781 VSS.n14191 VSS.n14190 11.636
R18782 VSS.n14190 VSS.n14189 11.636
R18783 VSS.n14189 VSS.n14161 11.636
R18784 VSS.n14183 VSS.n14161 11.636
R18785 VSS.n14183 VSS.n14182 11.636
R18786 VSS.n14182 VSS.n14181 11.636
R18787 VSS.n14181 VSS.n14165 11.636
R18788 VSS.n14175 VSS.n14165 11.636
R18789 VSS.n14175 VSS.n14174 11.636
R18790 VSS.n14174 VSS.n14173 11.636
R18791 VSS.n14173 VSS.n14169 11.636
R18792 VSS.n15393 VSS.n14204 11.636
R18793 VSS.n15394 VSS.n15393 11.636
R18794 VSS.n15395 VSS.n15394 11.636
R18795 VSS.n15395 VSS.n14200 11.636
R18796 VSS.n15401 VSS.n14200 11.636
R18797 VSS.n15402 VSS.n15401 11.636
R18798 VSS.n15403 VSS.n15402 11.636
R18799 VSS.n15403 VSS.n14196 11.636
R18800 VSS.n15409 VSS.n14196 11.636
R18801 VSS.n15410 VSS.n15409 11.636
R18802 VSS.n15411 VSS.n15410 11.636
R18803 VSS.n15360 VSS.n14219 11.636
R18804 VSS.n15366 VSS.n14219 11.636
R18805 VSS.n15367 VSS.n15366 11.636
R18806 VSS.n15368 VSS.n15367 11.636
R18807 VSS.n15368 VSS.n14215 11.636
R18808 VSS.n15374 VSS.n14215 11.636
R18809 VSS.n15375 VSS.n15374 11.636
R18810 VSS.n15377 VSS.n15375 11.636
R18811 VSS.n15377 VSS.n15376 11.636
R18812 VSS.n15376 VSS.n14211 11.636
R18813 VSS.n15384 VSS.n14211 11.636
R18814 VSS.n14831 VSS.n14321 11.636
R18815 VSS.n14831 VSS.n14830 11.636
R18816 VSS.n14830 VSS.n14829 11.636
R18817 VSS.n14829 VSS.n14803 11.636
R18818 VSS.n14823 VSS.n14803 11.636
R18819 VSS.n14823 VSS.n14822 11.636
R18820 VSS.n14822 VSS.n14821 11.636
R18821 VSS.n14821 VSS.n14808 11.636
R18822 VSS.n14815 VSS.n14808 11.636
R18823 VSS.n14815 VSS.n14814 11.636
R18824 VSS.n14814 VSS.n14223 11.636
R18825 VSS.n14781 VSS.n14780 11.636
R18826 VSS.n14781 VSS.n14331 11.636
R18827 VSS.n14787 VSS.n14331 11.636
R18828 VSS.n14788 VSS.n14787 11.636
R18829 VSS.n14789 VSS.n14788 11.636
R18830 VSS.n14789 VSS.n14327 11.636
R18831 VSS.n14795 VSS.n14327 11.636
R18832 VSS.n14796 VSS.n14795 11.636
R18833 VSS.n14797 VSS.n14796 11.636
R18834 VSS.n14797 VSS.n14322 11.636
R18835 VSS.n14838 VSS.n14322 11.636
R18836 VSS.n14753 VSS.n14752 11.636
R18837 VSS.n14754 VSS.n14753 11.636
R18838 VSS.n14754 VSS.n14346 11.636
R18839 VSS.n14760 VSS.n14346 11.636
R18840 VSS.n14761 VSS.n14760 11.636
R18841 VSS.n14762 VSS.n14761 11.636
R18842 VSS.n14762 VSS.n14342 11.636
R18843 VSS.n14769 VSS.n14342 11.636
R18844 VSS.n14770 VSS.n14769 11.636
R18845 VSS.n14771 VSS.n14770 11.636
R18846 VSS.n14771 VSS.n14335 11.636
R18847 VSS.n12789 VSS.n12724 11.636
R18848 VSS.n12729 VSS.n12724 11.636
R18849 VSS.n12782 VSS.n12729 11.636
R18850 VSS.n12782 VSS.n12781 11.636
R18851 VSS.n12781 VSS.n12780 11.636
R18852 VSS.n12780 VSS.n12730 11.636
R18853 VSS.n12774 VSS.n12730 11.636
R18854 VSS.n12774 VSS.n12773 11.636
R18855 VSS.n12773 VSS.n12772 11.636
R18856 VSS.n12772 VSS.n12734 11.636
R18857 VSS.n12766 VSS.n12734 11.636
R18858 VSS.n12212 VSS.n12064 11.636
R18859 VSS.n12206 VSS.n12064 11.636
R18860 VSS.n12206 VSS.n12205 11.636
R18861 VSS.n12205 VSS.n12204 11.636
R18862 VSS.n12204 VSS.n12068 11.636
R18863 VSS.n12198 VSS.n12068 11.636
R18864 VSS.n12198 VSS.n12197 11.636
R18865 VSS.n12197 VSS.n12196 11.636
R18866 VSS.n12196 VSS.n12072 11.636
R18867 VSS.n12190 VSS.n12072 11.636
R18868 VSS.n12190 VSS.n12189 11.636
R18869 VSS.n12166 VSS.n12165 11.636
R18870 VSS.n12166 VSS.n12084 11.636
R18871 VSS.n12172 VSS.n12084 11.636
R18872 VSS.n12173 VSS.n12172 11.636
R18873 VSS.n12174 VSS.n12173 11.636
R18874 VSS.n12174 VSS.n12080 11.636
R18875 VSS.n12180 VSS.n12080 11.636
R18876 VSS.n12181 VSS.n12180 11.636
R18877 VSS.n12182 VSS.n12181 11.636
R18878 VSS.n12182 VSS.n12076 11.636
R18879 VSS.n12188 VSS.n12076 11.636
R18880 VSS.n12138 VSS.n11528 11.636
R18881 VSS.n12139 VSS.n12138 11.636
R18882 VSS.n12139 VSS.n12132 11.636
R18883 VSS.n12145 VSS.n12132 11.636
R18884 VSS.n12146 VSS.n12145 11.636
R18885 VSS.n12147 VSS.n12146 11.636
R18886 VSS.n12147 VSS.n12128 11.636
R18887 VSS.n12154 VSS.n12128 11.636
R18888 VSS.n12155 VSS.n12154 11.636
R18889 VSS.n12156 VSS.n12155 11.636
R18890 VSS.n12156 VSS.n12088 11.636
R18891 VSS.n12458 VSS.n11515 11.636
R18892 VSS.n11519 VSS.n11515 11.636
R18893 VSS.n12451 VSS.n11519 11.636
R18894 VSS.n12451 VSS.n12450 11.636
R18895 VSS.n12450 VSS.n12449 11.636
R18896 VSS.n12449 VSS.n11520 11.636
R18897 VSS.n12443 VSS.n11520 11.636
R18898 VSS.n12443 VSS.n12442 11.636
R18899 VSS.n12442 VSS.n12441 11.636
R18900 VSS.n12441 VSS.n11524 11.636
R18901 VSS.n12435 VSS.n11524 11.636
R18902 VSS.n12485 VSS.n12484 11.636
R18903 VSS.n12484 VSS.n12483 11.636
R18904 VSS.n12483 VSS.n11500 11.636
R18905 VSS.n12477 VSS.n11500 11.636
R18906 VSS.n12477 VSS.n12476 11.636
R18907 VSS.n12476 VSS.n12475 11.636
R18908 VSS.n12475 VSS.n11504 11.636
R18909 VSS.n12469 VSS.n11504 11.636
R18910 VSS.n12469 VSS.n12468 11.636
R18911 VSS.n12468 VSS.n12467 11.636
R18912 VSS.n12467 VSS.n11508 11.636
R18913 VSS.n13349 VSS.n12498 11.636
R18914 VSS.n13350 VSS.n13349 11.636
R18915 VSS.n13351 VSS.n13350 11.636
R18916 VSS.n13351 VSS.n12494 11.636
R18917 VSS.n13357 VSS.n12494 11.636
R18918 VSS.n13358 VSS.n13357 11.636
R18919 VSS.n13359 VSS.n13358 11.636
R18920 VSS.n13359 VSS.n12490 11.636
R18921 VSS.n13365 VSS.n12490 11.636
R18922 VSS.n13366 VSS.n13365 11.636
R18923 VSS.n13367 VSS.n13366 11.636
R18924 VSS.n12626 VSS.n12625 11.636
R18925 VSS.n12625 VSS.n12624 11.636
R18926 VSS.n12624 VSS.n12601 11.636
R18927 VSS.n12618 VSS.n12601 11.636
R18928 VSS.n12618 VSS.n12617 11.636
R18929 VSS.n12617 VSS.n12616 11.636
R18930 VSS.n12616 VSS.n12605 11.636
R18931 VSS.n12610 VSS.n12605 11.636
R18932 VSS.n12610 VSS.n12609 11.636
R18933 VSS.n12609 VSS.n12504 11.636
R18934 VSS.n13342 VSS.n12504 11.636
R18935 VSS.n13100 VSS.n12639 11.636
R18936 VSS.n13101 VSS.n13100 11.636
R18937 VSS.n13102 VSS.n13101 11.636
R18938 VSS.n13102 VSS.n12635 11.636
R18939 VSS.n13108 VSS.n12635 11.636
R18940 VSS.n13109 VSS.n13108 11.636
R18941 VSS.n13110 VSS.n13109 11.636
R18942 VSS.n13110 VSS.n12631 11.636
R18943 VSS.n13116 VSS.n12631 11.636
R18944 VSS.n13117 VSS.n13116 11.636
R18945 VSS.n13118 VSS.n13117 11.636
R18946 VSS.n12765 VSS.n12764 11.636
R18947 VSS.n12764 VSS.n12738 11.636
R18948 VSS.n12758 VSS.n12738 11.636
R18949 VSS.n12758 VSS.n12757 11.636
R18950 VSS.n12757 VSS.n12756 11.636
R18951 VSS.n12756 VSS.n12742 11.636
R18952 VSS.n12750 VSS.n12742 11.636
R18953 VSS.n12750 VSS.n12749 11.636
R18954 VSS.n12749 VSS.n12748 11.636
R18955 VSS.n12748 VSS.n12645 11.636
R18956 VSS.n13093 VSS.n12645 11.636
R18957 VSS.n7843 VSS.n7842 11.636
R18958 VSS.n7843 VSS.n7667 11.636
R18959 VSS.n7849 VSS.n7667 11.636
R18960 VSS.n7850 VSS.n7849 11.636
R18961 VSS.n7851 VSS.n7850 11.636
R18962 VSS.n7851 VSS.n7663 11.636
R18963 VSS.n7857 VSS.n7663 11.636
R18964 VSS.n7858 VSS.n7857 11.636
R18965 VSS.n7859 VSS.n7858 11.636
R18966 VSS.n7859 VSS.n7659 11.636
R18967 VSS.n7865 VSS.n7659 11.636
R18968 VSS.n7180 VSS.n7179 11.636
R18969 VSS.n7180 VSS.n7001 11.636
R18970 VSS.n7186 VSS.n7001 11.636
R18971 VSS.n7187 VSS.n7186 11.636
R18972 VSS.n7188 VSS.n7187 11.636
R18973 VSS.n7188 VSS.n6997 11.636
R18974 VSS.n7194 VSS.n6997 11.636
R18975 VSS.n7195 VSS.n7194 11.636
R18976 VSS.n7196 VSS.n7195 11.636
R18977 VSS.n7196 VSS.n6993 11.636
R18978 VSS.n7202 VSS.n6993 11.636
R18979 VSS.n7226 VSS.n6981 11.636
R18980 VSS.n7220 VSS.n6981 11.636
R18981 VSS.n7220 VSS.n7219 11.636
R18982 VSS.n7219 VSS.n7218 11.636
R18983 VSS.n7218 VSS.n6985 11.636
R18984 VSS.n7212 VSS.n6985 11.636
R18985 VSS.n7212 VSS.n7211 11.636
R18986 VSS.n7211 VSS.n7210 11.636
R18987 VSS.n7210 VSS.n6989 11.636
R18988 VSS.n7204 VSS.n6989 11.636
R18989 VSS.n7204 VSS.n7203 11.636
R18990 VSS.n8805 VSS.n8804 11.636
R18991 VSS.n8805 VSS.n7235 11.636
R18992 VSS.n8811 VSS.n7235 11.636
R18993 VSS.n8812 VSS.n8811 11.636
R18994 VSS.n8813 VSS.n8812 11.636
R18995 VSS.n8813 VSS.n7231 11.636
R18996 VSS.n8819 VSS.n7231 11.636
R18997 VSS.n8820 VSS.n8819 11.636
R18998 VSS.n8821 VSS.n8820 11.636
R18999 VSS.n8821 VSS.n7227 11.636
R19000 VSS.n8827 VSS.n7227 11.636
R19001 VSS.n7366 VSS.n7337 11.636
R19002 VSS.n7360 VSS.n7337 11.636
R19003 VSS.n7360 VSS.n7359 11.636
R19004 VSS.n7359 VSS.n7358 11.636
R19005 VSS.n7358 VSS.n7341 11.636
R19006 VSS.n7352 VSS.n7341 11.636
R19007 VSS.n7352 VSS.n7351 11.636
R19008 VSS.n7351 VSS.n7350 11.636
R19009 VSS.n7350 VSS.n7345 11.636
R19010 VSS.n7345 VSS.n7240 11.636
R19011 VSS.n8802 VSS.n7240 11.636
R19012 VSS.n8583 VSS.n8582 11.636
R19013 VSS.n8583 VSS.n7375 11.636
R19014 VSS.n8589 VSS.n7375 11.636
R19015 VSS.n8590 VSS.n8589 11.636
R19016 VSS.n8591 VSS.n8590 11.636
R19017 VSS.n8591 VSS.n7371 11.636
R19018 VSS.n8597 VSS.n7371 11.636
R19019 VSS.n8598 VSS.n8597 11.636
R19020 VSS.n8599 VSS.n8598 11.636
R19021 VSS.n8599 VSS.n7367 11.636
R19022 VSS.n8605 VSS.n7367 11.636
R19023 VSS.n7506 VSS.n7477 11.636
R19024 VSS.n7500 VSS.n7477 11.636
R19025 VSS.n7500 VSS.n7499 11.636
R19026 VSS.n7499 VSS.n7498 11.636
R19027 VSS.n7498 VSS.n7481 11.636
R19028 VSS.n7492 VSS.n7481 11.636
R19029 VSS.n7492 VSS.n7491 11.636
R19030 VSS.n7491 VSS.n7490 11.636
R19031 VSS.n7490 VSS.n7485 11.636
R19032 VSS.n7485 VSS.n7380 11.636
R19033 VSS.n8580 VSS.n7380 11.636
R19034 VSS.n8225 VSS.n8224 11.636
R19035 VSS.n8225 VSS.n7515 11.636
R19036 VSS.n8231 VSS.n7515 11.636
R19037 VSS.n8232 VSS.n8231 11.636
R19038 VSS.n8233 VSS.n8232 11.636
R19039 VSS.n8233 VSS.n7511 11.636
R19040 VSS.n8239 VSS.n7511 11.636
R19041 VSS.n8240 VSS.n8239 11.636
R19042 VSS.n8241 VSS.n8240 11.636
R19043 VSS.n8241 VSS.n7507 11.636
R19044 VSS.n8247 VSS.n7507 11.636
R19045 VSS.n7646 VSS.n7617 11.636
R19046 VSS.n7640 VSS.n7617 11.636
R19047 VSS.n7640 VSS.n7639 11.636
R19048 VSS.n7639 VSS.n7638 11.636
R19049 VSS.n7638 VSS.n7621 11.636
R19050 VSS.n7632 VSS.n7621 11.636
R19051 VSS.n7632 VSS.n7631 11.636
R19052 VSS.n7631 VSS.n7630 11.636
R19053 VSS.n7630 VSS.n7625 11.636
R19054 VSS.n7625 VSS.n7520 11.636
R19055 VSS.n8222 VSS.n7520 11.636
R19056 VSS.n7867 VSS.n7866 11.636
R19057 VSS.n7867 VSS.n7655 11.636
R19058 VSS.n7873 VSS.n7655 11.636
R19059 VSS.n7874 VSS.n7873 11.636
R19060 VSS.n7875 VSS.n7874 11.636
R19061 VSS.n7875 VSS.n7651 11.636
R19062 VSS.n7881 VSS.n7651 11.636
R19063 VSS.n7882 VSS.n7881 11.636
R19064 VSS.n7883 VSS.n7882 11.636
R19065 VSS.n7883 VSS.n7647 11.636
R19066 VSS.n7889 VSS.n7647 11.636
R19067 VSS.n6832 VSS.n6831 11.636
R19068 VSS.n6833 VSS.n6832 11.636
R19069 VSS.n6833 VSS.n6752 11.636
R19070 VSS.n6839 VSS.n6752 11.636
R19071 VSS.n6840 VSS.n6839 11.636
R19072 VSS.n6841 VSS.n6840 11.636
R19073 VSS.n6841 VSS.n6748 11.636
R19074 VSS.n6847 VSS.n6748 11.636
R19075 VSS.n6848 VSS.n6847 11.636
R19076 VSS.n6849 VSS.n6848 11.636
R19077 VSS.n6849 VSS.n6744 11.636
R19078 VSS.n6825 VSS.n6824 11.636
R19079 VSS.n6824 VSS.n6823 11.636
R19080 VSS.n6823 VSS.n6761 11.636
R19081 VSS.n6817 VSS.n6816 11.636
R19082 VSS.n6816 VSS.n6815 11.636
R19083 VSS.n6809 VSS.n6768 11.636
R19084 VSS.n6809 VSS.n6808 11.636
R19085 VSS.n6808 VSS.n6807 11.636
R19086 VSS.n6807 VSS.n6769 11.636
R19087 VSS.n6800 VSS.n6799 11.636
R19088 VSS.n6799 VSS.n6773 11.636
R19089 VSS.n6793 VSS.n6773 11.636
R19090 VSS.n6793 VSS.n6792 11.636
R19091 VSS.n6792 VSS.n6791 11.636
R19092 VSS.n6791 VSS.n6777 11.636
R19093 VSS.n6785 VSS.n6777 11.636
R19094 VSS.n6785 VSS.n6784 11.636
R19095 VSS.n6784 VSS.n6783 11.636
R19096 VSS.n6783 VSS.n6730 11.636
R19097 VSS.n6879 VSS.n6730 11.636
R19098 VSS.n6856 VSS.n6855 11.636
R19099 VSS.n6857 VSS.n6856 11.636
R19100 VSS.n6857 VSS.n6740 11.636
R19101 VSS.n6863 VSS.n6740 11.636
R19102 VSS.n6864 VSS.n6863 11.636
R19103 VSS.n6865 VSS.n6864 11.636
R19104 VSS.n6865 VSS.n6736 11.636
R19105 VSS.n6871 VSS.n6736 11.636
R19106 VSS.n6872 VSS.n6871 11.636
R19107 VSS.n6873 VSS.n6872 11.636
R19108 VSS.n6873 VSS.n6729 11.636
R19109 VSS.n4242 VSS.n4177 11.636
R19110 VSS.n4182 VSS.n4177 11.636
R19111 VSS.n4235 VSS.n4182 11.636
R19112 VSS.n4235 VSS.n4234 11.636
R19113 VSS.n4234 VSS.n4233 11.636
R19114 VSS.n4233 VSS.n4183 11.636
R19115 VSS.n4227 VSS.n4183 11.636
R19116 VSS.n4227 VSS.n4226 11.636
R19117 VSS.n4226 VSS.n4225 11.636
R19118 VSS.n4225 VSS.n4187 11.636
R19119 VSS.n4219 VSS.n4187 11.636
R19120 VSS.n5655 VSS.n5654 11.636
R19121 VSS.n5654 VSS.n5653 11.636
R19122 VSS.n5653 VSS.n3649 11.636
R19123 VSS.n5647 VSS.n3649 11.636
R19124 VSS.n5647 VSS.n5646 11.636
R19125 VSS.n5646 VSS.n5645 11.636
R19126 VSS.n5645 VSS.n3653 11.636
R19127 VSS.n5639 VSS.n3653 11.636
R19128 VSS.n5639 VSS.n5638 11.636
R19129 VSS.n5638 VSS.n5637 11.636
R19130 VSS.n5637 VSS.n3657 11.636
R19131 VSS.n5613 VSS.n3669 11.636
R19132 VSS.n5614 VSS.n5613 11.636
R19133 VSS.n5615 VSS.n5614 11.636
R19134 VSS.n5615 VSS.n3665 11.636
R19135 VSS.n5621 VSS.n3665 11.636
R19136 VSS.n5622 VSS.n5621 11.636
R19137 VSS.n5623 VSS.n5622 11.636
R19138 VSS.n5623 VSS.n3661 11.636
R19139 VSS.n5629 VSS.n3661 11.636
R19140 VSS.n5630 VSS.n5629 11.636
R19141 VSS.n5631 VSS.n5630 11.636
R19142 VSS.n3797 VSS.n3796 11.636
R19143 VSS.n3796 VSS.n3795 11.636
R19144 VSS.n3795 VSS.n3772 11.636
R19145 VSS.n3789 VSS.n3772 11.636
R19146 VSS.n3789 VSS.n3788 11.636
R19147 VSS.n3788 VSS.n3787 11.636
R19148 VSS.n3787 VSS.n3776 11.636
R19149 VSS.n3781 VSS.n3776 11.636
R19150 VSS.n3781 VSS.n3780 11.636
R19151 VSS.n3780 VSS.n3675 11.636
R19152 VSS.n5606 VSS.n3675 11.636
R19153 VSS.n5267 VSS.n3810 11.636
R19154 VSS.n5268 VSS.n5267 11.636
R19155 VSS.n5269 VSS.n5268 11.636
R19156 VSS.n5269 VSS.n3806 11.636
R19157 VSS.n5275 VSS.n3806 11.636
R19158 VSS.n5276 VSS.n5275 11.636
R19159 VSS.n5277 VSS.n5276 11.636
R19160 VSS.n5277 VSS.n3802 11.636
R19161 VSS.n5283 VSS.n3802 11.636
R19162 VSS.n5284 VSS.n5283 11.636
R19163 VSS.n5285 VSS.n5284 11.636
R19164 VSS.n3938 VSS.n3937 11.636
R19165 VSS.n3937 VSS.n3936 11.636
R19166 VSS.n3936 VSS.n3913 11.636
R19167 VSS.n3930 VSS.n3913 11.636
R19168 VSS.n3930 VSS.n3929 11.636
R19169 VSS.n3929 VSS.n3928 11.636
R19170 VSS.n3928 VSS.n3917 11.636
R19171 VSS.n3922 VSS.n3917 11.636
R19172 VSS.n3922 VSS.n3921 11.636
R19173 VSS.n3921 VSS.n3816 11.636
R19174 VSS.n5260 VSS.n3816 11.636
R19175 VSS.n4910 VSS.n3951 11.636
R19176 VSS.n4911 VSS.n4910 11.636
R19177 VSS.n4912 VSS.n4911 11.636
R19178 VSS.n4912 VSS.n3947 11.636
R19179 VSS.n4918 VSS.n3947 11.636
R19180 VSS.n4919 VSS.n4918 11.636
R19181 VSS.n4920 VSS.n4919 11.636
R19182 VSS.n4920 VSS.n3943 11.636
R19183 VSS.n4926 VSS.n3943 11.636
R19184 VSS.n4927 VSS.n4926 11.636
R19185 VSS.n4928 VSS.n4927 11.636
R19186 VSS.n4079 VSS.n4078 11.636
R19187 VSS.n4078 VSS.n4077 11.636
R19188 VSS.n4077 VSS.n4054 11.636
R19189 VSS.n4071 VSS.n4054 11.636
R19190 VSS.n4071 VSS.n4070 11.636
R19191 VSS.n4070 VSS.n4069 11.636
R19192 VSS.n4069 VSS.n4058 11.636
R19193 VSS.n4063 VSS.n4058 11.636
R19194 VSS.n4063 VSS.n4062 11.636
R19195 VSS.n4062 VSS.n3957 11.636
R19196 VSS.n4903 VSS.n3957 11.636
R19197 VSS.n4553 VSS.n4092 11.636
R19198 VSS.n4554 VSS.n4553 11.636
R19199 VSS.n4555 VSS.n4554 11.636
R19200 VSS.n4555 VSS.n4088 11.636
R19201 VSS.n4561 VSS.n4088 11.636
R19202 VSS.n4562 VSS.n4561 11.636
R19203 VSS.n4563 VSS.n4562 11.636
R19204 VSS.n4563 VSS.n4084 11.636
R19205 VSS.n4569 VSS.n4084 11.636
R19206 VSS.n4570 VSS.n4569 11.636
R19207 VSS.n4571 VSS.n4570 11.636
R19208 VSS.n4218 VSS.n4217 11.636
R19209 VSS.n4217 VSS.n4191 11.636
R19210 VSS.n4211 VSS.n4191 11.636
R19211 VSS.n4211 VSS.n4210 11.636
R19212 VSS.n4210 VSS.n4209 11.636
R19213 VSS.n4209 VSS.n4195 11.636
R19214 VSS.n4203 VSS.n4195 11.636
R19215 VSS.n4203 VSS.n4202 11.636
R19216 VSS.n4202 VSS.n4201 11.636
R19217 VSS.n4201 VSS.n4098 11.636
R19218 VSS.n4546 VSS.n4098 11.636
R19219 VSS.n1970 VSS.n1969 11.636
R19220 VSS.n1971 VSS.n1970 11.636
R19221 VSS.n1971 VSS.n1599 11.636
R19222 VSS.n1977 VSS.n1599 11.636
R19223 VSS.n1978 VSS.n1977 11.636
R19224 VSS.n1979 VSS.n1978 11.636
R19225 VSS.n1979 VSS.n1595 11.636
R19226 VSS.n1985 VSS.n1595 11.636
R19227 VSS.n1986 VSS.n1985 11.636
R19228 VSS.n1987 VSS.n1986 11.636
R19229 VSS.n1987 VSS.n1591 11.636
R19230 VSS.n2997 VSS.n2996 11.636
R19231 VSS.n2998 VSS.n2997 11.636
R19232 VSS.n2998 VSS.n1291 11.636
R19233 VSS.n3004 VSS.n1291 11.636
R19234 VSS.n3005 VSS.n3004 11.636
R19235 VSS.n3006 VSS.n3005 11.636
R19236 VSS.n3006 VSS.n1287 11.636
R19237 VSS.n3012 VSS.n1287 11.636
R19238 VSS.n3013 VSS.n3012 11.636
R19239 VSS.n3014 VSS.n3013 11.636
R19240 VSS.n3014 VSS.n1283 11.636
R19241 VSS.n3038 VSS.n1268 11.636
R19242 VSS.n3038 VSS.n3037 11.636
R19243 VSS.n3037 VSS.n3036 11.636
R19244 VSS.n3036 VSS.n1275 11.636
R19245 VSS.n3030 VSS.n1275 11.636
R19246 VSS.n3030 VSS.n3029 11.636
R19247 VSS.n3029 VSS.n3028 11.636
R19248 VSS.n3028 VSS.n1279 11.636
R19249 VSS.n3022 VSS.n1279 11.636
R19250 VSS.n3022 VSS.n3021 11.636
R19251 VSS.n3021 VSS.n3020 11.636
R19252 VSS.n1432 VSS.n1431 11.636
R19253 VSS.n1431 VSS.n1430 11.636
R19254 VSS.n1430 VSS.n1402 11.636
R19255 VSS.n1424 VSS.n1402 11.636
R19256 VSS.n1424 VSS.n1423 11.636
R19257 VSS.n1423 VSS.n1422 11.636
R19258 VSS.n1422 VSS.n1406 11.636
R19259 VSS.n1416 VSS.n1406 11.636
R19260 VSS.n1416 VSS.n1415 11.636
R19261 VSS.n1415 VSS.n1414 11.636
R19262 VSS.n1414 VSS.n1410 11.636
R19263 VSS.n2634 VSS.n1445 11.636
R19264 VSS.n2635 VSS.n2634 11.636
R19265 VSS.n2636 VSS.n2635 11.636
R19266 VSS.n2636 VSS.n1441 11.636
R19267 VSS.n2642 VSS.n1441 11.636
R19268 VSS.n2643 VSS.n2642 11.636
R19269 VSS.n2644 VSS.n2643 11.636
R19270 VSS.n2644 VSS.n1437 11.636
R19271 VSS.n2650 VSS.n1437 11.636
R19272 VSS.n2651 VSS.n2650 11.636
R19273 VSS.n2652 VSS.n2651 11.636
R19274 VSS.n2601 VSS.n1460 11.636
R19275 VSS.n2607 VSS.n1460 11.636
R19276 VSS.n2608 VSS.n2607 11.636
R19277 VSS.n2609 VSS.n2608 11.636
R19278 VSS.n2609 VSS.n1456 11.636
R19279 VSS.n2615 VSS.n1456 11.636
R19280 VSS.n2616 VSS.n2615 11.636
R19281 VSS.n2618 VSS.n2616 11.636
R19282 VSS.n2618 VSS.n2617 11.636
R19283 VSS.n2617 VSS.n1452 11.636
R19284 VSS.n2625 VSS.n1452 11.636
R19285 VSS.n2072 VSS.n1562 11.636
R19286 VSS.n2072 VSS.n2071 11.636
R19287 VSS.n2071 VSS.n2070 11.636
R19288 VSS.n2070 VSS.n2044 11.636
R19289 VSS.n2064 VSS.n2044 11.636
R19290 VSS.n2064 VSS.n2063 11.636
R19291 VSS.n2063 VSS.n2062 11.636
R19292 VSS.n2062 VSS.n2049 11.636
R19293 VSS.n2056 VSS.n2049 11.636
R19294 VSS.n2056 VSS.n2055 11.636
R19295 VSS.n2055 VSS.n1464 11.636
R19296 VSS.n2022 VSS.n2021 11.636
R19297 VSS.n2022 VSS.n1572 11.636
R19298 VSS.n2028 VSS.n1572 11.636
R19299 VSS.n2029 VSS.n2028 11.636
R19300 VSS.n2030 VSS.n2029 11.636
R19301 VSS.n2030 VSS.n1568 11.636
R19302 VSS.n2036 VSS.n1568 11.636
R19303 VSS.n2037 VSS.n2036 11.636
R19304 VSS.n2038 VSS.n2037 11.636
R19305 VSS.n2038 VSS.n1563 11.636
R19306 VSS.n2079 VSS.n1563 11.636
R19307 VSS.n1994 VSS.n1993 11.636
R19308 VSS.n1995 VSS.n1994 11.636
R19309 VSS.n1995 VSS.n1587 11.636
R19310 VSS.n2001 VSS.n1587 11.636
R19311 VSS.n2002 VSS.n2001 11.636
R19312 VSS.n2003 VSS.n2002 11.636
R19313 VSS.n2003 VSS.n1583 11.636
R19314 VSS.n2010 VSS.n1583 11.636
R19315 VSS.n2011 VSS.n2010 11.636
R19316 VSS.n2012 VSS.n2011 11.636
R19317 VSS.n2012 VSS.n1576 11.636
R19318 sky130_asc_res_xhigh_po_2p85_1_16/VGND VSS.n17485 10.79
R19319 sky130_asc_res_xhigh_po_2p85_1_17/VGND VSS.n13965 10.79
R19320 sky130_asc_pnp_05v5_W3p40L3p40_1_0/Collector VSS.n6761 10.731
R19321 VSS.n10372 VSS.n10371 10.438
R19322 VSS.n6768 sky130_asc_pnp_05v5_W3p40L3p40_1_0/xm1/Collector 10.343
R19323 VSS.n6881 VSS.n6728 10.299
R19324 VSS.n17393 VSS.n17391 9.955
R19325 VSS.n17457 VSS.n16048 9.955
R19326 VSS.n17450 VSS.n17449 9.955
R19327 VSS.n17403 VSS.n17400 9.955
R19328 VSS.n17437 VSS.n17406 9.955
R19329 VSS.n17431 VSS.n17410 9.955
R19330 VSS.n17425 VSS.n17414 9.955
R19331 VSS.n17419 VSS.n17417 9.955
R19332 VSS.n17301 VSS.n16091 9.955
R19333 VSS.n17294 VSS.n17293 9.955
R19334 VSS.n17234 VSS.n17231 9.955
R19335 VSS.n17281 VSS.n17237 9.955
R19336 VSS.n17275 VSS.n17241 9.955
R19337 VSS.n17269 VSS.n17245 9.955
R19338 VSS.n17263 VSS.n17248 9.955
R19339 VSS.n17258 VSS.n17251 9.955
R19340 VSS.n17211 VSS.n16181 9.955
R19341 VSS.n17204 VSS.n17203 9.955
R19342 VSS.n17144 VSS.n17141 9.955
R19343 VSS.n17191 VSS.n17147 9.955
R19344 VSS.n17185 VSS.n17151 9.955
R19345 VSS.n17179 VSS.n17155 9.955
R19346 VSS.n17173 VSS.n17158 9.955
R19347 VSS.n17168 VSS.n17161 9.955
R19348 VSS.n17121 VSS.n16271 9.955
R19349 VSS.n17114 VSS.n17113 9.955
R19350 VSS.n17054 VSS.n17051 9.955
R19351 VSS.n17101 VSS.n17057 9.955
R19352 VSS.n17095 VSS.n17061 9.955
R19353 VSS.n17089 VSS.n17065 9.955
R19354 VSS.n17083 VSS.n17068 9.955
R19355 VSS.n17078 VSS.n17071 9.955
R19356 VSS.n17031 VSS.n16361 9.955
R19357 VSS.n17024 VSS.n17023 9.955
R19358 VSS.n16964 VSS.n16961 9.955
R19359 VSS.n17011 VSS.n16967 9.955
R19360 VSS.n17005 VSS.n16971 9.955
R19361 VSS.n16999 VSS.n16975 9.955
R19362 VSS.n16993 VSS.n16978 9.955
R19363 VSS.n16988 VSS.n16981 9.955
R19364 VSS.n16941 VSS.n16451 9.955
R19365 VSS.n16934 VSS.n16933 9.955
R19366 VSS.n16874 VSS.n16871 9.955
R19367 VSS.n16921 VSS.n16877 9.955
R19368 VSS.n16915 VSS.n16881 9.955
R19369 VSS.n16909 VSS.n16885 9.955
R19370 VSS.n16903 VSS.n16888 9.955
R19371 VSS.n16898 VSS.n16891 9.955
R19372 VSS.n16851 VSS.n16541 9.955
R19373 VSS.n16844 VSS.n16843 9.955
R19374 VSS.n16784 VSS.n16781 9.955
R19375 VSS.n16831 VSS.n16787 9.955
R19376 VSS.n16825 VSS.n16791 9.955
R19377 VSS.n16819 VSS.n16795 9.955
R19378 VSS.n16813 VSS.n16798 9.955
R19379 VSS.n16808 VSS.n16801 9.955
R19380 VSS.n16761 VSS.n16631 9.955
R19381 VSS.n16754 VSS.n16753 9.955
R19382 VSS.n16694 VSS.n16691 9.955
R19383 VSS.n16741 VSS.n16697 9.955
R19384 VSS.n16735 VSS.n16701 9.955
R19385 VSS.n16729 VSS.n16705 9.955
R19386 VSS.n16723 VSS.n16708 9.955
R19387 VSS.n16718 VSS.n16711 9.955
R19388 VSS.n11229 VSS.n11098 9.955
R19389 VSS.n11222 VSS.n11221 9.955
R19390 VSS.n11161 VSS.n11158 9.955
R19391 VSS.n11209 VSS.n11164 9.955
R19392 VSS.n11203 VSS.n11168 9.955
R19393 VSS.n11197 VSS.n11171 9.955
R19394 VSS.n11192 VSS.n11174 9.955
R19395 VSS.n11186 VSS.n11177 9.955
R19396 VSS.n11319 VSS.n11008 9.955
R19397 VSS.n11312 VSS.n11311 9.955
R19398 VSS.n11251 VSS.n11248 9.955
R19399 VSS.n11299 VSS.n11254 9.955
R19400 VSS.n11293 VSS.n11258 9.955
R19401 VSS.n11287 VSS.n11261 9.955
R19402 VSS.n11282 VSS.n11264 9.955
R19403 VSS.n11276 VSS.n11267 9.955
R19404 VSS.n11409 VSS.n10918 9.955
R19405 VSS.n11402 VSS.n11401 9.955
R19406 VSS.n11341 VSS.n11338 9.955
R19407 VSS.n11389 VSS.n11344 9.955
R19408 VSS.n11383 VSS.n11348 9.955
R19409 VSS.n11377 VSS.n11351 9.955
R19410 VSS.n11372 VSS.n11354 9.955
R19411 VSS.n11366 VSS.n11357 9.955
R19412 VSS.n13529 VSS.n10828 9.955
R19413 VSS.n13522 VSS.n13521 9.955
R19414 VSS.n13460 VSS.n11428 9.955
R19415 VSS.n13508 VSS.n13463 9.955
R19416 VSS.n13502 VSS.n13467 9.955
R19417 VSS.n13496 VSS.n13470 9.955
R19418 VSS.n13491 VSS.n13473 9.955
R19419 VSS.n13485 VSS.n13476 9.955
R19420 VSS.n13619 VSS.n10738 9.955
R19421 VSS.n13612 VSS.n13611 9.955
R19422 VSS.n13551 VSS.n13548 9.955
R19423 VSS.n13599 VSS.n13554 9.955
R19424 VSS.n13593 VSS.n13558 9.955
R19425 VSS.n13587 VSS.n13561 9.955
R19426 VSS.n13582 VSS.n13564 9.955
R19427 VSS.n13576 VSS.n13567 9.955
R19428 VSS.n13709 VSS.n10648 9.955
R19429 VSS.n13702 VSS.n13701 9.955
R19430 VSS.n13641 VSS.n13638 9.955
R19431 VSS.n13689 VSS.n13644 9.955
R19432 VSS.n13683 VSS.n13648 9.955
R19433 VSS.n13677 VSS.n13651 9.955
R19434 VSS.n13672 VSS.n13654 9.955
R19435 VSS.n13666 VSS.n13657 9.955
R19436 VSS.n13799 VSS.n10558 9.955
R19437 VSS.n13792 VSS.n13791 9.955
R19438 VSS.n13731 VSS.n13728 9.955
R19439 VSS.n13779 VSS.n13734 9.955
R19440 VSS.n13773 VSS.n13738 9.955
R19441 VSS.n13767 VSS.n13741 9.955
R19442 VSS.n13762 VSS.n13744 9.955
R19443 VSS.n13756 VSS.n13747 9.955
R19444 VSS.n13893 VSS.n13891 9.955
R19445 VSS.n13949 VSS.n10515 9.955
R19446 VSS.n13942 VSS.n13941 9.955
R19447 VSS.n13903 VSS.n13900 9.955
R19448 VSS.n13929 VSS.n13906 9.955
R19449 VSS.n13923 VSS.n13910 9.955
R19450 VSS.n13917 VSS.n13915 9.955
R19451 VSS.n13957 VSS.n13956 9.955
R19452 VSS.n9039 VSS.n9038 9.955
R19453 VSS.n9047 VSS.n9046 9.955
R19454 VSS.n9055 VSS.n9054 9.955
R19455 VSS.n9063 VSS.n9062 9.955
R19456 VSS.n9071 VSS.n9070 9.955
R19457 VSS.n9079 VSS.n9078 9.955
R19458 VSS.n9087 VSS.n9086 9.955
R19459 VSS.n9095 VSS.n9094 9.955
R19460 VSS.n10256 VSS.n9226 9.955
R19461 VSS.n10249 VSS.n10248 9.955
R19462 VSS.n10189 VSS.n10186 9.955
R19463 VSS.n10236 VSS.n10192 9.955
R19464 VSS.n10230 VSS.n10196 9.955
R19465 VSS.n10224 VSS.n10200 9.955
R19466 VSS.n10218 VSS.n10203 9.955
R19467 VSS.n10213 VSS.n10206 9.955
R19468 VSS.n10166 VSS.n9316 9.955
R19469 VSS.n10159 VSS.n10158 9.955
R19470 VSS.n10099 VSS.n10096 9.955
R19471 VSS.n10146 VSS.n10102 9.955
R19472 VSS.n10140 VSS.n10106 9.955
R19473 VSS.n10134 VSS.n10110 9.955
R19474 VSS.n10128 VSS.n10113 9.955
R19475 VSS.n10123 VSS.n10116 9.955
R19476 VSS.n10076 VSS.n9406 9.955
R19477 VSS.n10069 VSS.n10068 9.955
R19478 VSS.n10009 VSS.n10006 9.955
R19479 VSS.n10056 VSS.n10012 9.955
R19480 VSS.n10050 VSS.n10016 9.955
R19481 VSS.n10044 VSS.n10020 9.955
R19482 VSS.n10038 VSS.n10023 9.955
R19483 VSS.n10033 VSS.n10026 9.955
R19484 VSS.n9986 VSS.n9496 9.955
R19485 VSS.n9979 VSS.n9978 9.955
R19486 VSS.n9919 VSS.n9916 9.955
R19487 VSS.n9966 VSS.n9922 9.955
R19488 VSS.n9960 VSS.n9926 9.955
R19489 VSS.n9954 VSS.n9930 9.955
R19490 VSS.n9948 VSS.n9933 9.955
R19491 VSS.n9943 VSS.n9936 9.955
R19492 VSS.n9896 VSS.n9586 9.955
R19493 VSS.n9889 VSS.n9888 9.955
R19494 VSS.n9829 VSS.n9826 9.955
R19495 VSS.n9876 VSS.n9832 9.955
R19496 VSS.n9870 VSS.n9836 9.955
R19497 VSS.n9864 VSS.n9840 9.955
R19498 VSS.n9858 VSS.n9843 9.955
R19499 VSS.n9853 VSS.n9846 9.955
R19500 VSS.n9806 VSS.n9676 9.955
R19501 VSS.n9799 VSS.n9798 9.955
R19502 VSS.n9739 VSS.n9736 9.955
R19503 VSS.n9786 VSS.n9742 9.955
R19504 VSS.n9780 VSS.n9746 9.955
R19505 VSS.n9774 VSS.n9750 9.955
R19506 VSS.n9768 VSS.n9753 9.955
R19507 VSS.n9763 VSS.n9756 9.955
R19508 VSS.n9185 VSS.n9184 9.955
R19509 VSS.n10365 VSS.n8937 9.955
R19510 VSS.n10359 VSS.n8942 9.955
R19511 VSS.n10353 VSS.n8948 9.955
R19512 VSS.n10347 VSS.n8954 9.955
R19513 VSS.n10341 VSS.n8959 9.955
R19514 VSS.n10335 VSS.n8966 9.955
R19515 VSS.n10329 VSS.n8972 9.955
R19516 VSS.n5780 VSS.n3584 9.955
R19517 VSS.n5774 VSS.n3589 9.955
R19518 VSS.n5768 VSS.n3595 9.955
R19519 VSS.n5762 VSS.n3601 9.955
R19520 VSS.n5756 VSS.n3607 9.955
R19521 VSS.n5750 VSS.n3612 9.955
R19522 VSS.n5744 VSS.n3619 9.955
R19523 VSS.n5738 VSS.n3625 9.955
R19524 VSS.n5902 VSS.n3526 9.955
R19525 VSS.n5896 VSS.n3531 9.955
R19526 VSS.n5890 VSS.n3537 9.955
R19527 VSS.n5884 VSS.n3543 9.955
R19528 VSS.n5878 VSS.n3549 9.955
R19529 VSS.n5872 VSS.n3554 9.955
R19530 VSS.n5866 VSS.n3561 9.955
R19531 VSS.n5860 VSS.n3567 9.955
R19532 VSS.n6024 VSS.n3468 9.955
R19533 VSS.n6018 VSS.n3473 9.955
R19534 VSS.n6012 VSS.n3479 9.955
R19535 VSS.n6006 VSS.n3485 9.955
R19536 VSS.n6000 VSS.n3491 9.955
R19537 VSS.n5994 VSS.n3496 9.955
R19538 VSS.n5988 VSS.n3503 9.955
R19539 VSS.n5982 VSS.n3509 9.955
R19540 VSS.n6146 VSS.n3410 9.955
R19541 VSS.n6140 VSS.n3415 9.955
R19542 VSS.n6134 VSS.n3421 9.955
R19543 VSS.n6128 VSS.n3427 9.955
R19544 VSS.n6122 VSS.n3433 9.955
R19545 VSS.n6116 VSS.n3438 9.955
R19546 VSS.n6110 VSS.n3445 9.955
R19547 VSS.n6104 VSS.n3451 9.955
R19548 VSS.n6268 VSS.n3352 9.955
R19549 VSS.n6262 VSS.n3357 9.955
R19550 VSS.n6256 VSS.n3363 9.955
R19551 VSS.n6250 VSS.n3369 9.955
R19552 VSS.n6244 VSS.n3375 9.955
R19553 VSS.n6238 VSS.n3380 9.955
R19554 VSS.n6232 VSS.n3387 9.955
R19555 VSS.n6226 VSS.n3393 9.955
R19556 VSS.n6390 VSS.n3294 9.955
R19557 VSS.n6384 VSS.n3299 9.955
R19558 VSS.n6378 VSS.n3305 9.955
R19559 VSS.n6372 VSS.n3311 9.955
R19560 VSS.n6366 VSS.n3317 9.955
R19561 VSS.n6360 VSS.n3322 9.955
R19562 VSS.n6354 VSS.n3329 9.955
R19563 VSS.n6348 VSS.n3335 9.955
R19564 VSS.n6512 VSS.n3236 9.955
R19565 VSS.n6506 VSS.n3241 9.955
R19566 VSS.n6500 VSS.n3247 9.955
R19567 VSS.n6494 VSS.n3253 9.955
R19568 VSS.n6488 VSS.n3259 9.955
R19569 VSS.n6482 VSS.n3264 9.955
R19570 VSS.n6476 VSS.n3271 9.955
R19571 VSS.n6470 VSS.n3277 9.955
R19572 VSS.n6602 VSS.n6601 9.955
R19573 VSS.n3179 VSS.n3178 9.955
R19574 VSS.n3187 VSS.n3186 9.955
R19575 VSS.n3195 VSS.n3194 9.955
R19576 VSS.n3203 VSS.n3202 9.955
R19577 VSS.n3211 VSS.n3210 9.955
R19578 VSS.n3219 VSS.n3218 9.955
R19579 VSS.n3227 VSS.n3226 9.955
R19580 VSS.n1249 VSS.n43 9.955
R19581 VSS.n1242 VSS.n1241 9.955
R19582 VSS.n1187 VSS.n1184 9.955
R19583 VSS.n1229 VSS.n1190 9.955
R19584 VSS.n1223 VSS.n1194 9.955
R19585 VSS.n1217 VSS.n1198 9.955
R19586 VSS.n1211 VSS.n1201 9.955
R19587 VSS.n1206 VSS.n1204 9.955
R19588 VSS.n1164 VSS.n134 9.955
R19589 VSS.n1157 VSS.n1156 9.955
R19590 VSS.n1097 VSS.n1094 9.955
R19591 VSS.n1144 VSS.n1100 9.955
R19592 VSS.n1138 VSS.n1104 9.955
R19593 VSS.n1132 VSS.n1108 9.955
R19594 VSS.n1126 VSS.n1111 9.955
R19595 VSS.n1121 VSS.n1114 9.955
R19596 VSS.n1074 VSS.n224 9.955
R19597 VSS.n1067 VSS.n1066 9.955
R19598 VSS.n1007 VSS.n1004 9.955
R19599 VSS.n1054 VSS.n1010 9.955
R19600 VSS.n1048 VSS.n1014 9.955
R19601 VSS.n1042 VSS.n1018 9.955
R19602 VSS.n1036 VSS.n1021 9.955
R19603 VSS.n1031 VSS.n1024 9.955
R19604 VSS.n984 VSS.n314 9.955
R19605 VSS.n977 VSS.n976 9.955
R19606 VSS.n917 VSS.n914 9.955
R19607 VSS.n964 VSS.n920 9.955
R19608 VSS.n958 VSS.n924 9.955
R19609 VSS.n952 VSS.n928 9.955
R19610 VSS.n946 VSS.n931 9.955
R19611 VSS.n941 VSS.n934 9.955
R19612 VSS.n894 VSS.n404 9.955
R19613 VSS.n887 VSS.n886 9.955
R19614 VSS.n827 VSS.n824 9.955
R19615 VSS.n874 VSS.n830 9.955
R19616 VSS.n868 VSS.n834 9.955
R19617 VSS.n862 VSS.n838 9.955
R19618 VSS.n856 VSS.n841 9.955
R19619 VSS.n851 VSS.n844 9.955
R19620 VSS.n804 VSS.n494 9.955
R19621 VSS.n797 VSS.n796 9.955
R19622 VSS.n737 VSS.n734 9.955
R19623 VSS.n784 VSS.n740 9.955
R19624 VSS.n778 VSS.n744 9.955
R19625 VSS.n772 VSS.n748 9.955
R19626 VSS.n766 VSS.n751 9.955
R19627 VSS.n761 VSS.n754 9.955
R19628 VSS.n714 VSS.n584 9.955
R19629 VSS.n707 VSS.n706 9.955
R19630 VSS.n647 VSS.n644 9.955
R19631 VSS.n694 VSS.n650 9.955
R19632 VSS.n688 VSS.n654 9.955
R19633 VSS.n682 VSS.n658 9.955
R19634 VSS.n676 VSS.n661 9.955
R19635 VSS.n671 VSS.n664 9.955
R19636 VSS.n17600 sky130_asc_res_xhigh_po_2p85_1_19/VGND 9.905
R19637 sky130_asc_res_xhigh_po_2p85_1_8/VGND VSS.n10372 9.523
R19638 VSS.n16014 VSS.n16013 9.3
R19639 VSS.n16014 VSS.n14003 9.3
R19640 VSS.n14003 VSS.n14002 9.3
R19641 VSS.n14007 VSS.n14006 9.3
R19642 VSS.n16022 VSS.n16021 9.3
R19643 VSS.n16021 VSS.n16020 9.3
R19644 VSS.n16020 VSS.n16019 9.3
R19645 VSS.n15733 VSS.n15724 9.3
R19646 VSS.n15734 VSS.n15733 9.3
R19647 VSS.n15735 VSS.n15734 9.3
R19648 VSS.n15741 VSS.n15740 9.3
R19649 VSS.n15744 VSS.n15743 9.3
R19650 VSS.n15744 VSS.n15719 9.3
R19651 VSS.n15719 VSS.n15718 9.3
R19652 VSS.n15751 sky130_asc_pnp_05v5_W3p40L3p40_8_3/xm1/Collector 9.3
R19653 sky130_asc_pnp_05v5_W3p40L3p40_8_3/xm1/Collector VSS.n15750 9.3
R19654 VSS.n15750 VSS.n15749 9.3
R19655 VSS.n15752 VSS.n15710 9.3
R19656 VSS.n15755 VSS.n15705 9.3
R19657 VSS.n15756 VSS.n15755 9.3
R19658 VSS.n15757 VSS.n15756 9.3
R19659 VSS.n15766 VSS.n15765 9.3
R19660 VSS.n15766 VSS.n15700 9.3
R19661 VSS.n15700 VSS.n15699 9.3
R19662 VSS.n15704 VSS.n15703 9.3
R19663 VSS.n15774 VSS.n15773 9.3
R19664 VSS.n15773 VSS.n15772 9.3
R19665 VSS.n15772 VSS.n15771 9.3
R19666 VSS.n15778 VSS.n15686 9.3
R19667 VSS.n15779 VSS.n15778 9.3
R19668 VSS.n15780 VSS.n15779 9.3
R19669 VSS.n15786 VSS.n15785 9.3
R19670 VSS.n15789 VSS.n15788 9.3
R19671 VSS.n15789 VSS.n15681 9.3
R19672 VSS.n15681 VSS.n15680 9.3
R19673 VSS.n15797 VSS.n15796 9.3
R19674 VSS.n15796 VSS.n15795 9.3
R19675 VSS.n15795 VSS.n15794 9.3
R19676 VSS.n16011 VSS.n16010 9.3
R19677 VSS.n15730 VSS.n13995 9.3
R19678 VSS.n15723 VSS.n15722 9.3
R19679 VSS.n15763 VSS.n15762 9.3
R19680 VSS.n15775 VSS.n15691 9.3
R19681 VSS.n15685 VSS.n15684 9.3
R19682 VSS.n15799 VSS.n15636 9.3
R19683 VSS.n15802 VSS.n15631 9.3
R19684 VSS.n15803 VSS.n15802 9.3
R19685 VSS.n15804 VSS.n15803 9.3
R19686 VSS.n15810 VSS.n15809 9.3
R19687 VSS.n15813 VSS.n15812 9.3
R19688 VSS.n15813 VSS.n15626 9.3
R19689 VSS.n15626 VSS.n15625 9.3
R19690 VSS.n15630 VSS.n15629 9.3
R19691 VSS.n15821 VSS.n15820 9.3
R19692 VSS.n15820 VSS.n15819 9.3
R19693 VSS.n15819 VSS.n15818 9.3
R19694 VSS.n15822 VSS.n15617 9.3
R19695 VSS.n15825 VSS.n15612 9.3
R19696 VSS.n15826 VSS.n15825 9.3
R19697 VSS.n15827 VSS.n15826 9.3
R19698 VSS.n15833 VSS.n15832 9.3
R19699 VSS.n15836 VSS.n15835 9.3
R19700 VSS.n15836 VSS.n15607 9.3
R19701 VSS.n15607 VSS.n15606 9.3
R19702 VSS.n15611 VSS.n15610 9.3
R19703 VSS.n15843 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector 9.3
R19704 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector VSS.n15842 9.3
R19705 VSS.n15842 VSS.n15841 9.3
R19706 VSS.n15844 VSS.n15598 9.3
R19707 VSS.n15847 VSS.n15593 9.3
R19708 VSS.n15848 VSS.n15847 9.3
R19709 VSS.n15849 VSS.n15848 9.3
R19710 VSS.n15855 VSS.n15854 9.3
R19711 VSS.n15858 VSS.n15857 9.3
R19712 VSS.n15858 VSS.n15588 9.3
R19713 VSS.n15588 VSS.n15587 9.3
R19714 VSS.n15592 VSS.n15591 9.3
R19715 VSS.n15866 VSS.n15865 9.3
R19716 VSS.n15865 VSS.n15864 9.3
R19717 VSS.n15864 VSS.n15863 9.3
R19718 VSS.n15867 VSS.n15579 9.3
R19719 VSS.n15870 VSS.n15574 9.3
R19720 VSS.n15871 VSS.n15870 9.3
R19721 VSS.n15872 VSS.n15871 9.3
R19722 VSS.n15878 VSS.n15877 9.3
R19723 VSS.n15881 VSS.n15880 9.3
R19724 VSS.n15881 VSS.n15569 9.3
R19725 VSS.n15569 VSS.n15568 9.3
R19726 VSS.n15573 VSS.n15572 9.3
R19727 VSS.n15889 VSS.n15888 9.3
R19728 VSS.n15888 VSS.n15887 9.3
R19729 VSS.n15887 VSS.n15886 9.3
R19730 VSS.n15559 VSS.n14072 9.3
R19731 VSS.n15556 VSS.n14073 9.3
R19732 VSS.n15556 VSS.n15555 9.3
R19733 VSS.n15555 VSS.n15554 9.3
R19734 VSS.n15549 VSS.n15548 9.3
R19735 VSS.n15546 VSS.n15545 9.3
R19736 VSS.n15545 VSS.n14077 9.3
R19737 VSS.n14077 VSS.n14076 9.3
R19738 VSS.n14085 VSS.n14079 9.3
R19739 VSS.n15538 VSS.n15537 9.3
R19740 VSS.n15539 VSS.n15538 9.3
R19741 VSS.n15540 VSS.n15539 9.3
R19742 VSS.n15535 VSS.n15534 9.3
R19743 VSS.n15526 VSS.n15525 9.3
R19744 VSS.n15526 VSS.n14089 9.3
R19745 VSS.n15530 VSS.n14089 9.3
R19746 VSS.n15524 VSS.n15523 9.3
R19747 VSS.n15521 VSS.n14095 9.3
R19748 VSS.n15521 VSS.n15520 9.3
R19749 VSS.n15520 VSS.n15519 9.3
R19750 VSS.n15514 VSS.n15513 9.3
R19751 VSS.n15511 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector 9.3
R19752 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector VSS.n14098 9.3
R19753 VSS.n14098 VSS.n14097 9.3
R19754 VSS.n14106 VSS.n14100 9.3
R19755 VSS.n15504 VSS.n15503 9.3
R19756 VSS.n15505 VSS.n15504 9.3
R19757 VSS.n15506 VSS.n15505 9.3
R19758 VSS.n15501 VSS.n15500 9.3
R19759 VSS.n15492 VSS.n15491 9.3
R19760 VSS.n15492 VSS.n14110 9.3
R19761 VSS.n15496 VSS.n14110 9.3
R19762 VSS.n15490 VSS.n15489 9.3
R19763 VSS.n15487 VSS.n14116 9.3
R19764 VSS.n15487 VSS.n15486 9.3
R19765 VSS.n15486 VSS.n15485 9.3
R19766 VSS.n15480 VSS.n15479 9.3
R19767 VSS.n15477 VSS.n15476 9.3
R19768 VSS.n15476 VSS.n14119 9.3
R19769 VSS.n14119 VSS.n14118 9.3
R19770 VSS.n14127 VSS.n14121 9.3
R19771 VSS.n15469 VSS.n15468 9.3
R19772 VSS.n15470 VSS.n15469 9.3
R19773 VSS.n15471 VSS.n15470 9.3
R19774 VSS.n15466 VSS.n15465 9.3
R19775 VSS.n15457 VSS.n15456 9.3
R19776 VSS.n15457 VSS.n14131 9.3
R19777 VSS.n15461 VSS.n14131 9.3
R19778 VSS.n15453 VSS.n14135 9.3
R19779 VSS.n15450 VSS.n14137 9.3
R19780 VSS.n15442 VSS.n14137 9.3
R19781 VSS.n15443 VSS.n15442 9.3
R19782 VSS.n15449 VSS.n15448 9.3
R19783 VSS.n15154 VSS.n15153 9.3
R19784 VSS.n15154 VSS.n14141 9.3
R19785 VSS.n14143 VSS.n14141 9.3
R19786 VSS.n15152 VSS.n15151 9.3
R19787 VSS.n15162 VSS.n15161 9.3
R19788 VSS.n15161 VSS.n15160 9.3
R19789 VSS.n15160 VSS.n15159 9.3
R19790 VSS.n15163 VSS.n15142 9.3
R19791 VSS.n15166 VSS.n15137 9.3
R19792 VSS.n15167 VSS.n15166 9.3
R19793 VSS.n15168 VSS.n15167 9.3
R19794 VSS.n15174 VSS.n15173 9.3
R19795 VSS.n15177 VSS.n15176 9.3
R19796 VSS.n15177 VSS.n15132 9.3
R19797 VSS.n15132 VSS.n15131 9.3
R19798 VSS.n15136 VSS.n15135 9.3
R19799 VSS.n15184 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector 9.3
R19800 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector VSS.n15183 9.3
R19801 VSS.n15183 VSS.n15182 9.3
R19802 VSS.n15185 VSS.n15123 9.3
R19803 VSS.n15188 VSS.n15118 9.3
R19804 VSS.n15189 VSS.n15188 9.3
R19805 VSS.n15190 VSS.n15189 9.3
R19806 VSS.n15196 VSS.n15195 9.3
R19807 VSS.n15199 VSS.n15198 9.3
R19808 VSS.n15199 VSS.n15113 9.3
R19809 VSS.n15113 VSS.n15112 9.3
R19810 VSS.n15117 VSS.n15116 9.3
R19811 VSS.n15207 VSS.n15206 9.3
R19812 VSS.n15206 VSS.n15205 9.3
R19813 VSS.n15205 VSS.n15204 9.3
R19814 VSS.n15208 VSS.n15104 9.3
R19815 VSS.n15211 VSS.n15099 9.3
R19816 VSS.n15212 VSS.n15211 9.3
R19817 VSS.n15213 VSS.n15212 9.3
R19818 VSS.n15219 VSS.n15218 9.3
R19819 VSS.n15222 VSS.n15221 9.3
R19820 VSS.n15222 VSS.n15094 9.3
R19821 VSS.n15094 VSS.n15093 9.3
R19822 VSS.n15098 VSS.n15097 9.3
R19823 VSS.n15230 VSS.n15229 9.3
R19824 VSS.n15229 VSS.n15228 9.3
R19825 VSS.n15228 VSS.n15227 9.3
R19826 VSS.n15232 VSS.n15049 9.3
R19827 VSS.n15235 VSS.n15044 9.3
R19828 VSS.n15236 VSS.n15235 9.3
R19829 VSS.n15237 VSS.n15236 9.3
R19830 VSS.n15243 VSS.n15242 9.3
R19831 VSS.n15246 VSS.n15245 9.3
R19832 VSS.n15246 VSS.n15039 9.3
R19833 VSS.n15039 VSS.n15038 9.3
R19834 VSS.n15043 VSS.n15042 9.3
R19835 VSS.n15254 VSS.n15253 9.3
R19836 VSS.n15253 VSS.n15252 9.3
R19837 VSS.n15252 VSS.n15251 9.3
R19838 VSS.n15255 VSS.n15030 9.3
R19839 VSS.n15258 VSS.n15025 9.3
R19840 VSS.n15259 VSS.n15258 9.3
R19841 VSS.n15260 VSS.n15259 9.3
R19842 VSS.n15266 VSS.n15265 9.3
R19843 VSS.n15269 VSS.n15268 9.3
R19844 VSS.n15269 VSS.n15020 9.3
R19845 VSS.n15020 VSS.n15019 9.3
R19846 VSS.n15024 VSS.n15023 9.3
R19847 VSS.n15276 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector 9.3
R19848 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector VSS.n15275 9.3
R19849 VSS.n15275 VSS.n15274 9.3
R19850 VSS.n15277 VSS.n15011 9.3
R19851 VSS.n15280 VSS.n15006 9.3
R19852 VSS.n15281 VSS.n15280 9.3
R19853 VSS.n15282 VSS.n15281 9.3
R19854 VSS.n15288 VSS.n15287 9.3
R19855 VSS.n15291 VSS.n15290 9.3
R19856 VSS.n15291 VSS.n15001 9.3
R19857 VSS.n15001 VSS.n15000 9.3
R19858 VSS.n15005 VSS.n15004 9.3
R19859 VSS.n15299 VSS.n15298 9.3
R19860 VSS.n15298 VSS.n15297 9.3
R19861 VSS.n15297 VSS.n15296 9.3
R19862 VSS.n15300 VSS.n14992 9.3
R19863 VSS.n15303 VSS.n14987 9.3
R19864 VSS.n15304 VSS.n15303 9.3
R19865 VSS.n15305 VSS.n15304 9.3
R19866 VSS.n15311 VSS.n15310 9.3
R19867 VSS.n15314 VSS.n15313 9.3
R19868 VSS.n15314 VSS.n14982 9.3
R19869 VSS.n14982 VSS.n14981 9.3
R19870 VSS.n14986 VSS.n14985 9.3
R19871 VSS.n15322 VSS.n15321 9.3
R19872 VSS.n15321 VSS.n15320 9.3
R19873 VSS.n15320 VSS.n15319 9.3
R19874 VSS.n15325 VSS.n15324 9.3
R19875 VSS.n15328 VSS.n15327 9.3
R19876 VSS.n15329 VSS.n15328 9.3
R19877 VSS.n15330 VSS.n15329 9.3
R19878 VSS.n14972 VSS.n14971 9.3
R19879 VSS.n14963 VSS.n14962 9.3
R19880 VSS.n14963 VSS.n14245 9.3
R19881 VSS.n14967 VSS.n14245 9.3
R19882 VSS.n14961 VSS.n14960 9.3
R19883 VSS.n14958 VSS.n14251 9.3
R19884 VSS.n14958 VSS.n14957 9.3
R19885 VSS.n14957 VSS.n14956 9.3
R19886 VSS.n14951 VSS.n14950 9.3
R19887 VSS.n14948 VSS.n14947 9.3
R19888 VSS.n14947 VSS.n14254 9.3
R19889 VSS.n14254 VSS.n14253 9.3
R19890 VSS.n14262 VSS.n14256 9.3
R19891 VSS.n14940 VSS.n14939 9.3
R19892 VSS.n14941 VSS.n14940 9.3
R19893 VSS.n14942 VSS.n14941 9.3
R19894 VSS.n14937 VSS.n14936 9.3
R19895 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector VSS.n14928 9.3
R19896 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector VSS.n14266 9.3
R19897 VSS.n14932 VSS.n14266 9.3
R19898 VSS.n14927 VSS.n14926 9.3
R19899 VSS.n14924 VSS.n14272 9.3
R19900 VSS.n14924 VSS.n14923 9.3
R19901 VSS.n14923 VSS.n14922 9.3
R19902 VSS.n14917 VSS.n14916 9.3
R19903 VSS.n14914 VSS.n14913 9.3
R19904 VSS.n14913 VSS.n14275 9.3
R19905 VSS.n14275 VSS.n14274 9.3
R19906 VSS.n14283 VSS.n14277 9.3
R19907 VSS.n14906 VSS.n14905 9.3
R19908 VSS.n14907 VSS.n14906 9.3
R19909 VSS.n14908 VSS.n14907 9.3
R19910 VSS.n14903 VSS.n14902 9.3
R19911 VSS.n14894 VSS.n14893 9.3
R19912 VSS.n14894 VSS.n14287 9.3
R19913 VSS.n14898 VSS.n14287 9.3
R19914 VSS.n14892 VSS.n14891 9.3
R19915 VSS.n14889 VSS.n14293 9.3
R19916 VSS.n14889 VSS.n14888 9.3
R19917 VSS.n14888 VSS.n14887 9.3
R19918 VSS.n14882 VSS.n14881 9.3
R19919 VSS.n14879 VSS.n14878 9.3
R19920 VSS.n14878 VSS.n14296 9.3
R19921 VSS.n14296 VSS.n14295 9.3
R19922 VSS.n14867 VSS.n14866 9.3
R19923 VSS.n14870 VSS.n14869 9.3
R19924 VSS.n14871 VSS.n14870 9.3
R19925 VSS.n14872 VSS.n14871 9.3
R19926 VSS.n14547 VSS.n14307 9.3
R19927 VSS.n14553 VSS.n14552 9.3
R19928 VSS.n14553 VSS.n14542 9.3
R19929 VSS.n14542 VSS.n14541 9.3
R19930 VSS.n14550 VSS.n14549 9.3
R19931 VSS.n14561 VSS.n14560 9.3
R19932 VSS.n14560 VSS.n14559 9.3
R19933 VSS.n14559 VSS.n14558 9.3
R19934 VSS.n14562 VSS.n14533 9.3
R19935 VSS.n14565 VSS.n14528 9.3
R19936 VSS.n14566 VSS.n14565 9.3
R19937 VSS.n14567 VSS.n14566 9.3
R19938 VSS.n14573 VSS.n14572 9.3
R19939 VSS.n14576 VSS.n14575 9.3
R19940 VSS.n14576 VSS.n14523 9.3
R19941 VSS.n14523 VSS.n14522 9.3
R19942 VSS.n14527 VSS.n14526 9.3
R19943 VSS.n14583 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector 9.3
R19944 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector VSS.n14582 9.3
R19945 VSS.n14582 VSS.n14581 9.3
R19946 VSS.n14584 VSS.n14514 9.3
R19947 VSS.n14587 VSS.n14509 9.3
R19948 VSS.n14588 VSS.n14587 9.3
R19949 VSS.n14589 VSS.n14588 9.3
R19950 VSS.n14595 VSS.n14594 9.3
R19951 VSS.n14598 VSS.n14597 9.3
R19952 VSS.n14598 VSS.n14504 9.3
R19953 VSS.n14504 VSS.n14503 9.3
R19954 VSS.n14508 VSS.n14507 9.3
R19955 VSS.n14606 VSS.n14605 9.3
R19956 VSS.n14605 VSS.n14604 9.3
R19957 VSS.n14604 VSS.n14603 9.3
R19958 VSS.n14607 VSS.n14495 9.3
R19959 VSS.n14610 VSS.n14490 9.3
R19960 VSS.n14611 VSS.n14610 9.3
R19961 VSS.n14612 VSS.n14611 9.3
R19962 VSS.n14618 VSS.n14617 9.3
R19963 VSS.n14621 VSS.n14620 9.3
R19964 VSS.n14621 VSS.n14485 9.3
R19965 VSS.n14485 VSS.n14484 9.3
R19966 VSS.n14489 VSS.n14488 9.3
R19967 VSS.n14629 VSS.n14628 9.3
R19968 VSS.n14628 VSS.n14627 9.3
R19969 VSS.n14627 VSS.n14626 9.3
R19970 VSS.n14631 VSS.n14440 9.3
R19971 VSS.n14634 VSS.n14435 9.3
R19972 VSS.n14635 VSS.n14634 9.3
R19973 VSS.n14636 VSS.n14635 9.3
R19974 VSS.n14642 VSS.n14641 9.3
R19975 VSS.n14645 VSS.n14644 9.3
R19976 VSS.n14645 VSS.n14430 9.3
R19977 VSS.n14430 VSS.n14429 9.3
R19978 VSS.n14434 VSS.n14433 9.3
R19979 VSS.n14653 VSS.n14652 9.3
R19980 VSS.n14652 VSS.n14651 9.3
R19981 VSS.n14651 VSS.n14650 9.3
R19982 VSS.n14654 VSS.n14421 9.3
R19983 VSS.n14657 VSS.n14416 9.3
R19984 VSS.n14658 VSS.n14657 9.3
R19985 VSS.n14659 VSS.n14658 9.3
R19986 VSS.n14665 VSS.n14664 9.3
R19987 VSS.n14668 VSS.n14667 9.3
R19988 VSS.n14668 VSS.n14411 9.3
R19989 VSS.n14411 VSS.n14410 9.3
R19990 VSS.n14415 VSS.n14414 9.3
R19991 VSS.n14675 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Collector 9.3
R19992 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Collector VSS.n14674 9.3
R19993 VSS.n14674 VSS.n14673 9.3
R19994 VSS.n14676 VSS.n14402 9.3
R19995 VSS.n14679 VSS.n14397 9.3
R19996 VSS.n14680 VSS.n14679 9.3
R19997 VSS.n14681 VSS.n14680 9.3
R19998 VSS.n14687 VSS.n14686 9.3
R19999 VSS.n14690 VSS.n14689 9.3
R20000 VSS.n14690 VSS.n14392 9.3
R20001 VSS.n14392 VSS.n14391 9.3
R20002 VSS.n14396 VSS.n14395 9.3
R20003 VSS.n14698 VSS.n14697 9.3
R20004 VSS.n14697 VSS.n14696 9.3
R20005 VSS.n14696 VSS.n14695 9.3
R20006 VSS.n14699 VSS.n14383 9.3
R20007 VSS.n14702 VSS.n14378 9.3
R20008 VSS.n14703 VSS.n14702 9.3
R20009 VSS.n14704 VSS.n14703 9.3
R20010 VSS.n14710 VSS.n14709 9.3
R20011 VSS.n14713 VSS.n14712 9.3
R20012 VSS.n14713 VSS.n14372 9.3
R20013 VSS.n14372 VSS.n14371 9.3
R20014 VSS.n14377 VSS.n14376 9.3
R20015 VSS.n14720 VSS.n14369 9.3
R20016 VSS.n14720 VSS.n14719 9.3
R20017 VSS.n14719 VSS.n14718 9.3
R20018 VSS.n16003 VSS.n14008 9.3
R20019 VSS.n16004 VSS.n16003 9.3
R20020 VSS.n16005 VSS.n16004 9.3
R20021 VSS.n16000 VSS.n14013 9.3
R20022 VSS.n16721 VSS.n16720 9.3
R20023 VSS.n16720 VSS.n16620 9.3
R20024 VSS.n16723 VSS.n16722 9.3
R20025 VSS.n16727 VSS.n16726 9.3
R20026 VSS.n16726 VSS.n16725 9.3
R20027 VSS.n16733 VSS.n16732 9.3
R20028 VSS.n16732 VSS.n16731 9.3
R20029 VSS.n16735 VSS.n16734 9.3
R20030 VSS.n16739 VSS.n16738 9.3
R20031 VSS.n16738 VSS.n16737 9.3
R20032 VSS.n16745 VSS.n16744 9.3
R20033 VSS.n16744 VSS.n16743 9.3
R20034 VSS.n16746 VSS.n16691 9.3
R20035 VSS.n16750 VSS.n16690 9.3
R20036 VSS.n16750 VSS.n16749 9.3
R20037 VSS.n16759 VSS.n16757 9.3
R20038 VSS.n16759 VSS.n16758 9.3
R20039 VSS.n16689 VSS.n16631 9.3
R20040 VSS.n16686 VSS.n16633 9.3
R20041 VSS.n16686 VSS.n16630 9.3
R20042 VSS.n16718 VSS.n16717 9.3
R20043 VSS.n16729 VSS.n16728 9.3
R20044 VSS.n16741 VSS.n16740 9.3
R20045 VSS.n16755 VSS.n16754 9.3
R20046 VSS.n16716 VSS.n16715 9.3
R20047 VSS.n16715 VSS.n16595 9.3
R20048 VSS.n16593 VSS.n16592 9.3
R20049 VSS.n16811 VSS.n16810 9.3
R20050 VSS.n16810 VSS.n16530 9.3
R20051 VSS.n16813 VSS.n16812 9.3
R20052 VSS.n16817 VSS.n16816 9.3
R20053 VSS.n16816 VSS.n16815 9.3
R20054 VSS.n16823 VSS.n16822 9.3
R20055 VSS.n16822 VSS.n16821 9.3
R20056 VSS.n16825 VSS.n16824 9.3
R20057 VSS.n16829 VSS.n16828 9.3
R20058 VSS.n16828 VSS.n16827 9.3
R20059 VSS.n16835 VSS.n16834 9.3
R20060 VSS.n16834 VSS.n16833 9.3
R20061 VSS.n16836 VSS.n16781 9.3
R20062 VSS.n16840 VSS.n16780 9.3
R20063 VSS.n16840 VSS.n16839 9.3
R20064 VSS.n16849 VSS.n16847 9.3
R20065 VSS.n16849 VSS.n16848 9.3
R20066 VSS.n16779 VSS.n16541 9.3
R20067 VSS.n16776 VSS.n16543 9.3
R20068 VSS.n16776 VSS.n16540 9.3
R20069 VSS.n16808 VSS.n16807 9.3
R20070 VSS.n16819 VSS.n16818 9.3
R20071 VSS.n16831 VSS.n16830 9.3
R20072 VSS.n16845 VSS.n16844 9.3
R20073 VSS.n16806 VSS.n16805 9.3
R20074 VSS.n16805 VSS.n16505 9.3
R20075 VSS.n16503 VSS.n16502 9.3
R20076 VSS.n16901 VSS.n16900 9.3
R20077 VSS.n16900 VSS.n16440 9.3
R20078 VSS.n16903 VSS.n16902 9.3
R20079 VSS.n16907 VSS.n16906 9.3
R20080 VSS.n16906 VSS.n16905 9.3
R20081 VSS.n16913 VSS.n16912 9.3
R20082 VSS.n16912 VSS.n16911 9.3
R20083 VSS.n16915 VSS.n16914 9.3
R20084 VSS.n16919 VSS.n16918 9.3
R20085 VSS.n16918 VSS.n16917 9.3
R20086 VSS.n16925 VSS.n16924 9.3
R20087 VSS.n16924 VSS.n16923 9.3
R20088 VSS.n16926 VSS.n16871 9.3
R20089 VSS.n16930 VSS.n16870 9.3
R20090 VSS.n16930 VSS.n16929 9.3
R20091 VSS.n16939 VSS.n16937 9.3
R20092 VSS.n16939 VSS.n16938 9.3
R20093 VSS.n16869 VSS.n16451 9.3
R20094 VSS.n16866 VSS.n16453 9.3
R20095 VSS.n16866 VSS.n16450 9.3
R20096 VSS.n16898 VSS.n16897 9.3
R20097 VSS.n16909 VSS.n16908 9.3
R20098 VSS.n16921 VSS.n16920 9.3
R20099 VSS.n16935 VSS.n16934 9.3
R20100 VSS.n16896 VSS.n16895 9.3
R20101 VSS.n16895 VSS.n16415 9.3
R20102 VSS.n16413 VSS.n16412 9.3
R20103 VSS.n16991 VSS.n16990 9.3
R20104 VSS.n16990 VSS.n16350 9.3
R20105 VSS.n16993 VSS.n16992 9.3
R20106 VSS.n16997 VSS.n16996 9.3
R20107 VSS.n16996 VSS.n16995 9.3
R20108 VSS.n17003 VSS.n17002 9.3
R20109 VSS.n17002 VSS.n17001 9.3
R20110 VSS.n17005 VSS.n17004 9.3
R20111 VSS.n17009 VSS.n17008 9.3
R20112 VSS.n17008 VSS.n17007 9.3
R20113 VSS.n17015 VSS.n17014 9.3
R20114 VSS.n17014 VSS.n17013 9.3
R20115 VSS.n17016 VSS.n16961 9.3
R20116 VSS.n17020 VSS.n16960 9.3
R20117 VSS.n17020 VSS.n17019 9.3
R20118 VSS.n17029 VSS.n17027 9.3
R20119 VSS.n17029 VSS.n17028 9.3
R20120 VSS.n16959 VSS.n16361 9.3
R20121 VSS.n16956 VSS.n16363 9.3
R20122 VSS.n16956 VSS.n16360 9.3
R20123 VSS.n16988 VSS.n16987 9.3
R20124 VSS.n16999 VSS.n16998 9.3
R20125 VSS.n17011 VSS.n17010 9.3
R20126 VSS.n17025 VSS.n17024 9.3
R20127 VSS.n16986 VSS.n16985 9.3
R20128 VSS.n16985 VSS.n16325 9.3
R20129 VSS.n16323 VSS.n16322 9.3
R20130 VSS.n17081 VSS.n17080 9.3
R20131 VSS.n17080 VSS.n16260 9.3
R20132 VSS.n17083 VSS.n17082 9.3
R20133 VSS.n17087 VSS.n17086 9.3
R20134 VSS.n17086 VSS.n17085 9.3
R20135 VSS.n17093 VSS.n17092 9.3
R20136 VSS.n17092 VSS.n17091 9.3
R20137 VSS.n17095 VSS.n17094 9.3
R20138 VSS.n17099 VSS.n17098 9.3
R20139 VSS.n17098 VSS.n17097 9.3
R20140 VSS.n17105 VSS.n17104 9.3
R20141 VSS.n17104 VSS.n17103 9.3
R20142 VSS.n17106 VSS.n17051 9.3
R20143 VSS.n17110 VSS.n17050 9.3
R20144 VSS.n17110 VSS.n17109 9.3
R20145 VSS.n17119 VSS.n17117 9.3
R20146 VSS.n17119 VSS.n17118 9.3
R20147 VSS.n17049 VSS.n16271 9.3
R20148 VSS.n17046 VSS.n16273 9.3
R20149 VSS.n17046 VSS.n16270 9.3
R20150 VSS.n17078 VSS.n17077 9.3
R20151 VSS.n17089 VSS.n17088 9.3
R20152 VSS.n17101 VSS.n17100 9.3
R20153 VSS.n17115 VSS.n17114 9.3
R20154 VSS.n17076 VSS.n17075 9.3
R20155 VSS.n17075 VSS.n16235 9.3
R20156 VSS.n16233 VSS.n16232 9.3
R20157 VSS.n17171 VSS.n17170 9.3
R20158 VSS.n17170 VSS.n16170 9.3
R20159 VSS.n17173 VSS.n17172 9.3
R20160 VSS.n17177 VSS.n17176 9.3
R20161 VSS.n17176 VSS.n17175 9.3
R20162 VSS.n17183 VSS.n17182 9.3
R20163 VSS.n17182 VSS.n17181 9.3
R20164 VSS.n17185 VSS.n17184 9.3
R20165 VSS.n17189 VSS.n17188 9.3
R20166 VSS.n17188 VSS.n17187 9.3
R20167 VSS.n17195 VSS.n17194 9.3
R20168 VSS.n17194 VSS.n17193 9.3
R20169 VSS.n17196 VSS.n17141 9.3
R20170 VSS.n17200 VSS.n17140 9.3
R20171 VSS.n17200 VSS.n17199 9.3
R20172 VSS.n17209 VSS.n17207 9.3
R20173 VSS.n17209 VSS.n17208 9.3
R20174 VSS.n17139 VSS.n16181 9.3
R20175 VSS.n17136 VSS.n16183 9.3
R20176 VSS.n17136 VSS.n16180 9.3
R20177 VSS.n17168 VSS.n17167 9.3
R20178 VSS.n17179 VSS.n17178 9.3
R20179 VSS.n17191 VSS.n17190 9.3
R20180 VSS.n17205 VSS.n17204 9.3
R20181 VSS.n17166 VSS.n17165 9.3
R20182 VSS.n17165 VSS.n16145 9.3
R20183 VSS.n16143 VSS.n16142 9.3
R20184 VSS.n17261 VSS.n17260 9.3
R20185 VSS.n17260 VSS.n16080 9.3
R20186 VSS.n17263 VSS.n17262 9.3
R20187 VSS.n17267 VSS.n17266 9.3
R20188 VSS.n17266 VSS.n17265 9.3
R20189 VSS.n17273 VSS.n17272 9.3
R20190 VSS.n17272 VSS.n17271 9.3
R20191 VSS.n17275 VSS.n17274 9.3
R20192 VSS.n17279 VSS.n17278 9.3
R20193 VSS.n17278 VSS.n17277 9.3
R20194 VSS.n17285 VSS.n17284 9.3
R20195 VSS.n17284 VSS.n17283 9.3
R20196 VSS.n17286 VSS.n17231 9.3
R20197 VSS.n17290 VSS.n17230 9.3
R20198 VSS.n17290 VSS.n17289 9.3
R20199 VSS.n17299 VSS.n17297 9.3
R20200 VSS.n17299 VSS.n17298 9.3
R20201 VSS.n17229 VSS.n16091 9.3
R20202 VSS.n17226 VSS.n16093 9.3
R20203 VSS.n17226 VSS.n16090 9.3
R20204 VSS.n17258 VSS.n17257 9.3
R20205 VSS.n17269 VSS.n17268 9.3
R20206 VSS.n17281 VSS.n17280 9.3
R20207 VSS.n17295 VSS.n17294 9.3
R20208 VSS.n17256 VSS.n17255 9.3
R20209 VSS.n17255 VSS.n16055 9.3
R20210 VSS.n16053 VSS.n16052 9.3
R20211 VSS.n17429 VSS.n17428 9.3
R20212 VSS.n17428 VSS.n17427 9.3
R20213 VSS.n17431 VSS.n17430 9.3
R20214 VSS.n17435 VSS.n17434 9.3
R20215 VSS.n17434 VSS.n17433 9.3
R20216 VSS.n17441 VSS.n17440 9.3
R20217 VSS.n17440 VSS.n17439 9.3
R20218 VSS.n17442 VSS.n17400 9.3
R20219 VSS.n17446 VSS.n17399 9.3
R20220 VSS.n17446 VSS.n17445 9.3
R20221 VSS.n17455 VSS.n17453 9.3
R20222 VSS.n17455 VSS.n17454 9.3
R20223 VSS.n17398 VSS.n16048 9.3
R20224 VSS.n17395 VSS.n16050 9.3
R20225 VSS.n17395 VSS.n16047 9.3
R20226 VSS.n17388 VSS.n17387 9.3
R20227 VSS.n17387 VSS.n17386 9.3
R20228 VSS.n17463 VSS.n17462 9.3
R20229 VSS.n17462 VSS.n17461 9.3
R20230 VSS.n17461 VSS.n17460 9.3
R20231 VSS.n17332 VSS.n17331 9.3
R20232 VSS.n17425 VSS.n17424 9.3
R20233 VSS.n17437 VSS.n17436 9.3
R20234 VSS.n17451 VSS.n17450 9.3
R20235 VSS.n17391 VSS.n17390 9.3
R20236 VSS.n17423 VSS.n17422 9.3
R20237 VSS.n17422 VSS.n17421 9.3
R20238 VSS.n17419 VSS.n17418 9.3
R20239 VSS.n12229 VSS.n12228 9.3
R20240 VSS.n12229 VSS.n12052 9.3
R20241 VSS.n12052 VSS.n12051 9.3
R20242 VSS.n12056 VSS.n12055 9.3
R20243 VSS.n12237 VSS.n12236 9.3
R20244 VSS.n12236 VSS.n12235 9.3
R20245 VSS.n12235 VSS.n12234 9.3
R20246 VSS.n12241 VSS.n12038 9.3
R20247 VSS.n12242 VSS.n12241 9.3
R20248 VSS.n12243 VSS.n12242 9.3
R20249 VSS.n12249 VSS.n12248 9.3
R20250 VSS.n12252 VSS.n12251 9.3
R20251 VSS.n12252 VSS.n12033 9.3
R20252 VSS.n12033 VSS.n12032 9.3
R20253 VSS.n12259 sky130_asc_pnp_05v5_W3p40L3p40_8_0/xm1/Collector 9.3
R20254 sky130_asc_pnp_05v5_W3p40L3p40_8_0/xm1/Collector VSS.n12258 9.3
R20255 VSS.n12258 VSS.n12257 9.3
R20256 VSS.n12260 VSS.n12024 9.3
R20257 VSS.n12263 VSS.n12019 9.3
R20258 VSS.n12264 VSS.n12263 9.3
R20259 VSS.n12265 VSS.n12264 9.3
R20260 VSS.n12274 VSS.n12273 9.3
R20261 VSS.n12274 VSS.n12014 9.3
R20262 VSS.n12014 VSS.n12013 9.3
R20263 VSS.n12018 VSS.n12017 9.3
R20264 VSS.n12282 VSS.n12281 9.3
R20265 VSS.n12281 VSS.n12280 9.3
R20266 VSS.n12280 VSS.n12279 9.3
R20267 VSS.n12286 VSS.n12000 9.3
R20268 VSS.n12287 VSS.n12286 9.3
R20269 VSS.n12288 VSS.n12287 9.3
R20270 VSS.n12294 VSS.n12293 9.3
R20271 VSS.n12297 VSS.n12296 9.3
R20272 VSS.n12297 VSS.n11995 9.3
R20273 VSS.n11995 VSS.n11994 9.3
R20274 VSS.n12305 VSS.n12304 9.3
R20275 VSS.n12304 VSS.n12303 9.3
R20276 VSS.n12303 VSS.n12302 9.3
R20277 VSS.n12226 VSS.n12225 9.3
R20278 VSS.n12238 VSS.n12043 9.3
R20279 VSS.n12037 VSS.n12036 9.3
R20280 VSS.n12271 VSS.n12270 9.3
R20281 VSS.n12283 VSS.n12005 9.3
R20282 VSS.n11999 VSS.n11998 9.3
R20283 VSS.n12307 VSS.n11983 9.3
R20284 VSS.n12310 VSS.n11978 9.3
R20285 VSS.n12311 VSS.n12310 9.3
R20286 VSS.n12312 VSS.n12311 9.3
R20287 VSS.n12318 VSS.n12317 9.3
R20288 VSS.n12321 VSS.n12320 9.3
R20289 VSS.n12321 VSS.n11973 9.3
R20290 VSS.n11973 VSS.n11972 9.3
R20291 VSS.n11977 VSS.n11976 9.3
R20292 VSS.n12329 VSS.n12328 9.3
R20293 VSS.n12328 VSS.n12327 9.3
R20294 VSS.n12327 VSS.n12326 9.3
R20295 VSS.n12330 VSS.n11964 9.3
R20296 VSS.n12333 VSS.n11959 9.3
R20297 VSS.n12334 VSS.n12333 9.3
R20298 VSS.n12335 VSS.n12334 9.3
R20299 VSS.n12341 VSS.n12340 9.3
R20300 VSS.n12344 VSS.n12343 9.3
R20301 VSS.n12344 VSS.n11954 9.3
R20302 VSS.n11954 VSS.n11953 9.3
R20303 VSS.n11958 VSS.n11957 9.3
R20304 VSS.n12351 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector 9.3
R20305 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector VSS.n12350 9.3
R20306 VSS.n12350 VSS.n12349 9.3
R20307 VSS.n12352 VSS.n11945 9.3
R20308 VSS.n12355 VSS.n11940 9.3
R20309 VSS.n12356 VSS.n12355 9.3
R20310 VSS.n12357 VSS.n12356 9.3
R20311 VSS.n12363 VSS.n12362 9.3
R20312 VSS.n12366 VSS.n12365 9.3
R20313 VSS.n12366 VSS.n11935 9.3
R20314 VSS.n11935 VSS.n11934 9.3
R20315 VSS.n11939 VSS.n11938 9.3
R20316 VSS.n12374 VSS.n12373 9.3
R20317 VSS.n12373 VSS.n12372 9.3
R20318 VSS.n12372 VSS.n12371 9.3
R20319 VSS.n12375 VSS.n11926 9.3
R20320 VSS.n12378 VSS.n11921 9.3
R20321 VSS.n12379 VSS.n12378 9.3
R20322 VSS.n12380 VSS.n12379 9.3
R20323 VSS.n12386 VSS.n12385 9.3
R20324 VSS.n12389 VSS.n12388 9.3
R20325 VSS.n12389 VSS.n11916 9.3
R20326 VSS.n11916 VSS.n11915 9.3
R20327 VSS.n11920 VSS.n11919 9.3
R20328 VSS.n12397 VSS.n12396 9.3
R20329 VSS.n12396 VSS.n12395 9.3
R20330 VSS.n12395 VSS.n12394 9.3
R20331 VSS.n12400 VSS.n12399 9.3
R20332 VSS.n12403 VSS.n12402 9.3
R20333 VSS.n12404 VSS.n12403 9.3
R20334 VSS.n12405 VSS.n12404 9.3
R20335 VSS.n11906 VSS.n11905 9.3
R20336 VSS.n11897 VSS.n11896 9.3
R20337 VSS.n11897 VSS.n11550 9.3
R20338 VSS.n11901 VSS.n11550 9.3
R20339 VSS.n11895 VSS.n11894 9.3
R20340 VSS.n11892 VSS.n11556 9.3
R20341 VSS.n11892 VSS.n11891 9.3
R20342 VSS.n11891 VSS.n11890 9.3
R20343 VSS.n11885 VSS.n11884 9.3
R20344 VSS.n11882 VSS.n11881 9.3
R20345 VSS.n11881 VSS.n11559 9.3
R20346 VSS.n11559 VSS.n11558 9.3
R20347 VSS.n11567 VSS.n11561 9.3
R20348 VSS.n11874 VSS.n11873 9.3
R20349 VSS.n11875 VSS.n11874 9.3
R20350 VSS.n11876 VSS.n11875 9.3
R20351 VSS.n11871 VSS.n11870 9.3
R20352 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector VSS.n11862 9.3
R20353 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector VSS.n11571 9.3
R20354 VSS.n11866 VSS.n11571 9.3
R20355 VSS.n11861 VSS.n11860 9.3
R20356 VSS.n11858 VSS.n11577 9.3
R20357 VSS.n11858 VSS.n11857 9.3
R20358 VSS.n11857 VSS.n11856 9.3
R20359 VSS.n11851 VSS.n11850 9.3
R20360 VSS.n11848 VSS.n11847 9.3
R20361 VSS.n11847 VSS.n11580 9.3
R20362 VSS.n11580 VSS.n11579 9.3
R20363 VSS.n11588 VSS.n11582 9.3
R20364 VSS.n11840 VSS.n11839 9.3
R20365 VSS.n11841 VSS.n11840 9.3
R20366 VSS.n11842 VSS.n11841 9.3
R20367 VSS.n11837 VSS.n11836 9.3
R20368 VSS.n11828 VSS.n11827 9.3
R20369 VSS.n11828 VSS.n11592 9.3
R20370 VSS.n11832 VSS.n11592 9.3
R20371 VSS.n11826 VSS.n11825 9.3
R20372 VSS.n11823 VSS.n11598 9.3
R20373 VSS.n11823 VSS.n11822 9.3
R20374 VSS.n11822 VSS.n11821 9.3
R20375 VSS.n11816 VSS.n11815 9.3
R20376 VSS.n11813 VSS.n11812 9.3
R20377 VSS.n11812 VSS.n11601 9.3
R20378 VSS.n11601 VSS.n11600 9.3
R20379 VSS.n11774 VSS.n11773 9.3
R20380 VSS.n11771 VSS.n11770 9.3
R20381 VSS.n11770 VSS.n11769 9.3
R20382 VSS.n11769 VSS.n11606 9.3
R20383 VSS.n11618 VSS.n11611 9.3
R20384 VSS.n11763 VSS.n11762 9.3
R20385 VSS.n11764 VSS.n11763 9.3
R20386 VSS.n11765 VSS.n11764 9.3
R20387 VSS.n11760 VSS.n11759 9.3
R20388 VSS.n11751 VSS.n11750 9.3
R20389 VSS.n11751 VSS.n11622 9.3
R20390 VSS.n11755 VSS.n11622 9.3
R20391 VSS.n11749 VSS.n11748 9.3
R20392 VSS.n11746 VSS.n11628 9.3
R20393 VSS.n11746 VSS.n11745 9.3
R20394 VSS.n11745 VSS.n11744 9.3
R20395 VSS.n11739 VSS.n11738 9.3
R20396 VSS.n11736 VSS.n11735 9.3
R20397 VSS.n11735 VSS.n11631 9.3
R20398 VSS.n11631 VSS.n11630 9.3
R20399 VSS.n11639 VSS.n11633 9.3
R20400 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector VSS.n11728 9.3
R20401 VSS.n11729 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector 9.3
R20402 VSS.n11730 VSS.n11729 9.3
R20403 VSS.n11726 VSS.n11725 9.3
R20404 VSS.n11717 VSS.n11716 9.3
R20405 VSS.n11717 VSS.n11643 9.3
R20406 VSS.n11721 VSS.n11643 9.3
R20407 VSS.n11715 VSS.n11714 9.3
R20408 VSS.n11712 VSS.n11649 9.3
R20409 VSS.n11712 VSS.n11711 9.3
R20410 VSS.n11711 VSS.n11710 9.3
R20411 VSS.n11705 VSS.n11704 9.3
R20412 VSS.n11702 VSS.n11701 9.3
R20413 VSS.n11701 VSS.n11652 9.3
R20414 VSS.n11652 VSS.n11651 9.3
R20415 VSS.n11660 VSS.n11654 9.3
R20416 VSS.n11694 VSS.n11693 9.3
R20417 VSS.n11695 VSS.n11694 9.3
R20418 VSS.n11696 VSS.n11695 9.3
R20419 VSS.n11691 VSS.n11690 9.3
R20420 VSS.n11682 VSS.n11681 9.3
R20421 VSS.n11682 VSS.n11664 9.3
R20422 VSS.n11686 VSS.n11664 9.3
R20423 VSS.n11680 VSS.n11679 9.3
R20424 VSS.n11677 VSS.n11670 9.3
R20425 VSS.n11677 VSS.n11676 9.3
R20426 VSS.n11676 VSS.n11675 9.3
R20427 VSS.n13400 VSS.n13399 9.3
R20428 VSS.n13403 VSS.n13402 9.3
R20429 VSS.n13403 VSS.n11475 9.3
R20430 VSS.n11475 VSS.n11474 9.3
R20431 VSS.n11479 VSS.n11478 9.3
R20432 VSS.n13411 VSS.n13410 9.3
R20433 VSS.n13410 VSS.n13409 9.3
R20434 VSS.n13409 VSS.n13408 9.3
R20435 VSS.n13412 VSS.n11466 9.3
R20436 VSS.n13415 VSS.n11461 9.3
R20437 VSS.n13416 VSS.n13415 9.3
R20438 VSS.n13417 VSS.n13416 9.3
R20439 VSS.n13423 VSS.n13422 9.3
R20440 VSS.n13426 VSS.n13425 9.3
R20441 VSS.n13426 VSS.n11456 9.3
R20442 VSS.n11456 VSS.n11455 9.3
R20443 VSS.n11460 VSS.n11459 9.3
R20444 VSS.n13434 VSS.n13433 9.3
R20445 VSS.n13433 VSS.n13432 9.3
R20446 VSS.n13432 VSS.n13431 9.3
R20447 VSS.n13435 VSS.n11447 9.3
R20448 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector VSS.n11442 9.3
R20449 VSS.n13438 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector 9.3
R20450 VSS.n13439 VSS.n13438 9.3
R20451 VSS.n13445 VSS.n13444 9.3
R20452 VSS.n13448 VSS.n13447 9.3
R20453 VSS.n13448 VSS.n11437 9.3
R20454 VSS.n11437 VSS.n11436 9.3
R20455 VSS.n11441 VSS.n11440 9.3
R20456 VSS.n13456 VSS.n13455 9.3
R20457 VSS.n13455 VSS.n13454 9.3
R20458 VSS.n13454 VSS.n13453 9.3
R20459 VSS.n13272 VSS.n11429 9.3
R20460 VSS.n13278 VSS.n13277 9.3
R20461 VSS.n13278 VSS.n13267 9.3
R20462 VSS.n13267 VSS.n13266 9.3
R20463 VSS.n13275 VSS.n13274 9.3
R20464 VSS.n13286 VSS.n13285 9.3
R20465 VSS.n13285 VSS.n13284 9.3
R20466 VSS.n13284 VSS.n13283 9.3
R20467 VSS.n13287 VSS.n13258 9.3
R20468 VSS.n13290 VSS.n13252 9.3
R20469 VSS.n13291 VSS.n13290 9.3
R20470 VSS.n13292 VSS.n13291 9.3
R20471 VSS.n13298 VSS.n13297 9.3
R20472 VSS.n13301 VSS.n13300 9.3
R20473 VSS.n13301 VSS.n13250 9.3
R20474 VSS.n13255 VSS.n13250 9.3
R20475 VSS.n13313 VSS.n13312 9.3
R20476 VSS.n13310 VSS.n13309 9.3
R20477 VSS.n13309 VSS.n13308 9.3
R20478 VSS.n13308 VSS.n13307 9.3
R20479 VSS.n13244 VSS.n12520 9.3
R20480 VSS.n13241 VSS.n12526 9.3
R20481 VSS.n12526 VSS.n12525 9.3
R20482 VSS.n12525 VSS.n12524 9.3
R20483 VSS.n13240 VSS.n13239 9.3
R20484 VSS.n13230 VSS.n13229 9.3
R20485 VSS.n13230 VSS.n12530 9.3
R20486 VSS.n13234 VSS.n12530 9.3
R20487 VSS.n13228 VSS.n13227 9.3
R20488 VSS.n13225 VSS.n12537 9.3
R20489 VSS.n13225 VSS.n13224 9.3
R20490 VSS.n13224 VSS.n13223 9.3
R20491 VSS.n13218 VSS.n13217 9.3
R20492 VSS.n13215 VSS.n13214 9.3
R20493 VSS.n13214 VSS.n12540 9.3
R20494 VSS.n12540 VSS.n12539 9.3
R20495 VSS.n12548 VSS.n12542 9.3
R20496 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector VSS.n13207 9.3
R20497 VSS.n13208 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector 9.3
R20498 VSS.n13209 VSS.n13208 9.3
R20499 VSS.n13205 VSS.n13204 9.3
R20500 VSS.n13196 VSS.n13195 9.3
R20501 VSS.n13196 VSS.n12552 9.3
R20502 VSS.n13200 VSS.n12552 9.3
R20503 VSS.n13194 VSS.n13193 9.3
R20504 VSS.n13191 VSS.n12558 9.3
R20505 VSS.n13191 VSS.n13190 9.3
R20506 VSS.n13190 VSS.n13189 9.3
R20507 VSS.n13184 VSS.n13183 9.3
R20508 VSS.n13181 VSS.n13180 9.3
R20509 VSS.n13180 VSS.n12561 9.3
R20510 VSS.n12561 VSS.n12560 9.3
R20511 VSS.n12569 VSS.n12563 9.3
R20512 VSS.n13173 VSS.n13172 9.3
R20513 VSS.n13174 VSS.n13173 9.3
R20514 VSS.n13175 VSS.n13174 9.3
R20515 VSS.n13170 VSS.n13169 9.3
R20516 VSS.n13161 VSS.n13160 9.3
R20517 VSS.n13161 VSS.n12573 9.3
R20518 VSS.n13165 VSS.n12573 9.3
R20519 VSS.n13159 VSS.n13158 9.3
R20520 VSS.n13156 VSS.n12579 9.3
R20521 VSS.n13156 VSS.n13155 9.3
R20522 VSS.n13155 VSS.n13154 9.3
R20523 VSS.n12959 VSS.n12583 9.3
R20524 VSS.n12969 VSS.n12968 9.3
R20525 VSS.n12968 VSS.n12967 9.3
R20526 VSS.n12967 VSS.n12966 9.3
R20527 VSS.n12970 VSS.n12958 9.3
R20528 VSS.n12973 VSS.n12953 9.3
R20529 VSS.n12974 VSS.n12973 9.3
R20530 VSS.n12975 VSS.n12974 9.3
R20531 VSS.n12981 VSS.n12980 9.3
R20532 VSS.n12984 VSS.n12983 9.3
R20533 VSS.n12984 VSS.n12948 9.3
R20534 VSS.n12948 VSS.n12947 9.3
R20535 VSS.n12952 VSS.n12951 9.3
R20536 VSS.n12992 VSS.n12991 9.3
R20537 VSS.n12991 VSS.n12990 9.3
R20538 VSS.n12990 VSS.n12989 9.3
R20539 VSS.n12993 VSS.n12939 9.3
R20540 VSS.n12996 VSS.n12934 9.3
R20541 VSS.n12997 VSS.n12996 9.3
R20542 VSS.n12998 VSS.n12997 9.3
R20543 VSS.n13004 VSS.n13003 9.3
R20544 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector VSS.n13006 9.3
R20545 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector VSS.n12929 9.3
R20546 VSS.n12929 VSS.n12928 9.3
R20547 VSS.n12933 VSS.n12932 9.3
R20548 VSS.n13014 VSS.n13013 9.3
R20549 VSS.n13013 VSS.n13012 9.3
R20550 VSS.n13012 VSS.n13011 9.3
R20551 VSS.n13015 VSS.n12920 9.3
R20552 VSS.n13018 VSS.n12915 9.3
R20553 VSS.n13019 VSS.n13018 9.3
R20554 VSS.n13020 VSS.n13019 9.3
R20555 VSS.n13026 VSS.n13025 9.3
R20556 VSS.n13029 VSS.n13028 9.3
R20557 VSS.n13029 VSS.n12910 9.3
R20558 VSS.n12910 VSS.n12909 9.3
R20559 VSS.n12914 VSS.n12913 9.3
R20560 VSS.n13037 VSS.n13036 9.3
R20561 VSS.n13036 VSS.n13035 9.3
R20562 VSS.n13035 VSS.n13034 9.3
R20563 VSS.n13038 VSS.n12901 9.3
R20564 VSS.n13041 VSS.n12895 9.3
R20565 VSS.n13042 VSS.n13041 9.3
R20566 VSS.n13043 VSS.n13042 9.3
R20567 VSS.n13049 VSS.n13048 9.3
R20568 VSS.n13052 VSS.n13051 9.3
R20569 VSS.n13052 VSS.n12893 9.3
R20570 VSS.n12898 VSS.n12893 9.3
R20571 VSS.n13064 VSS.n13063 9.3
R20572 VSS.n13061 VSS.n13060 9.3
R20573 VSS.n13060 VSS.n13059 9.3
R20574 VSS.n13059 VSS.n13058 9.3
R20575 VSS.n12887 VSS.n12661 9.3
R20576 VSS.n12884 VSS.n12667 9.3
R20577 VSS.n12667 VSS.n12666 9.3
R20578 VSS.n12666 VSS.n12665 9.3
R20579 VSS.n12883 VSS.n12882 9.3
R20580 VSS.n12873 VSS.n12872 9.3
R20581 VSS.n12873 VSS.n12671 9.3
R20582 VSS.n12877 VSS.n12671 9.3
R20583 VSS.n12871 VSS.n12870 9.3
R20584 VSS.n12868 VSS.n12678 9.3
R20585 VSS.n12868 VSS.n12867 9.3
R20586 VSS.n12867 VSS.n12866 9.3
R20587 VSS.n12861 VSS.n12860 9.3
R20588 VSS.n12858 VSS.n12857 9.3
R20589 VSS.n12857 VSS.n12681 9.3
R20590 VSS.n12681 VSS.n12680 9.3
R20591 VSS.n12689 VSS.n12683 9.3
R20592 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Collector VSS.n12850 9.3
R20593 VSS.n12851 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Collector 9.3
R20594 VSS.n12852 VSS.n12851 9.3
R20595 VSS.n12848 VSS.n12847 9.3
R20596 VSS.n12839 VSS.n12838 9.3
R20597 VSS.n12839 VSS.n12693 9.3
R20598 VSS.n12843 VSS.n12693 9.3
R20599 VSS.n12837 VSS.n12836 9.3
R20600 VSS.n12834 VSS.n12699 9.3
R20601 VSS.n12834 VSS.n12833 9.3
R20602 VSS.n12833 VSS.n12832 9.3
R20603 VSS.n12827 VSS.n12826 9.3
R20604 VSS.n12824 VSS.n12823 9.3
R20605 VSS.n12823 VSS.n12702 9.3
R20606 VSS.n12702 VSS.n12701 9.3
R20607 VSS.n12710 VSS.n12704 9.3
R20608 VSS.n12816 VSS.n12815 9.3
R20609 VSS.n12817 VSS.n12816 9.3
R20610 VSS.n12818 VSS.n12817 9.3
R20611 VSS.n12813 VSS.n12812 9.3
R20612 VSS.n12804 VSS.n12803 9.3
R20613 VSS.n12804 VSS.n12714 9.3
R20614 VSS.n12808 VSS.n12714 9.3
R20615 VSS.n12802 VSS.n12801 9.3
R20616 VSS.n12799 VSS.n12720 9.3
R20617 VSS.n12799 VSS.n12798 9.3
R20618 VSS.n12798 VSS.n12797 9.3
R20619 VSS.n12218 VSS.n12057 9.3
R20620 VSS.n12219 VSS.n12218 9.3
R20621 VSS.n12220 VSS.n12219 9.3
R20622 VSS.n12215 VSS.n12062 9.3
R20623 VSS.n13921 VSS.n13920 9.3
R20624 VSS.n13920 VSS.n13919 9.3
R20625 VSS.n13923 VSS.n13922 9.3
R20626 VSS.n13927 VSS.n13926 9.3
R20627 VSS.n13926 VSS.n13925 9.3
R20628 VSS.n13933 VSS.n13932 9.3
R20629 VSS.n13932 VSS.n13931 9.3
R20630 VSS.n13934 VSS.n13900 9.3
R20631 VSS.n13938 VSS.n13899 9.3
R20632 VSS.n13938 VSS.n13937 9.3
R20633 VSS.n13947 VSS.n13945 9.3
R20634 VSS.n13947 VSS.n13946 9.3
R20635 VSS.n13898 VSS.n10515 9.3
R20636 VSS.n13895 VSS.n10517 9.3
R20637 VSS.n13895 VSS.n10514 9.3
R20638 VSS.n13888 VSS.n13887 9.3
R20639 VSS.n13887 VSS.n13886 9.3
R20640 VSS.n13891 VSS.n13890 9.3
R20641 VSS.n13929 VSS.n13928 9.3
R20642 VSS.n13943 VSS.n13942 9.3
R20643 VSS.n13917 VSS.n13916 9.3
R20644 VSS.n13829 VSS.n10498 9.3
R20645 VSS.n13953 VSS.n10498 9.3
R20646 VSS.n13953 VSS.n13952 9.3
R20647 VSS.n13832 VSS.n13828 9.3
R20648 VSS.n13754 VSS.n13753 9.3
R20649 VSS.n13753 VSS.n10522 9.3
R20650 VSS.n13802 VSS.n10522 9.3
R20651 VSS.n13765 VSS.n13764 9.3
R20652 VSS.n13764 VSS.n10547 9.3
R20653 VSS.n13767 VSS.n13766 9.3
R20654 VSS.n13771 VSS.n13770 9.3
R20655 VSS.n13770 VSS.n13769 9.3
R20656 VSS.n13777 VSS.n13776 9.3
R20657 VSS.n13776 VSS.n13775 9.3
R20658 VSS.n13779 VSS.n13778 9.3
R20659 VSS.n13783 VSS.n13782 9.3
R20660 VSS.n13782 VSS.n13781 9.3
R20661 VSS.n13788 VSS.n13727 9.3
R20662 VSS.n13788 VSS.n13787 9.3
R20663 VSS.n13793 VSS.n13792 9.3
R20664 VSS.n13797 VSS.n13795 9.3
R20665 VSS.n13797 VSS.n13796 9.3
R20666 VSS.n13723 VSS.n10560 9.3
R20667 VSS.n13723 VSS.n10557 9.3
R20668 VSS.n13726 VSS.n10558 9.3
R20669 VSS.n13762 VSS.n13761 9.3
R20670 VSS.n13773 VSS.n13772 9.3
R20671 VSS.n13784 VSS.n13728 9.3
R20672 VSS.n13664 VSS.n13663 9.3
R20673 VSS.n13663 VSS.n10612 9.3
R20674 VSS.n13712 VSS.n10612 9.3
R20675 VSS.n13675 VSS.n13674 9.3
R20676 VSS.n13674 VSS.n10637 9.3
R20677 VSS.n13677 VSS.n13676 9.3
R20678 VSS.n13681 VSS.n13680 9.3
R20679 VSS.n13680 VSS.n13679 9.3
R20680 VSS.n13687 VSS.n13686 9.3
R20681 VSS.n13686 VSS.n13685 9.3
R20682 VSS.n13689 VSS.n13688 9.3
R20683 VSS.n13693 VSS.n13692 9.3
R20684 VSS.n13692 VSS.n13691 9.3
R20685 VSS.n13698 VSS.n13637 9.3
R20686 VSS.n13698 VSS.n13697 9.3
R20687 VSS.n13703 VSS.n13702 9.3
R20688 VSS.n13707 VSS.n13705 9.3
R20689 VSS.n13707 VSS.n13706 9.3
R20690 VSS.n13633 VSS.n10650 9.3
R20691 VSS.n13633 VSS.n10647 9.3
R20692 VSS.n13636 VSS.n10648 9.3
R20693 VSS.n13672 VSS.n13671 9.3
R20694 VSS.n13683 VSS.n13682 9.3
R20695 VSS.n13694 VSS.n13638 9.3
R20696 VSS.n13574 VSS.n13573 9.3
R20697 VSS.n13573 VSS.n10702 9.3
R20698 VSS.n13622 VSS.n10702 9.3
R20699 VSS.n13585 VSS.n13584 9.3
R20700 VSS.n13584 VSS.n10727 9.3
R20701 VSS.n13587 VSS.n13586 9.3
R20702 VSS.n13591 VSS.n13590 9.3
R20703 VSS.n13590 VSS.n13589 9.3
R20704 VSS.n13597 VSS.n13596 9.3
R20705 VSS.n13596 VSS.n13595 9.3
R20706 VSS.n13599 VSS.n13598 9.3
R20707 VSS.n13603 VSS.n13602 9.3
R20708 VSS.n13602 VSS.n13601 9.3
R20709 VSS.n13608 VSS.n13547 9.3
R20710 VSS.n13608 VSS.n13607 9.3
R20711 VSS.n13613 VSS.n13612 9.3
R20712 VSS.n13617 VSS.n13615 9.3
R20713 VSS.n13617 VSS.n13616 9.3
R20714 VSS.n13543 VSS.n10740 9.3
R20715 VSS.n13543 VSS.n10737 9.3
R20716 VSS.n13546 VSS.n10738 9.3
R20717 VSS.n13582 VSS.n13581 9.3
R20718 VSS.n13593 VSS.n13592 9.3
R20719 VSS.n13604 VSS.n13548 9.3
R20720 VSS.n13483 VSS.n13482 9.3
R20721 VSS.n13482 VSS.n10792 9.3
R20722 VSS.n13532 VSS.n10792 9.3
R20723 VSS.n13494 VSS.n13493 9.3
R20724 VSS.n13493 VSS.n10817 9.3
R20725 VSS.n13496 VSS.n13495 9.3
R20726 VSS.n13500 VSS.n13499 9.3
R20727 VSS.n13499 VSS.n13498 9.3
R20728 VSS.n13506 VSS.n13505 9.3
R20729 VSS.n13505 VSS.n13504 9.3
R20730 VSS.n13508 VSS.n13507 9.3
R20731 VSS.n13512 VSS.n13511 9.3
R20732 VSS.n13511 VSS.n13510 9.3
R20733 VSS.n13518 VSS.n11427 9.3
R20734 VSS.n13518 VSS.n13517 9.3
R20735 VSS.n13523 VSS.n13522 9.3
R20736 VSS.n13527 VSS.n13525 9.3
R20737 VSS.n13527 VSS.n13526 9.3
R20738 VSS.n11423 VSS.n10830 9.3
R20739 VSS.n11423 VSS.n10827 9.3
R20740 VSS.n11426 VSS.n10828 9.3
R20741 VSS.n13491 VSS.n13490 9.3
R20742 VSS.n13502 VSS.n13501 9.3
R20743 VSS.n13514 VSS.n11428 9.3
R20744 VSS.n11364 VSS.n11363 9.3
R20745 VSS.n11363 VSS.n10882 9.3
R20746 VSS.n11412 VSS.n10882 9.3
R20747 VSS.n11375 VSS.n11374 9.3
R20748 VSS.n11374 VSS.n10907 9.3
R20749 VSS.n11377 VSS.n11376 9.3
R20750 VSS.n11381 VSS.n11380 9.3
R20751 VSS.n11380 VSS.n11379 9.3
R20752 VSS.n11387 VSS.n11386 9.3
R20753 VSS.n11386 VSS.n11385 9.3
R20754 VSS.n11389 VSS.n11388 9.3
R20755 VSS.n11393 VSS.n11392 9.3
R20756 VSS.n11392 VSS.n11391 9.3
R20757 VSS.n11398 VSS.n11337 9.3
R20758 VSS.n11398 VSS.n11397 9.3
R20759 VSS.n11403 VSS.n11402 9.3
R20760 VSS.n11407 VSS.n11405 9.3
R20761 VSS.n11407 VSS.n11406 9.3
R20762 VSS.n11333 VSS.n10920 9.3
R20763 VSS.n11333 VSS.n10917 9.3
R20764 VSS.n11336 VSS.n10918 9.3
R20765 VSS.n11372 VSS.n11371 9.3
R20766 VSS.n11383 VSS.n11382 9.3
R20767 VSS.n11394 VSS.n11338 9.3
R20768 VSS.n11274 VSS.n11273 9.3
R20769 VSS.n11273 VSS.n10972 9.3
R20770 VSS.n11322 VSS.n10972 9.3
R20771 VSS.n11285 VSS.n11284 9.3
R20772 VSS.n11284 VSS.n10997 9.3
R20773 VSS.n11287 VSS.n11286 9.3
R20774 VSS.n11291 VSS.n11290 9.3
R20775 VSS.n11290 VSS.n11289 9.3
R20776 VSS.n11297 VSS.n11296 9.3
R20777 VSS.n11296 VSS.n11295 9.3
R20778 VSS.n11299 VSS.n11298 9.3
R20779 VSS.n11303 VSS.n11302 9.3
R20780 VSS.n11302 VSS.n11301 9.3
R20781 VSS.n11308 VSS.n11247 9.3
R20782 VSS.n11308 VSS.n11307 9.3
R20783 VSS.n11313 VSS.n11312 9.3
R20784 VSS.n11317 VSS.n11315 9.3
R20785 VSS.n11317 VSS.n11316 9.3
R20786 VSS.n11243 VSS.n11010 9.3
R20787 VSS.n11243 VSS.n11007 9.3
R20788 VSS.n11246 VSS.n11008 9.3
R20789 VSS.n11282 VSS.n11281 9.3
R20790 VSS.n11293 VSS.n11292 9.3
R20791 VSS.n11304 VSS.n11248 9.3
R20792 VSS.n11184 VSS.n11183 9.3
R20793 VSS.n11183 VSS.n11062 9.3
R20794 VSS.n11232 VSS.n11062 9.3
R20795 VSS.n11195 VSS.n11194 9.3
R20796 VSS.n11194 VSS.n11087 9.3
R20797 VSS.n11197 VSS.n11196 9.3
R20798 VSS.n11201 VSS.n11200 9.3
R20799 VSS.n11200 VSS.n11199 9.3
R20800 VSS.n11207 VSS.n11206 9.3
R20801 VSS.n11206 VSS.n11205 9.3
R20802 VSS.n11209 VSS.n11208 9.3
R20803 VSS.n11213 VSS.n11212 9.3
R20804 VSS.n11212 VSS.n11211 9.3
R20805 VSS.n11218 VSS.n11157 9.3
R20806 VSS.n11218 VSS.n11217 9.3
R20807 VSS.n11223 VSS.n11222 9.3
R20808 VSS.n11227 VSS.n11225 9.3
R20809 VSS.n11227 VSS.n11226 9.3
R20810 VSS.n11153 VSS.n11100 9.3
R20811 VSS.n11153 VSS.n11097 9.3
R20812 VSS.n11156 VSS.n11098 9.3
R20813 VSS.n11192 VSS.n11191 9.3
R20814 VSS.n11203 VSS.n11202 9.3
R20815 VSS.n11214 VSS.n11158 9.3
R20816 VSS.n11190 VSS.n11189 9.3
R20817 VSS.n11189 VSS.n11188 9.3
R20818 VSS.n11186 VSS.n11185 9.3
R20819 VSS.n11060 VSS.n11059 9.3
R20820 VSS.n11280 VSS.n11279 9.3
R20821 VSS.n11279 VSS.n11278 9.3
R20822 VSS.n11276 VSS.n11275 9.3
R20823 VSS.n10970 VSS.n10969 9.3
R20824 VSS.n11370 VSS.n11369 9.3
R20825 VSS.n11369 VSS.n11368 9.3
R20826 VSS.n11366 VSS.n11365 9.3
R20827 VSS.n10880 VSS.n10879 9.3
R20828 VSS.n13489 VSS.n13488 9.3
R20829 VSS.n13488 VSS.n13487 9.3
R20830 VSS.n13485 VSS.n13484 9.3
R20831 VSS.n10790 VSS.n10789 9.3
R20832 VSS.n13580 VSS.n13579 9.3
R20833 VSS.n13579 VSS.n13578 9.3
R20834 VSS.n13576 VSS.n13575 9.3
R20835 VSS.n10700 VSS.n10699 9.3
R20836 VSS.n13670 VSS.n13669 9.3
R20837 VSS.n13669 VSS.n13668 9.3
R20838 VSS.n13666 VSS.n13665 9.3
R20839 VSS.n10610 VSS.n10609 9.3
R20840 VSS.n13760 VSS.n13759 9.3
R20841 VSS.n13759 VSS.n13758 9.3
R20842 VSS.n13756 VSS.n13755 9.3
R20843 VSS.n10520 VSS.n10519 9.3
R20844 VSS.n10493 VSS.n10491 9.3
R20845 VSS.n10499 VSS.n10493 9.3
R20846 VSS.n13957 VSS.n10492 9.3
R20847 VSS.n10483 VSS.n10419 9.3
R20848 VSS.n10478 VSS.n10421 9.3
R20849 VSS.n10473 VSS.n10423 9.3
R20850 VSS.n10468 VSS.n10425 9.3
R20851 VSS.n10443 VSS.n10442 9.3
R20852 VSS.n10448 VSS.n10441 9.3
R20853 VSS.n10453 VSS.n10440 9.3
R20854 VSS.n10458 VSS.n10439 9.3
R20855 VSS.n10460 VSS.n10459 9.3
R20856 VSS.n10457 VSS.n10456 9.3
R20857 VSS.n10455 VSS.n10454 9.3
R20858 VSS.n10452 VSS.n10451 9.3
R20859 VSS.n10450 VSS.n10449 9.3
R20860 VSS.n10447 VSS.n10446 9.3
R20861 VSS.n10445 VSS.n10444 9.3
R20862 VSS.n10428 VSS.n10427 9.3
R20863 VSS.n10467 VSS.n10466 9.3
R20864 VSS.n10470 VSS.n10469 9.3
R20865 VSS.n10472 VSS.n10471 9.3
R20866 VSS.n10475 VSS.n10474 9.3
R20867 VSS.n10477 VSS.n10476 9.3
R20868 VSS.n10480 VSS.n10479 9.3
R20869 VSS.n10482 VSS.n10481 9.3
R20870 VSS.n10485 VSS.n10484 9.3
R20871 VSS.n7162 VSS.n7161 9.3
R20872 VSS.n7161 VSS.n7012 9.3
R20873 VSS.n7012 VSS.n7011 9.3
R20874 VSS.n7020 VSS.n7014 9.3
R20875 VSS.n7154 VSS.n7153 9.3
R20876 VSS.n7155 VSS.n7154 9.3
R20877 VSS.n7156 VSS.n7155 9.3
R20878 VSS.n7142 VSS.n7141 9.3
R20879 VSS.n7142 VSS.n7024 9.3
R20880 VSS.n7146 VSS.n7024 9.3
R20881 VSS.n7140 VSS.n7139 9.3
R20882 VSS.n7137 VSS.n7030 9.3
R20883 VSS.n7137 VSS.n7136 9.3
R20884 VSS.n7136 VSS.n7135 9.3
R20885 VSS.n7127 sky130_asc_pnp_05v5_W3p40L3p40_8_1/xm1/Collector 9.3
R20886 sky130_asc_pnp_05v5_W3p40L3p40_8_1/xm1/Collector VSS.n7033 9.3
R20887 VSS.n7033 VSS.n7032 9.3
R20888 VSS.n7041 VSS.n7035 9.3
R20889 VSS.n7120 VSS.n7119 9.3
R20890 VSS.n7121 VSS.n7120 9.3
R20891 VSS.n7122 VSS.n7121 9.3
R20892 VSS.n7108 VSS.n7107 9.3
R20893 VSS.n7108 VSS.n7045 9.3
R20894 VSS.n7112 VSS.n7045 9.3
R20895 VSS.n7106 VSS.n7105 9.3
R20896 VSS.n7103 VSS.n7051 9.3
R20897 VSS.n7103 VSS.n7102 9.3
R20898 VSS.n7102 VSS.n7101 9.3
R20899 VSS.n7093 VSS.n7092 9.3
R20900 VSS.n7092 VSS.n7054 9.3
R20901 VSS.n7054 VSS.n7053 9.3
R20902 VSS.n7062 VSS.n7056 9.3
R20903 VSS.n7085 VSS.n7084 9.3
R20904 VSS.n7086 VSS.n7085 9.3
R20905 VSS.n7087 VSS.n7086 9.3
R20906 VSS.n7073 VSS.n7072 9.3
R20907 VSS.n7073 VSS.n7066 9.3
R20908 VSS.n7077 VSS.n7066 9.3
R20909 VSS.n7165 VSS.n7164 9.3
R20910 VSS.n7151 VSS.n7150 9.3
R20911 VSS.n7130 VSS.n7129 9.3
R20912 VSS.n7117 VSS.n7116 9.3
R20913 VSS.n7096 VSS.n7095 9.3
R20914 VSS.n7082 VSS.n7081 9.3
R20915 VSS.n7070 VSS.n7069 9.3
R20916 VSS.n8860 VSS.n8859 9.3
R20917 VSS.n8859 VSS.n8858 9.3
R20918 VSS.n8858 VSS.n8857 9.3
R20919 VSS.n8861 VSS.n6957 9.3
R20920 VSS.n8864 VSS.n6952 9.3
R20921 VSS.n8865 VSS.n8864 9.3
R20922 VSS.n8866 VSS.n8865 9.3
R20923 VSS.n8872 VSS.n8871 9.3
R20924 VSS.n8875 VSS.n8874 9.3
R20925 VSS.n8875 VSS.n6947 9.3
R20926 VSS.n6947 VSS.n6946 9.3
R20927 VSS.n6951 VSS.n6950 9.3
R20928 VSS.n8883 VSS.n8882 9.3
R20929 VSS.n8882 VSS.n8881 9.3
R20930 VSS.n8881 VSS.n8880 9.3
R20931 VSS.n8884 VSS.n6938 9.3
R20932 VSS.n8887 VSS.n6933 9.3
R20933 VSS.n8888 VSS.n8887 9.3
R20934 VSS.n8889 VSS.n8888 9.3
R20935 VSS.n8895 VSS.n8894 9.3
R20936 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector VSS.n8897 9.3
R20937 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector VSS.n6928 9.3
R20938 VSS.n6928 VSS.n6927 9.3
R20939 VSS.n6932 VSS.n6931 9.3
R20940 VSS.n8905 VSS.n8904 9.3
R20941 VSS.n8904 VSS.n8903 9.3
R20942 VSS.n8903 VSS.n8902 9.3
R20943 VSS.n8906 VSS.n6919 9.3
R20944 VSS.n8909 VSS.n6914 9.3
R20945 VSS.n8910 VSS.n8909 9.3
R20946 VSS.n8911 VSS.n8910 9.3
R20947 VSS.n8917 VSS.n8916 9.3
R20948 VSS.n8920 VSS.n8919 9.3
R20949 VSS.n8920 VSS.n6909 9.3
R20950 VSS.n6909 VSS.n6908 9.3
R20951 VSS.n6913 VSS.n6912 9.3
R20952 VSS.n8928 VSS.n8927 9.3
R20953 VSS.n8927 VSS.n8926 9.3
R20954 VSS.n8926 VSS.n8925 9.3
R20955 VSS.n8748 VSS.n6901 9.3
R20956 VSS.n8754 VSS.n8747 9.3
R20957 VSS.n8754 VSS.n8753 9.3
R20958 VSS.n8753 VSS.n8752 9.3
R20959 VSS.n8745 VSS.n8739 9.3
R20960 VSS.n8742 VSS.n8741 9.3
R20961 VSS.n8742 VSS.n8736 9.3
R20962 VSS.n8759 VSS.n8736 9.3
R20963 VSS.n8766 VSS.n8765 9.3
R20964 VSS.n8769 VSS.n8768 9.3
R20965 VSS.n8770 VSS.n8769 9.3
R20966 VSS.n8771 VSS.n8770 9.3
R20967 VSS.n8733 VSS.n8732 9.3
R20968 VSS.n8724 VSS.n8723 9.3
R20969 VSS.n8724 VSS.n7264 9.3
R20970 VSS.n8728 VSS.n7264 9.3
R20971 VSS.n8722 VSS.n8721 9.3
R20972 VSS.n8719 VSS.n7270 9.3
R20973 VSS.n8719 VSS.n8718 9.3
R20974 VSS.n8718 VSS.n8717 9.3
R20975 VSS.n8712 VSS.n8711 9.3
R20976 VSS.n8709 VSS.n8708 9.3
R20977 VSS.n8708 VSS.n7273 9.3
R20978 VSS.n7273 VSS.n7272 9.3
R20979 VSS.n7281 VSS.n7275 9.3
R20980 VSS.n8701 VSS.n8700 9.3
R20981 VSS.n8702 VSS.n8701 9.3
R20982 VSS.n8703 VSS.n8702 9.3
R20983 VSS.n8698 VSS.n8697 9.3
R20984 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector VSS.n8689 9.3
R20985 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector VSS.n7285 9.3
R20986 VSS.n8693 VSS.n7285 9.3
R20987 VSS.n8688 VSS.n8687 9.3
R20988 VSS.n8685 VSS.n7291 9.3
R20989 VSS.n8685 VSS.n8684 9.3
R20990 VSS.n8684 VSS.n8683 9.3
R20991 VSS.n8678 VSS.n8677 9.3
R20992 VSS.n8675 VSS.n8674 9.3
R20993 VSS.n8674 VSS.n7294 9.3
R20994 VSS.n7294 VSS.n7293 9.3
R20995 VSS.n7302 VSS.n7296 9.3
R20996 VSS.n8667 VSS.n8666 9.3
R20997 VSS.n8668 VSS.n8667 9.3
R20998 VSS.n8669 VSS.n8668 9.3
R20999 VSS.n8664 VSS.n8663 9.3
R21000 VSS.n8655 VSS.n8654 9.3
R21001 VSS.n8655 VSS.n7306 9.3
R21002 VSS.n8659 VSS.n7306 9.3
R21003 VSS.n8653 VSS.n8652 9.3
R21004 VSS.n8650 VSS.n7312 9.3
R21005 VSS.n8650 VSS.n8649 9.3
R21006 VSS.n8649 VSS.n8648 9.3
R21007 VSS.n8643 VSS.n8642 9.3
R21008 VSS.n8640 VSS.n8639 9.3
R21009 VSS.n8639 VSS.n7315 9.3
R21010 VSS.n7315 VSS.n7314 9.3
R21011 VSS.n8454 VSS.n8453 9.3
R21012 VSS.n8457 VSS.n8456 9.3
R21013 VSS.n8457 VSS.n8448 9.3
R21014 VSS.n8448 VSS.n7320 9.3
R21015 VSS.n8452 VSS.n8451 9.3
R21016 VSS.n8465 VSS.n8464 9.3
R21017 VSS.n8464 VSS.n8463 9.3
R21018 VSS.n8463 VSS.n8462 9.3
R21019 VSS.n8466 VSS.n8440 9.3
R21020 VSS.n8469 VSS.n8435 9.3
R21021 VSS.n8470 VSS.n8469 9.3
R21022 VSS.n8471 VSS.n8470 9.3
R21023 VSS.n8477 VSS.n8476 9.3
R21024 VSS.n8480 VSS.n8479 9.3
R21025 VSS.n8480 VSS.n8430 9.3
R21026 VSS.n8430 VSS.n8429 9.3
R21027 VSS.n8434 VSS.n8433 9.3
R21028 VSS.n8488 VSS.n8487 9.3
R21029 VSS.n8487 VSS.n8486 9.3
R21030 VSS.n8486 VSS.n8485 9.3
R21031 VSS.n8489 VSS.n8421 9.3
R21032 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector VSS.n8416 9.3
R21033 VSS.n8492 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector 9.3
R21034 VSS.n8493 VSS.n8492 9.3
R21035 VSS.n8499 VSS.n8498 9.3
R21036 VSS.n8502 VSS.n8501 9.3
R21037 VSS.n8502 VSS.n8411 9.3
R21038 VSS.n8411 VSS.n8410 9.3
R21039 VSS.n8415 VSS.n8414 9.3
R21040 VSS.n8510 VSS.n8509 9.3
R21041 VSS.n8509 VSS.n8508 9.3
R21042 VSS.n8508 VSS.n8507 9.3
R21043 VSS.n8511 VSS.n8402 9.3
R21044 VSS.n8514 VSS.n8397 9.3
R21045 VSS.n8515 VSS.n8514 9.3
R21046 VSS.n8516 VSS.n8515 9.3
R21047 VSS.n8522 VSS.n8521 9.3
R21048 VSS.n8525 VSS.n8524 9.3
R21049 VSS.n8525 VSS.n8391 9.3
R21050 VSS.n8391 VSS.n8390 9.3
R21051 VSS.n8396 VSS.n8395 9.3
R21052 VSS.n8532 VSS.n8388 9.3
R21053 VSS.n8532 VSS.n8531 9.3
R21054 VSS.n8531 VSS.n8530 9.3
R21055 VSS.n8387 VSS.n8381 9.3
R21056 VSS.n8384 VSS.n8383 9.3
R21057 VSS.n8384 VSS.n8378 9.3
R21058 VSS.n8537 VSS.n8378 9.3
R21059 VSS.n8544 VSS.n8543 9.3
R21060 VSS.n8547 VSS.n8546 9.3
R21061 VSS.n8548 VSS.n8547 9.3
R21062 VSS.n8549 VSS.n8548 9.3
R21063 VSS.n8375 VSS.n8374 9.3
R21064 VSS.n8366 VSS.n8365 9.3
R21065 VSS.n8366 VSS.n7404 9.3
R21066 VSS.n8370 VSS.n7404 9.3
R21067 VSS.n8364 VSS.n8363 9.3
R21068 VSS.n8361 VSS.n7410 9.3
R21069 VSS.n8361 VSS.n8360 9.3
R21070 VSS.n8360 VSS.n8359 9.3
R21071 VSS.n8354 VSS.n8353 9.3
R21072 VSS.n8351 VSS.n8350 9.3
R21073 VSS.n8350 VSS.n7413 9.3
R21074 VSS.n7413 VSS.n7412 9.3
R21075 VSS.n7421 VSS.n7415 9.3
R21076 VSS.n8343 VSS.n8342 9.3
R21077 VSS.n8344 VSS.n8343 9.3
R21078 VSS.n8345 VSS.n8344 9.3
R21079 VSS.n8340 VSS.n8339 9.3
R21080 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector VSS.n8331 9.3
R21081 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector VSS.n7425 9.3
R21082 VSS.n8335 VSS.n7425 9.3
R21083 VSS.n8330 VSS.n8329 9.3
R21084 VSS.n8327 VSS.n7431 9.3
R21085 VSS.n8327 VSS.n8326 9.3
R21086 VSS.n8326 VSS.n8325 9.3
R21087 VSS.n8320 VSS.n8319 9.3
R21088 VSS.n8317 VSS.n8316 9.3
R21089 VSS.n8316 VSS.n7434 9.3
R21090 VSS.n7434 VSS.n7433 9.3
R21091 VSS.n7442 VSS.n7436 9.3
R21092 VSS.n8309 VSS.n8308 9.3
R21093 VSS.n8310 VSS.n8309 9.3
R21094 VSS.n8311 VSS.n8310 9.3
R21095 VSS.n8306 VSS.n8305 9.3
R21096 VSS.n8297 VSS.n8296 9.3
R21097 VSS.n8297 VSS.n7446 9.3
R21098 VSS.n8301 VSS.n7446 9.3
R21099 VSS.n8295 VSS.n8294 9.3
R21100 VSS.n8292 VSS.n7452 9.3
R21101 VSS.n8292 VSS.n8291 9.3
R21102 VSS.n8291 VSS.n8290 9.3
R21103 VSS.n8285 VSS.n8284 9.3
R21104 VSS.n8282 VSS.n8281 9.3
R21105 VSS.n8281 VSS.n7455 9.3
R21106 VSS.n7455 VSS.n7454 9.3
R21107 VSS.n8096 VSS.n8095 9.3
R21108 VSS.n8099 VSS.n8098 9.3
R21109 VSS.n8099 VSS.n8090 9.3
R21110 VSS.n8090 VSS.n7460 9.3
R21111 VSS.n8094 VSS.n8093 9.3
R21112 VSS.n8107 VSS.n8106 9.3
R21113 VSS.n8106 VSS.n8105 9.3
R21114 VSS.n8105 VSS.n8104 9.3
R21115 VSS.n8108 VSS.n8082 9.3
R21116 VSS.n8111 VSS.n8077 9.3
R21117 VSS.n8112 VSS.n8111 9.3
R21118 VSS.n8113 VSS.n8112 9.3
R21119 VSS.n8119 VSS.n8118 9.3
R21120 VSS.n8122 VSS.n8121 9.3
R21121 VSS.n8122 VSS.n8072 9.3
R21122 VSS.n8072 VSS.n8071 9.3
R21123 VSS.n8076 VSS.n8075 9.3
R21124 VSS.n8130 VSS.n8129 9.3
R21125 VSS.n8129 VSS.n8128 9.3
R21126 VSS.n8128 VSS.n8127 9.3
R21127 VSS.n8131 VSS.n8063 9.3
R21128 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector VSS.n8058 9.3
R21129 VSS.n8134 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector 9.3
R21130 VSS.n8135 VSS.n8134 9.3
R21131 VSS.n8141 VSS.n8140 9.3
R21132 VSS.n8144 VSS.n8143 9.3
R21133 VSS.n8144 VSS.n8053 9.3
R21134 VSS.n8053 VSS.n8052 9.3
R21135 VSS.n8057 VSS.n8056 9.3
R21136 VSS.n8152 VSS.n8151 9.3
R21137 VSS.n8151 VSS.n8150 9.3
R21138 VSS.n8150 VSS.n8149 9.3
R21139 VSS.n8153 VSS.n8044 9.3
R21140 VSS.n8156 VSS.n8039 9.3
R21141 VSS.n8157 VSS.n8156 9.3
R21142 VSS.n8158 VSS.n8157 9.3
R21143 VSS.n8164 VSS.n8163 9.3
R21144 VSS.n8167 VSS.n8166 9.3
R21145 VSS.n8167 VSS.n8033 9.3
R21146 VSS.n8033 VSS.n8032 9.3
R21147 VSS.n8038 VSS.n8037 9.3
R21148 VSS.n8174 VSS.n8030 9.3
R21149 VSS.n8174 VSS.n8173 9.3
R21150 VSS.n8173 VSS.n8172 9.3
R21151 VSS.n8029 VSS.n8023 9.3
R21152 VSS.n8026 VSS.n8025 9.3
R21153 VSS.n8026 VSS.n8020 9.3
R21154 VSS.n8179 VSS.n8020 9.3
R21155 VSS.n8186 VSS.n8185 9.3
R21156 VSS.n8189 VSS.n8188 9.3
R21157 VSS.n8190 VSS.n8189 9.3
R21158 VSS.n8191 VSS.n8190 9.3
R21159 VSS.n8017 VSS.n8016 9.3
R21160 VSS.n8008 VSS.n8007 9.3
R21161 VSS.n8008 VSS.n7544 9.3
R21162 VSS.n8012 VSS.n7544 9.3
R21163 VSS.n8006 VSS.n8005 9.3
R21164 VSS.n8003 VSS.n7550 9.3
R21165 VSS.n8003 VSS.n8002 9.3
R21166 VSS.n8002 VSS.n8001 9.3
R21167 VSS.n7996 VSS.n7995 9.3
R21168 VSS.n7993 VSS.n7992 9.3
R21169 VSS.n7992 VSS.n7553 9.3
R21170 VSS.n7553 VSS.n7552 9.3
R21171 VSS.n7561 VSS.n7555 9.3
R21172 VSS.n7985 VSS.n7984 9.3
R21173 VSS.n7986 VSS.n7985 9.3
R21174 VSS.n7987 VSS.n7986 9.3
R21175 VSS.n7982 VSS.n7981 9.3
R21176 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector VSS.n7973 9.3
R21177 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector VSS.n7565 9.3
R21178 VSS.n7977 VSS.n7565 9.3
R21179 VSS.n7972 VSS.n7971 9.3
R21180 VSS.n7969 VSS.n7571 9.3
R21181 VSS.n7969 VSS.n7968 9.3
R21182 VSS.n7968 VSS.n7967 9.3
R21183 VSS.n7962 VSS.n7961 9.3
R21184 VSS.n7959 VSS.n7958 9.3
R21185 VSS.n7958 VSS.n7574 9.3
R21186 VSS.n7574 VSS.n7573 9.3
R21187 VSS.n7582 VSS.n7576 9.3
R21188 VSS.n7951 VSS.n7950 9.3
R21189 VSS.n7952 VSS.n7951 9.3
R21190 VSS.n7953 VSS.n7952 9.3
R21191 VSS.n7948 VSS.n7947 9.3
R21192 VSS.n7939 VSS.n7938 9.3
R21193 VSS.n7939 VSS.n7586 9.3
R21194 VSS.n7943 VSS.n7586 9.3
R21195 VSS.n7937 VSS.n7936 9.3
R21196 VSS.n7934 VSS.n7592 9.3
R21197 VSS.n7934 VSS.n7933 9.3
R21198 VSS.n7933 VSS.n7932 9.3
R21199 VSS.n7927 VSS.n7926 9.3
R21200 VSS.n7924 VSS.n7923 9.3
R21201 VSS.n7923 VSS.n7595 9.3
R21202 VSS.n7595 VSS.n7594 9.3
R21203 VSS.n7745 VSS.n7744 9.3
R21204 VSS.n7748 VSS.n7742 9.3
R21205 VSS.n7749 VSS.n7748 9.3
R21206 VSS.n7749 VSS.n7600 9.3
R21207 VSS.n7756 VSS.n7755 9.3
R21208 VSS.n7759 VSS.n7758 9.3
R21209 VSS.n7759 VSS.n7737 9.3
R21210 VSS.n7737 VSS.n7736 9.3
R21211 VSS.n7741 VSS.n7740 9.3
R21212 VSS.n7767 VSS.n7766 9.3
R21213 VSS.n7766 VSS.n7765 9.3
R21214 VSS.n7765 VSS.n7764 9.3
R21215 VSS.n7768 VSS.n7728 9.3
R21216 VSS.n7771 VSS.n7723 9.3
R21217 VSS.n7772 VSS.n7771 9.3
R21218 VSS.n7773 VSS.n7772 9.3
R21219 VSS.n7779 VSS.n7778 9.3
R21220 VSS.n7782 VSS.n7781 9.3
R21221 VSS.n7782 VSS.n7718 9.3
R21222 VSS.n7718 VSS.n7717 9.3
R21223 VSS.n7722 VSS.n7721 9.3
R21224 VSS.n7789 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Collector 9.3
R21225 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Collector VSS.n7788 9.3
R21226 VSS.n7788 VSS.n7787 9.3
R21227 VSS.n7790 VSS.n7709 9.3
R21228 VSS.n7793 VSS.n7704 9.3
R21229 VSS.n7794 VSS.n7793 9.3
R21230 VSS.n7795 VSS.n7794 9.3
R21231 VSS.n7801 VSS.n7800 9.3
R21232 VSS.n7804 VSS.n7803 9.3
R21233 VSS.n7804 VSS.n7699 9.3
R21234 VSS.n7699 VSS.n7698 9.3
R21235 VSS.n7703 VSS.n7702 9.3
R21236 VSS.n7812 VSS.n7811 9.3
R21237 VSS.n7811 VSS.n7810 9.3
R21238 VSS.n7810 VSS.n7809 9.3
R21239 VSS.n7813 VSS.n7690 9.3
R21240 VSS.n7816 VSS.n7685 9.3
R21241 VSS.n7817 VSS.n7816 9.3
R21242 VSS.n7818 VSS.n7817 9.3
R21243 VSS.n7824 VSS.n7823 9.3
R21244 VSS.n7827 VSS.n7826 9.3
R21245 VSS.n7827 VSS.n7679 9.3
R21246 VSS.n7679 VSS.n7678 9.3
R21247 VSS.n7684 VSS.n7683 9.3
R21248 VSS.n7834 VSS.n7676 9.3
R21249 VSS.n7834 VSS.n7833 9.3
R21250 VSS.n7833 VSS.n7832 9.3
R21251 VSS.n7173 VSS.n7008 9.3
R21252 VSS.n7173 VSS.n7172 9.3
R21253 VSS.n7172 VSS.n7171 9.3
R21254 VSS.n7176 VSS.n7175 9.3
R21255 VSS.n9766 VSS.n9765 9.3
R21256 VSS.n9765 VSS.n9665 9.3
R21257 VSS.n9768 VSS.n9767 9.3
R21258 VSS.n9772 VSS.n9771 9.3
R21259 VSS.n9771 VSS.n9770 9.3
R21260 VSS.n9778 VSS.n9777 9.3
R21261 VSS.n9777 VSS.n9776 9.3
R21262 VSS.n9780 VSS.n9779 9.3
R21263 VSS.n9784 VSS.n9783 9.3
R21264 VSS.n9783 VSS.n9782 9.3
R21265 VSS.n9790 VSS.n9789 9.3
R21266 VSS.n9789 VSS.n9788 9.3
R21267 VSS.n9791 VSS.n9736 9.3
R21268 VSS.n9795 VSS.n9735 9.3
R21269 VSS.n9795 VSS.n9794 9.3
R21270 VSS.n9804 VSS.n9802 9.3
R21271 VSS.n9804 VSS.n9803 9.3
R21272 VSS.n9734 VSS.n9676 9.3
R21273 VSS.n9731 VSS.n9678 9.3
R21274 VSS.n9731 VSS.n9675 9.3
R21275 VSS.n9763 VSS.n9762 9.3
R21276 VSS.n9774 VSS.n9773 9.3
R21277 VSS.n9786 VSS.n9785 9.3
R21278 VSS.n9800 VSS.n9799 9.3
R21279 VSS.n9761 VSS.n9760 9.3
R21280 VSS.n9760 VSS.n9640 9.3
R21281 VSS.n9638 VSS.n9637 9.3
R21282 VSS.n9856 VSS.n9855 9.3
R21283 VSS.n9855 VSS.n9575 9.3
R21284 VSS.n9858 VSS.n9857 9.3
R21285 VSS.n9862 VSS.n9861 9.3
R21286 VSS.n9861 VSS.n9860 9.3
R21287 VSS.n9868 VSS.n9867 9.3
R21288 VSS.n9867 VSS.n9866 9.3
R21289 VSS.n9870 VSS.n9869 9.3
R21290 VSS.n9874 VSS.n9873 9.3
R21291 VSS.n9873 VSS.n9872 9.3
R21292 VSS.n9880 VSS.n9879 9.3
R21293 VSS.n9879 VSS.n9878 9.3
R21294 VSS.n9881 VSS.n9826 9.3
R21295 VSS.n9885 VSS.n9825 9.3
R21296 VSS.n9885 VSS.n9884 9.3
R21297 VSS.n9894 VSS.n9892 9.3
R21298 VSS.n9894 VSS.n9893 9.3
R21299 VSS.n9824 VSS.n9586 9.3
R21300 VSS.n9821 VSS.n9588 9.3
R21301 VSS.n9821 VSS.n9585 9.3
R21302 VSS.n9853 VSS.n9852 9.3
R21303 VSS.n9864 VSS.n9863 9.3
R21304 VSS.n9876 VSS.n9875 9.3
R21305 VSS.n9890 VSS.n9889 9.3
R21306 VSS.n9851 VSS.n9850 9.3
R21307 VSS.n9850 VSS.n9550 9.3
R21308 VSS.n9548 VSS.n9547 9.3
R21309 VSS.n9946 VSS.n9945 9.3
R21310 VSS.n9945 VSS.n9485 9.3
R21311 VSS.n9948 VSS.n9947 9.3
R21312 VSS.n9952 VSS.n9951 9.3
R21313 VSS.n9951 VSS.n9950 9.3
R21314 VSS.n9958 VSS.n9957 9.3
R21315 VSS.n9957 VSS.n9956 9.3
R21316 VSS.n9960 VSS.n9959 9.3
R21317 VSS.n9964 VSS.n9963 9.3
R21318 VSS.n9963 VSS.n9962 9.3
R21319 VSS.n9970 VSS.n9969 9.3
R21320 VSS.n9969 VSS.n9968 9.3
R21321 VSS.n9971 VSS.n9916 9.3
R21322 VSS.n9975 VSS.n9915 9.3
R21323 VSS.n9975 VSS.n9974 9.3
R21324 VSS.n9984 VSS.n9982 9.3
R21325 VSS.n9984 VSS.n9983 9.3
R21326 VSS.n9914 VSS.n9496 9.3
R21327 VSS.n9911 VSS.n9498 9.3
R21328 VSS.n9911 VSS.n9495 9.3
R21329 VSS.n9943 VSS.n9942 9.3
R21330 VSS.n9954 VSS.n9953 9.3
R21331 VSS.n9966 VSS.n9965 9.3
R21332 VSS.n9980 VSS.n9979 9.3
R21333 VSS.n9941 VSS.n9940 9.3
R21334 VSS.n9940 VSS.n9460 9.3
R21335 VSS.n9458 VSS.n9457 9.3
R21336 VSS.n10036 VSS.n10035 9.3
R21337 VSS.n10035 VSS.n9395 9.3
R21338 VSS.n10038 VSS.n10037 9.3
R21339 VSS.n10042 VSS.n10041 9.3
R21340 VSS.n10041 VSS.n10040 9.3
R21341 VSS.n10048 VSS.n10047 9.3
R21342 VSS.n10047 VSS.n10046 9.3
R21343 VSS.n10050 VSS.n10049 9.3
R21344 VSS.n10054 VSS.n10053 9.3
R21345 VSS.n10053 VSS.n10052 9.3
R21346 VSS.n10060 VSS.n10059 9.3
R21347 VSS.n10059 VSS.n10058 9.3
R21348 VSS.n10061 VSS.n10006 9.3
R21349 VSS.n10065 VSS.n10005 9.3
R21350 VSS.n10065 VSS.n10064 9.3
R21351 VSS.n10074 VSS.n10072 9.3
R21352 VSS.n10074 VSS.n10073 9.3
R21353 VSS.n10004 VSS.n9406 9.3
R21354 VSS.n10001 VSS.n9408 9.3
R21355 VSS.n10001 VSS.n9405 9.3
R21356 VSS.n10033 VSS.n10032 9.3
R21357 VSS.n10044 VSS.n10043 9.3
R21358 VSS.n10056 VSS.n10055 9.3
R21359 VSS.n10070 VSS.n10069 9.3
R21360 VSS.n10031 VSS.n10030 9.3
R21361 VSS.n10030 VSS.n9370 9.3
R21362 VSS.n9368 VSS.n9367 9.3
R21363 VSS.n10126 VSS.n10125 9.3
R21364 VSS.n10125 VSS.n9305 9.3
R21365 VSS.n10128 VSS.n10127 9.3
R21366 VSS.n10132 VSS.n10131 9.3
R21367 VSS.n10131 VSS.n10130 9.3
R21368 VSS.n10138 VSS.n10137 9.3
R21369 VSS.n10137 VSS.n10136 9.3
R21370 VSS.n10140 VSS.n10139 9.3
R21371 VSS.n10144 VSS.n10143 9.3
R21372 VSS.n10143 VSS.n10142 9.3
R21373 VSS.n10150 VSS.n10149 9.3
R21374 VSS.n10149 VSS.n10148 9.3
R21375 VSS.n10151 VSS.n10096 9.3
R21376 VSS.n10155 VSS.n10095 9.3
R21377 VSS.n10155 VSS.n10154 9.3
R21378 VSS.n10164 VSS.n10162 9.3
R21379 VSS.n10164 VSS.n10163 9.3
R21380 VSS.n10094 VSS.n9316 9.3
R21381 VSS.n10091 VSS.n9318 9.3
R21382 VSS.n10091 VSS.n9315 9.3
R21383 VSS.n10123 VSS.n10122 9.3
R21384 VSS.n10134 VSS.n10133 9.3
R21385 VSS.n10146 VSS.n10145 9.3
R21386 VSS.n10160 VSS.n10159 9.3
R21387 VSS.n10121 VSS.n10120 9.3
R21388 VSS.n10120 VSS.n9280 9.3
R21389 VSS.n9278 VSS.n9277 9.3
R21390 VSS.n10216 VSS.n10215 9.3
R21391 VSS.n10215 VSS.n9215 9.3
R21392 VSS.n10218 VSS.n10217 9.3
R21393 VSS.n10222 VSS.n10221 9.3
R21394 VSS.n10221 VSS.n10220 9.3
R21395 VSS.n10228 VSS.n10227 9.3
R21396 VSS.n10227 VSS.n10226 9.3
R21397 VSS.n10230 VSS.n10229 9.3
R21398 VSS.n10234 VSS.n10233 9.3
R21399 VSS.n10233 VSS.n10232 9.3
R21400 VSS.n10240 VSS.n10239 9.3
R21401 VSS.n10239 VSS.n10238 9.3
R21402 VSS.n10241 VSS.n10186 9.3
R21403 VSS.n10245 VSS.n10185 9.3
R21404 VSS.n10245 VSS.n10244 9.3
R21405 VSS.n10254 VSS.n10252 9.3
R21406 VSS.n10254 VSS.n10253 9.3
R21407 VSS.n10184 VSS.n9226 9.3
R21408 VSS.n10181 VSS.n9228 9.3
R21409 VSS.n10181 VSS.n9225 9.3
R21410 VSS.n10213 VSS.n10212 9.3
R21411 VSS.n10224 VSS.n10223 9.3
R21412 VSS.n10236 VSS.n10235 9.3
R21413 VSS.n10250 VSS.n10249 9.3
R21414 VSS.n10211 VSS.n10210 9.3
R21415 VSS.n10210 VSS.n9190 9.3
R21416 VSS.n9188 VSS.n9187 9.3
R21417 VSS.n8980 VSS.n8978 9.3
R21418 VSS.n8945 VSS.n8942 9.3
R21419 VSS.n8956 VSS.n8954 9.3
R21420 VSS.n8969 VSS.n8966 9.3
R21421 VSS.n9150 VSS.n9149 9.3
R21422 VSS.n9153 VSS.n9152 9.3
R21423 VSS.n9154 VSS.n9153 9.3
R21424 VSS.n9083 VSS.n9081 9.3
R21425 VSS.n9083 VSS.n9082 9.3
R21426 VSS.n9067 VSS.n9065 9.3
R21427 VSS.n9067 VSS.n9066 9.3
R21428 VSS.n9051 VSS.n9049 9.3
R21429 VSS.n9051 VSS.n9050 9.3
R21430 VSS.n9035 VSS.n8981 9.3
R21431 VSS.n9035 VSS.n9034 9.3
R21432 VSS.n9040 VSS.n9039 9.3
R21433 VSS.n9043 VSS.n9041 9.3
R21434 VSS.n9043 VSS.n9042 9.3
R21435 VSS.n9048 VSS.n9047 9.3
R21436 VSS.n9056 VSS.n9055 9.3
R21437 VSS.n9059 VSS.n9057 9.3
R21438 VSS.n9059 VSS.n9058 9.3
R21439 VSS.n9064 VSS.n9063 9.3
R21440 VSS.n9072 VSS.n9071 9.3
R21441 VSS.n9075 VSS.n9073 9.3
R21442 VSS.n9075 VSS.n9074 9.3
R21443 VSS.n9080 VSS.n9079 9.3
R21444 VSS.n9088 VSS.n9087 9.3
R21445 VSS.n9091 VSS.n9089 9.3
R21446 VSS.n9091 VSS.n9090 9.3
R21447 VSS.n9096 VSS.n9095 9.3
R21448 VSS.n10327 VSS.n8976 9.3
R21449 VSS.n10327 VSS.n10326 9.3
R21450 VSS.n10333 VSS.n8970 9.3
R21451 VSS.n10333 VSS.n10332 9.3
R21452 VSS.n8975 VSS.n8972 9.3
R21453 VSS.n10339 VSS.n8964 9.3
R21454 VSS.n10339 VSS.n10338 9.3
R21455 VSS.n10345 VSS.n8957 9.3
R21456 VSS.n10345 VSS.n10344 9.3
R21457 VSS.n8963 VSS.n8959 9.3
R21458 VSS.n10351 VSS.n8952 9.3
R21459 VSS.n10351 VSS.n10350 9.3
R21460 VSS.n10357 VSS.n8946 9.3
R21461 VSS.n10357 VSS.n10356 9.3
R21462 VSS.n8951 VSS.n8948 9.3
R21463 VSS.n10363 VSS.n8940 9.3
R21464 VSS.n10363 VSS.n10362 9.3
R21465 VSS.n8939 VSS.n8937 9.3
R21466 VSS.n10370 VSS.n10369 9.3
R21467 VSS.n10369 VSS.n10368 9.3
R21468 VSS.n10321 VSS.n10320 9.3
R21469 VSS.n10321 VSS.n9180 9.3
R21470 VSS.n9185 VSS.n8930 9.3
R21471 VSS.n5486 VSS.n5477 9.3
R21472 VSS.n5487 VSS.n5486 9.3
R21473 VSS.n5488 VSS.n5487 9.3
R21474 VSS.n5494 VSS.n5493 9.3
R21475 VSS.n5497 VSS.n5496 9.3
R21476 VSS.n5497 VSS.n5472 9.3
R21477 VSS.n5472 VSS.n5471 9.3
R21478 VSS.n5505 VSS.n5504 9.3
R21479 VSS.n5504 VSS.n5503 9.3
R21480 VSS.n5503 VSS.n5502 9.3
R21481 VSS.n5506 VSS.n5463 9.3
R21482 VSS.n5509 VSS.n5458 9.3
R21483 VSS.n5510 VSS.n5509 9.3
R21484 VSS.n5511 VSS.n5510 9.3
R21485 sky130_asc_pnp_05v5_W3p40L3p40_8_2/xm1/Collector VSS.n5519 9.3
R21486 sky130_asc_pnp_05v5_W3p40L3p40_8_2/xm1/Collector VSS.n5453 9.3
R21487 VSS.n5453 VSS.n5452 9.3
R21488 VSS.n5457 VSS.n5456 9.3
R21489 VSS.n5527 VSS.n5526 9.3
R21490 VSS.n5526 VSS.n5525 9.3
R21491 VSS.n5525 VSS.n5524 9.3
R21492 VSS.n5531 VSS.n5439 9.3
R21493 VSS.n5532 VSS.n5531 9.3
R21494 VSS.n5533 VSS.n5532 9.3
R21495 VSS.n5539 VSS.n5538 9.3
R21496 VSS.n5542 VSS.n5541 9.3
R21497 VSS.n5542 VSS.n5434 9.3
R21498 VSS.n5434 VSS.n5433 9.3
R21499 VSS.n5550 VSS.n5549 9.3
R21500 VSS.n5549 VSS.n5548 9.3
R21501 VSS.n5548 VSS.n5547 9.3
R21502 VSS.n5551 VSS.n5425 9.3
R21503 VSS.n5554 VSS.n5419 9.3
R21504 VSS.n5555 VSS.n5554 9.3
R21505 VSS.n5556 VSS.n5555 9.3
R21506 VSS.n5565 VSS.n5564 9.3
R21507 VSS.n5565 VSS.n5417 9.3
R21508 VSS.n5422 VSS.n5417 9.3
R21509 VSS.n5483 VSS.n3635 9.3
R21510 VSS.n5476 VSS.n5475 9.3
R21511 VSS.n5517 VSS.n5516 9.3
R21512 VSS.n5528 VSS.n5444 9.3
R21513 VSS.n5438 VSS.n5437 9.3
R21514 VSS.n5562 VSS.n5561 9.3
R21515 VSS.n5577 VSS.n5576 9.3
R21516 VSS.n5574 VSS.n5573 9.3
R21517 VSS.n5573 VSS.n5572 9.3
R21518 VSS.n5572 VSS.n5571 9.3
R21519 VSS.n5411 VSS.n3691 9.3
R21520 VSS.n5408 VSS.n3697 9.3
R21521 VSS.n3697 VSS.n3696 9.3
R21522 VSS.n3696 VSS.n3695 9.3
R21523 VSS.n5407 VSS.n5406 9.3
R21524 VSS.n5397 VSS.n5396 9.3
R21525 VSS.n5397 VSS.n3701 9.3
R21526 VSS.n5401 VSS.n3701 9.3
R21527 VSS.n5395 VSS.n5394 9.3
R21528 VSS.n5392 VSS.n3708 9.3
R21529 VSS.n5392 VSS.n5391 9.3
R21530 VSS.n5391 VSS.n5390 9.3
R21531 VSS.n5385 VSS.n5384 9.3
R21532 VSS.n5382 VSS.n5381 9.3
R21533 VSS.n5381 VSS.n3711 9.3
R21534 VSS.n3711 VSS.n3710 9.3
R21535 VSS.n3719 VSS.n3713 9.3
R21536 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector VSS.n5374 9.3
R21537 VSS.n5375 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector 9.3
R21538 VSS.n5376 VSS.n5375 9.3
R21539 VSS.n5372 VSS.n5371 9.3
R21540 VSS.n5363 VSS.n5362 9.3
R21541 VSS.n5363 VSS.n3723 9.3
R21542 VSS.n5367 VSS.n3723 9.3
R21543 VSS.n5361 VSS.n5360 9.3
R21544 VSS.n5358 VSS.n3729 9.3
R21545 VSS.n5358 VSS.n5357 9.3
R21546 VSS.n5357 VSS.n5356 9.3
R21547 VSS.n5351 VSS.n5350 9.3
R21548 VSS.n5348 VSS.n5347 9.3
R21549 VSS.n5347 VSS.n3732 9.3
R21550 VSS.n3732 VSS.n3731 9.3
R21551 VSS.n3740 VSS.n3734 9.3
R21552 VSS.n5340 VSS.n5339 9.3
R21553 VSS.n5341 VSS.n5340 9.3
R21554 VSS.n5342 VSS.n5341 9.3
R21555 VSS.n5337 VSS.n5336 9.3
R21556 VSS.n5328 VSS.n5327 9.3
R21557 VSS.n5328 VSS.n3744 9.3
R21558 VSS.n5332 VSS.n3744 9.3
R21559 VSS.n5326 VSS.n5325 9.3
R21560 VSS.n5323 VSS.n3750 9.3
R21561 VSS.n5323 VSS.n5322 9.3
R21562 VSS.n5322 VSS.n5321 9.3
R21563 VSS.n5126 VSS.n3754 9.3
R21564 VSS.n5136 VSS.n5135 9.3
R21565 VSS.n5135 VSS.n5134 9.3
R21566 VSS.n5134 VSS.n5133 9.3
R21567 VSS.n5137 VSS.n5125 9.3
R21568 VSS.n5140 VSS.n5120 9.3
R21569 VSS.n5141 VSS.n5140 9.3
R21570 VSS.n5142 VSS.n5141 9.3
R21571 VSS.n5148 VSS.n5147 9.3
R21572 VSS.n5151 VSS.n5150 9.3
R21573 VSS.n5151 VSS.n5115 9.3
R21574 VSS.n5115 VSS.n5114 9.3
R21575 VSS.n5119 VSS.n5118 9.3
R21576 VSS.n5159 VSS.n5158 9.3
R21577 VSS.n5158 VSS.n5157 9.3
R21578 VSS.n5157 VSS.n5156 9.3
R21579 VSS.n5160 VSS.n5106 9.3
R21580 VSS.n5163 VSS.n5101 9.3
R21581 VSS.n5164 VSS.n5163 9.3
R21582 VSS.n5165 VSS.n5164 9.3
R21583 VSS.n5171 VSS.n5170 9.3
R21584 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector VSS.n5173 9.3
R21585 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector VSS.n5096 9.3
R21586 VSS.n5096 VSS.n5095 9.3
R21587 VSS.n5100 VSS.n5099 9.3
R21588 VSS.n5181 VSS.n5180 9.3
R21589 VSS.n5180 VSS.n5179 9.3
R21590 VSS.n5179 VSS.n5178 9.3
R21591 VSS.n5182 VSS.n5087 9.3
R21592 VSS.n5185 VSS.n5082 9.3
R21593 VSS.n5186 VSS.n5185 9.3
R21594 VSS.n5187 VSS.n5186 9.3
R21595 VSS.n5193 VSS.n5192 9.3
R21596 VSS.n5196 VSS.n5195 9.3
R21597 VSS.n5196 VSS.n5077 9.3
R21598 VSS.n5077 VSS.n5076 9.3
R21599 VSS.n5081 VSS.n5080 9.3
R21600 VSS.n5204 VSS.n5203 9.3
R21601 VSS.n5203 VSS.n5202 9.3
R21602 VSS.n5202 VSS.n5201 9.3
R21603 VSS.n5205 VSS.n5068 9.3
R21604 VSS.n5208 VSS.n5062 9.3
R21605 VSS.n5209 VSS.n5208 9.3
R21606 VSS.n5210 VSS.n5209 9.3
R21607 VSS.n5216 VSS.n5215 9.3
R21608 VSS.n5219 VSS.n5218 9.3
R21609 VSS.n5219 VSS.n5060 9.3
R21610 VSS.n5065 VSS.n5060 9.3
R21611 VSS.n5231 VSS.n5230 9.3
R21612 VSS.n5228 VSS.n5227 9.3
R21613 VSS.n5227 VSS.n5226 9.3
R21614 VSS.n5226 VSS.n5225 9.3
R21615 VSS.n5054 VSS.n3832 9.3
R21616 VSS.n5051 VSS.n3838 9.3
R21617 VSS.n3838 VSS.n3837 9.3
R21618 VSS.n3837 VSS.n3836 9.3
R21619 VSS.n5050 VSS.n5049 9.3
R21620 VSS.n5040 VSS.n5039 9.3
R21621 VSS.n5040 VSS.n3842 9.3
R21622 VSS.n5044 VSS.n3842 9.3
R21623 VSS.n5038 VSS.n5037 9.3
R21624 VSS.n5035 VSS.n3849 9.3
R21625 VSS.n5035 VSS.n5034 9.3
R21626 VSS.n5034 VSS.n5033 9.3
R21627 VSS.n5028 VSS.n5027 9.3
R21628 VSS.n5025 VSS.n5024 9.3
R21629 VSS.n5024 VSS.n3852 9.3
R21630 VSS.n3852 VSS.n3851 9.3
R21631 VSS.n3860 VSS.n3854 9.3
R21632 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector VSS.n5017 9.3
R21633 VSS.n5018 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector 9.3
R21634 VSS.n5019 VSS.n5018 9.3
R21635 VSS.n5015 VSS.n5014 9.3
R21636 VSS.n5006 VSS.n5005 9.3
R21637 VSS.n5006 VSS.n3864 9.3
R21638 VSS.n5010 VSS.n3864 9.3
R21639 VSS.n5004 VSS.n5003 9.3
R21640 VSS.n5001 VSS.n3870 9.3
R21641 VSS.n5001 VSS.n5000 9.3
R21642 VSS.n5000 VSS.n4999 9.3
R21643 VSS.n4994 VSS.n4993 9.3
R21644 VSS.n4991 VSS.n4990 9.3
R21645 VSS.n4990 VSS.n3873 9.3
R21646 VSS.n3873 VSS.n3872 9.3
R21647 VSS.n3881 VSS.n3875 9.3
R21648 VSS.n4983 VSS.n4982 9.3
R21649 VSS.n4984 VSS.n4983 9.3
R21650 VSS.n4985 VSS.n4984 9.3
R21651 VSS.n4980 VSS.n4979 9.3
R21652 VSS.n4971 VSS.n4970 9.3
R21653 VSS.n4971 VSS.n3885 9.3
R21654 VSS.n4975 VSS.n3885 9.3
R21655 VSS.n4969 VSS.n4968 9.3
R21656 VSS.n4966 VSS.n3891 9.3
R21657 VSS.n4966 VSS.n4965 9.3
R21658 VSS.n4965 VSS.n4964 9.3
R21659 VSS.n4769 VSS.n3895 9.3
R21660 VSS.n4779 VSS.n4778 9.3
R21661 VSS.n4778 VSS.n4777 9.3
R21662 VSS.n4777 VSS.n4776 9.3
R21663 VSS.n4780 VSS.n4768 9.3
R21664 VSS.n4783 VSS.n4763 9.3
R21665 VSS.n4784 VSS.n4783 9.3
R21666 VSS.n4785 VSS.n4784 9.3
R21667 VSS.n4791 VSS.n4790 9.3
R21668 VSS.n4794 VSS.n4793 9.3
R21669 VSS.n4794 VSS.n4758 9.3
R21670 VSS.n4758 VSS.n4757 9.3
R21671 VSS.n4762 VSS.n4761 9.3
R21672 VSS.n4802 VSS.n4801 9.3
R21673 VSS.n4801 VSS.n4800 9.3
R21674 VSS.n4800 VSS.n4799 9.3
R21675 VSS.n4803 VSS.n4749 9.3
R21676 VSS.n4806 VSS.n4744 9.3
R21677 VSS.n4807 VSS.n4806 9.3
R21678 VSS.n4808 VSS.n4807 9.3
R21679 VSS.n4814 VSS.n4813 9.3
R21680 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector VSS.n4816 9.3
R21681 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector VSS.n4739 9.3
R21682 VSS.n4739 VSS.n4738 9.3
R21683 VSS.n4743 VSS.n4742 9.3
R21684 VSS.n4824 VSS.n4823 9.3
R21685 VSS.n4823 VSS.n4822 9.3
R21686 VSS.n4822 VSS.n4821 9.3
R21687 VSS.n4825 VSS.n4730 9.3
R21688 VSS.n4828 VSS.n4725 9.3
R21689 VSS.n4829 VSS.n4828 9.3
R21690 VSS.n4830 VSS.n4829 9.3
R21691 VSS.n4836 VSS.n4835 9.3
R21692 VSS.n4839 VSS.n4838 9.3
R21693 VSS.n4839 VSS.n4720 9.3
R21694 VSS.n4720 VSS.n4719 9.3
R21695 VSS.n4724 VSS.n4723 9.3
R21696 VSS.n4847 VSS.n4846 9.3
R21697 VSS.n4846 VSS.n4845 9.3
R21698 VSS.n4845 VSS.n4844 9.3
R21699 VSS.n4848 VSS.n4711 9.3
R21700 VSS.n4851 VSS.n4705 9.3
R21701 VSS.n4852 VSS.n4851 9.3
R21702 VSS.n4853 VSS.n4852 9.3
R21703 VSS.n4859 VSS.n4858 9.3
R21704 VSS.n4862 VSS.n4861 9.3
R21705 VSS.n4862 VSS.n4703 9.3
R21706 VSS.n4708 VSS.n4703 9.3
R21707 VSS.n4874 VSS.n4873 9.3
R21708 VSS.n4871 VSS.n4870 9.3
R21709 VSS.n4870 VSS.n4869 9.3
R21710 VSS.n4869 VSS.n4868 9.3
R21711 VSS.n4697 VSS.n3973 9.3
R21712 VSS.n4694 VSS.n3979 9.3
R21713 VSS.n3979 VSS.n3978 9.3
R21714 VSS.n3978 VSS.n3977 9.3
R21715 VSS.n4693 VSS.n4692 9.3
R21716 VSS.n4683 VSS.n4682 9.3
R21717 VSS.n4683 VSS.n3983 9.3
R21718 VSS.n4687 VSS.n3983 9.3
R21719 VSS.n4681 VSS.n4680 9.3
R21720 VSS.n4678 VSS.n3990 9.3
R21721 VSS.n4678 VSS.n4677 9.3
R21722 VSS.n4677 VSS.n4676 9.3
R21723 VSS.n4671 VSS.n4670 9.3
R21724 VSS.n4668 VSS.n4667 9.3
R21725 VSS.n4667 VSS.n3993 9.3
R21726 VSS.n3993 VSS.n3992 9.3
R21727 VSS.n4001 VSS.n3995 9.3
R21728 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector VSS.n4660 9.3
R21729 VSS.n4661 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector 9.3
R21730 VSS.n4662 VSS.n4661 9.3
R21731 VSS.n4658 VSS.n4657 9.3
R21732 VSS.n4649 VSS.n4648 9.3
R21733 VSS.n4649 VSS.n4005 9.3
R21734 VSS.n4653 VSS.n4005 9.3
R21735 VSS.n4647 VSS.n4646 9.3
R21736 VSS.n4644 VSS.n4011 9.3
R21737 VSS.n4644 VSS.n4643 9.3
R21738 VSS.n4643 VSS.n4642 9.3
R21739 VSS.n4637 VSS.n4636 9.3
R21740 VSS.n4634 VSS.n4633 9.3
R21741 VSS.n4633 VSS.n4014 9.3
R21742 VSS.n4014 VSS.n4013 9.3
R21743 VSS.n4022 VSS.n4016 9.3
R21744 VSS.n4626 VSS.n4625 9.3
R21745 VSS.n4627 VSS.n4626 9.3
R21746 VSS.n4628 VSS.n4627 9.3
R21747 VSS.n4623 VSS.n4622 9.3
R21748 VSS.n4614 VSS.n4613 9.3
R21749 VSS.n4614 VSS.n4026 9.3
R21750 VSS.n4618 VSS.n4026 9.3
R21751 VSS.n4612 VSS.n4611 9.3
R21752 VSS.n4609 VSS.n4032 9.3
R21753 VSS.n4609 VSS.n4608 9.3
R21754 VSS.n4608 VSS.n4607 9.3
R21755 VSS.n4412 VSS.n4036 9.3
R21756 VSS.n4422 VSS.n4421 9.3
R21757 VSS.n4421 VSS.n4420 9.3
R21758 VSS.n4420 VSS.n4419 9.3
R21759 VSS.n4423 VSS.n4411 9.3
R21760 VSS.n4426 VSS.n4406 9.3
R21761 VSS.n4427 VSS.n4426 9.3
R21762 VSS.n4428 VSS.n4427 9.3
R21763 VSS.n4434 VSS.n4433 9.3
R21764 VSS.n4437 VSS.n4436 9.3
R21765 VSS.n4437 VSS.n4401 9.3
R21766 VSS.n4401 VSS.n4400 9.3
R21767 VSS.n4405 VSS.n4404 9.3
R21768 VSS.n4445 VSS.n4444 9.3
R21769 VSS.n4444 VSS.n4443 9.3
R21770 VSS.n4443 VSS.n4442 9.3
R21771 VSS.n4446 VSS.n4392 9.3
R21772 VSS.n4449 VSS.n4387 9.3
R21773 VSS.n4450 VSS.n4449 9.3
R21774 VSS.n4451 VSS.n4450 9.3
R21775 VSS.n4457 VSS.n4456 9.3
R21776 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector VSS.n4459 9.3
R21777 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector VSS.n4382 9.3
R21778 VSS.n4382 VSS.n4381 9.3
R21779 VSS.n4386 VSS.n4385 9.3
R21780 VSS.n4467 VSS.n4466 9.3
R21781 VSS.n4466 VSS.n4465 9.3
R21782 VSS.n4465 VSS.n4464 9.3
R21783 VSS.n4468 VSS.n4373 9.3
R21784 VSS.n4471 VSS.n4368 9.3
R21785 VSS.n4472 VSS.n4471 9.3
R21786 VSS.n4473 VSS.n4472 9.3
R21787 VSS.n4479 VSS.n4478 9.3
R21788 VSS.n4482 VSS.n4481 9.3
R21789 VSS.n4482 VSS.n4363 9.3
R21790 VSS.n4363 VSS.n4362 9.3
R21791 VSS.n4367 VSS.n4366 9.3
R21792 VSS.n4490 VSS.n4489 9.3
R21793 VSS.n4489 VSS.n4488 9.3
R21794 VSS.n4488 VSS.n4487 9.3
R21795 VSS.n4491 VSS.n4354 9.3
R21796 VSS.n4494 VSS.n4348 9.3
R21797 VSS.n4495 VSS.n4494 9.3
R21798 VSS.n4496 VSS.n4495 9.3
R21799 VSS.n4502 VSS.n4501 9.3
R21800 VSS.n4505 VSS.n4504 9.3
R21801 VSS.n4505 VSS.n4346 9.3
R21802 VSS.n4351 VSS.n4346 9.3
R21803 VSS.n4517 VSS.n4516 9.3
R21804 VSS.n4514 VSS.n4513 9.3
R21805 VSS.n4513 VSS.n4512 9.3
R21806 VSS.n4512 VSS.n4511 9.3
R21807 VSS.n4340 VSS.n4114 9.3
R21808 VSS.n4337 VSS.n4120 9.3
R21809 VSS.n4120 VSS.n4119 9.3
R21810 VSS.n4119 VSS.n4118 9.3
R21811 VSS.n4336 VSS.n4335 9.3
R21812 VSS.n4326 VSS.n4325 9.3
R21813 VSS.n4326 VSS.n4124 9.3
R21814 VSS.n4330 VSS.n4124 9.3
R21815 VSS.n4324 VSS.n4323 9.3
R21816 VSS.n4321 VSS.n4131 9.3
R21817 VSS.n4321 VSS.n4320 9.3
R21818 VSS.n4320 VSS.n4319 9.3
R21819 VSS.n4314 VSS.n4313 9.3
R21820 VSS.n4311 VSS.n4310 9.3
R21821 VSS.n4310 VSS.n4134 9.3
R21822 VSS.n4134 VSS.n4133 9.3
R21823 VSS.n4142 VSS.n4136 9.3
R21824 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Collector VSS.n4303 9.3
R21825 VSS.n4304 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Collector 9.3
R21826 VSS.n4305 VSS.n4304 9.3
R21827 VSS.n4301 VSS.n4300 9.3
R21828 VSS.n4292 VSS.n4291 9.3
R21829 VSS.n4292 VSS.n4146 9.3
R21830 VSS.n4296 VSS.n4146 9.3
R21831 VSS.n4290 VSS.n4289 9.3
R21832 VSS.n4287 VSS.n4152 9.3
R21833 VSS.n4287 VSS.n4286 9.3
R21834 VSS.n4286 VSS.n4285 9.3
R21835 VSS.n4280 VSS.n4279 9.3
R21836 VSS.n4277 VSS.n4276 9.3
R21837 VSS.n4276 VSS.n4155 9.3
R21838 VSS.n4155 VSS.n4154 9.3
R21839 VSS.n4163 VSS.n4157 9.3
R21840 VSS.n4269 VSS.n4268 9.3
R21841 VSS.n4270 VSS.n4269 9.3
R21842 VSS.n4271 VSS.n4270 9.3
R21843 VSS.n4266 VSS.n4265 9.3
R21844 VSS.n4257 VSS.n4256 9.3
R21845 VSS.n4257 VSS.n4167 9.3
R21846 VSS.n4261 VSS.n4167 9.3
R21847 VSS.n4255 VSS.n4254 9.3
R21848 VSS.n4252 VSS.n4173 9.3
R21849 VSS.n4252 VSS.n4251 9.3
R21850 VSS.n4251 VSS.n4250 9.3
R21851 VSS.n5662 VSS.n5661 9.3
R21852 VSS.n5661 VSS.n5660 9.3
R21853 VSS.n5660 VSS.n5659 9.3
R21854 VSS.n3646 VSS.n3645 9.3
R21855 VSS.n3223 VSS.n3221 9.3
R21856 VSS.n3223 VSS.n3222 9.3
R21857 VSS.n3220 VSS.n3219 9.3
R21858 VSS.n3215 VSS.n3213 9.3
R21859 VSS.n3215 VSS.n3214 9.3
R21860 VSS.n3207 VSS.n3205 9.3
R21861 VSS.n3207 VSS.n3206 9.3
R21862 VSS.n3204 VSS.n3203 9.3
R21863 VSS.n3199 VSS.n3197 9.3
R21864 VSS.n3199 VSS.n3198 9.3
R21865 VSS.n3191 VSS.n3189 9.3
R21866 VSS.n3191 VSS.n3190 9.3
R21867 VSS.n3188 VSS.n3187 9.3
R21868 VSS.n3183 VSS.n3181 9.3
R21869 VSS.n3183 VSS.n3182 9.3
R21870 VSS.n3175 VSS.n3174 9.3
R21871 VSS.n3175 VSS.n3141 9.3
R21872 VSS.n6602 VSS.n3137 9.3
R21873 VSS.n3138 VSS.n3136 9.3
R21874 VSS.n6534 VSS.n3138 9.3
R21875 VSS.n3228 VSS.n3227 9.3
R21876 VSS.n3212 VSS.n3211 9.3
R21877 VSS.n3196 VSS.n3195 9.3
R21878 VSS.n3180 VSS.n3179 9.3
R21879 VSS.n6595 VSS.n6594 9.3
R21880 VSS.n6596 VSS.n6595 9.3
R21881 VSS.n6592 VSS.n6591 9.3
R21882 VSS.n6474 VSS.n3275 9.3
R21883 VSS.n6474 VSS.n6473 9.3
R21884 VSS.n3274 VSS.n3271 9.3
R21885 VSS.n6480 VSS.n3269 9.3
R21886 VSS.n6480 VSS.n6479 9.3
R21887 VSS.n6486 VSS.n3262 9.3
R21888 VSS.n6486 VSS.n6485 9.3
R21889 VSS.n3261 VSS.n3259 9.3
R21890 VSS.n6492 VSS.n3257 9.3
R21891 VSS.n6492 VSS.n6491 9.3
R21892 VSS.n6498 VSS.n3251 9.3
R21893 VSS.n6498 VSS.n6497 9.3
R21894 VSS.n3250 VSS.n3247 9.3
R21895 VSS.n6504 VSS.n3245 9.3
R21896 VSS.n6504 VSS.n6503 9.3
R21897 VSS.n6510 VSS.n3239 9.3
R21898 VSS.n6510 VSS.n6509 9.3
R21899 VSS.n3238 VSS.n3236 9.3
R21900 VSS.n6517 VSS.n6516 9.3
R21901 VSS.n6516 VSS.n6515 9.3
R21902 VSS.n3280 VSS.n3277 9.3
R21903 VSS.n3268 VSS.n3264 9.3
R21904 VSS.n3256 VSS.n3253 9.3
R21905 VSS.n3244 VSS.n3241 9.3
R21906 VSS.n6468 VSS.n3281 9.3
R21907 VSS.n6468 VSS.n6467 9.3
R21908 VSS.n3286 VSS.n3284 9.3
R21909 VSS.n6352 VSS.n3333 9.3
R21910 VSS.n6352 VSS.n6351 9.3
R21911 VSS.n3332 VSS.n3329 9.3
R21912 VSS.n6358 VSS.n3327 9.3
R21913 VSS.n6358 VSS.n6357 9.3
R21914 VSS.n6364 VSS.n3320 9.3
R21915 VSS.n6364 VSS.n6363 9.3
R21916 VSS.n3319 VSS.n3317 9.3
R21917 VSS.n6370 VSS.n3315 9.3
R21918 VSS.n6370 VSS.n6369 9.3
R21919 VSS.n6376 VSS.n3309 9.3
R21920 VSS.n6376 VSS.n6375 9.3
R21921 VSS.n3308 VSS.n3305 9.3
R21922 VSS.n6382 VSS.n3303 9.3
R21923 VSS.n6382 VSS.n6381 9.3
R21924 VSS.n6388 VSS.n3297 9.3
R21925 VSS.n6388 VSS.n6387 9.3
R21926 VSS.n3296 VSS.n3294 9.3
R21927 VSS.n6395 VSS.n6394 9.3
R21928 VSS.n6394 VSS.n6393 9.3
R21929 VSS.n3338 VSS.n3335 9.3
R21930 VSS.n3326 VSS.n3322 9.3
R21931 VSS.n3314 VSS.n3311 9.3
R21932 VSS.n3302 VSS.n3299 9.3
R21933 VSS.n6346 VSS.n3339 9.3
R21934 VSS.n6346 VSS.n6345 9.3
R21935 VSS.n3344 VSS.n3342 9.3
R21936 VSS.n6230 VSS.n3391 9.3
R21937 VSS.n6230 VSS.n6229 9.3
R21938 VSS.n3390 VSS.n3387 9.3
R21939 VSS.n6236 VSS.n3385 9.3
R21940 VSS.n6236 VSS.n6235 9.3
R21941 VSS.n6242 VSS.n3378 9.3
R21942 VSS.n6242 VSS.n6241 9.3
R21943 VSS.n3377 VSS.n3375 9.3
R21944 VSS.n6248 VSS.n3373 9.3
R21945 VSS.n6248 VSS.n6247 9.3
R21946 VSS.n6254 VSS.n3367 9.3
R21947 VSS.n6254 VSS.n6253 9.3
R21948 VSS.n3366 VSS.n3363 9.3
R21949 VSS.n6260 VSS.n3361 9.3
R21950 VSS.n6260 VSS.n6259 9.3
R21951 VSS.n6266 VSS.n3355 9.3
R21952 VSS.n6266 VSS.n6265 9.3
R21953 VSS.n3354 VSS.n3352 9.3
R21954 VSS.n6273 VSS.n6272 9.3
R21955 VSS.n6272 VSS.n6271 9.3
R21956 VSS.n3396 VSS.n3393 9.3
R21957 VSS.n3384 VSS.n3380 9.3
R21958 VSS.n3372 VSS.n3369 9.3
R21959 VSS.n3360 VSS.n3357 9.3
R21960 VSS.n6224 VSS.n3397 9.3
R21961 VSS.n6224 VSS.n6223 9.3
R21962 VSS.n3402 VSS.n3400 9.3
R21963 VSS.n6108 VSS.n3449 9.3
R21964 VSS.n6108 VSS.n6107 9.3
R21965 VSS.n3448 VSS.n3445 9.3
R21966 VSS.n6114 VSS.n3443 9.3
R21967 VSS.n6114 VSS.n6113 9.3
R21968 VSS.n6120 VSS.n3436 9.3
R21969 VSS.n6120 VSS.n6119 9.3
R21970 VSS.n3435 VSS.n3433 9.3
R21971 VSS.n6126 VSS.n3431 9.3
R21972 VSS.n6126 VSS.n6125 9.3
R21973 VSS.n6132 VSS.n3425 9.3
R21974 VSS.n6132 VSS.n6131 9.3
R21975 VSS.n3424 VSS.n3421 9.3
R21976 VSS.n6138 VSS.n3419 9.3
R21977 VSS.n6138 VSS.n6137 9.3
R21978 VSS.n6144 VSS.n3413 9.3
R21979 VSS.n6144 VSS.n6143 9.3
R21980 VSS.n3412 VSS.n3410 9.3
R21981 VSS.n6151 VSS.n6150 9.3
R21982 VSS.n6150 VSS.n6149 9.3
R21983 VSS.n3454 VSS.n3451 9.3
R21984 VSS.n3442 VSS.n3438 9.3
R21985 VSS.n3430 VSS.n3427 9.3
R21986 VSS.n3418 VSS.n3415 9.3
R21987 VSS.n6102 VSS.n3455 9.3
R21988 VSS.n6102 VSS.n6101 9.3
R21989 VSS.n3460 VSS.n3458 9.3
R21990 VSS.n5986 VSS.n3507 9.3
R21991 VSS.n5986 VSS.n5985 9.3
R21992 VSS.n3506 VSS.n3503 9.3
R21993 VSS.n5992 VSS.n3501 9.3
R21994 VSS.n5992 VSS.n5991 9.3
R21995 VSS.n5998 VSS.n3494 9.3
R21996 VSS.n5998 VSS.n5997 9.3
R21997 VSS.n3493 VSS.n3491 9.3
R21998 VSS.n6004 VSS.n3489 9.3
R21999 VSS.n6004 VSS.n6003 9.3
R22000 VSS.n6010 VSS.n3483 9.3
R22001 VSS.n6010 VSS.n6009 9.3
R22002 VSS.n3482 VSS.n3479 9.3
R22003 VSS.n6016 VSS.n3477 9.3
R22004 VSS.n6016 VSS.n6015 9.3
R22005 VSS.n6022 VSS.n3471 9.3
R22006 VSS.n6022 VSS.n6021 9.3
R22007 VSS.n3470 VSS.n3468 9.3
R22008 VSS.n6029 VSS.n6028 9.3
R22009 VSS.n6028 VSS.n6027 9.3
R22010 VSS.n3512 VSS.n3509 9.3
R22011 VSS.n3500 VSS.n3496 9.3
R22012 VSS.n3488 VSS.n3485 9.3
R22013 VSS.n3476 VSS.n3473 9.3
R22014 VSS.n5980 VSS.n3513 9.3
R22015 VSS.n5980 VSS.n5979 9.3
R22016 VSS.n3518 VSS.n3516 9.3
R22017 VSS.n5864 VSS.n3565 9.3
R22018 VSS.n5864 VSS.n5863 9.3
R22019 VSS.n3564 VSS.n3561 9.3
R22020 VSS.n5870 VSS.n3559 9.3
R22021 VSS.n5870 VSS.n5869 9.3
R22022 VSS.n5876 VSS.n3552 9.3
R22023 VSS.n5876 VSS.n5875 9.3
R22024 VSS.n3551 VSS.n3549 9.3
R22025 VSS.n5882 VSS.n3547 9.3
R22026 VSS.n5882 VSS.n5881 9.3
R22027 VSS.n5888 VSS.n3541 9.3
R22028 VSS.n5888 VSS.n5887 9.3
R22029 VSS.n3540 VSS.n3537 9.3
R22030 VSS.n5894 VSS.n3535 9.3
R22031 VSS.n5894 VSS.n5893 9.3
R22032 VSS.n5900 VSS.n3529 9.3
R22033 VSS.n5900 VSS.n5899 9.3
R22034 VSS.n3528 VSS.n3526 9.3
R22035 VSS.n5907 VSS.n5906 9.3
R22036 VSS.n5906 VSS.n5905 9.3
R22037 VSS.n3570 VSS.n3567 9.3
R22038 VSS.n3558 VSS.n3554 9.3
R22039 VSS.n3546 VSS.n3543 9.3
R22040 VSS.n3534 VSS.n3531 9.3
R22041 VSS.n5858 VSS.n3571 9.3
R22042 VSS.n5858 VSS.n5857 9.3
R22043 VSS.n3576 VSS.n3574 9.3
R22044 VSS.n5742 VSS.n3623 9.3
R22045 VSS.n5742 VSS.n5741 9.3
R22046 VSS.n3622 VSS.n3619 9.3
R22047 VSS.n5748 VSS.n3617 9.3
R22048 VSS.n5748 VSS.n5747 9.3
R22049 VSS.n5754 VSS.n3610 9.3
R22050 VSS.n5754 VSS.n5753 9.3
R22051 VSS.n3609 VSS.n3607 9.3
R22052 VSS.n5760 VSS.n3605 9.3
R22053 VSS.n5760 VSS.n5759 9.3
R22054 VSS.n5766 VSS.n3599 9.3
R22055 VSS.n5766 VSS.n5765 9.3
R22056 VSS.n3598 VSS.n3595 9.3
R22057 VSS.n5772 VSS.n3593 9.3
R22058 VSS.n5772 VSS.n5771 9.3
R22059 VSS.n5778 VSS.n3587 9.3
R22060 VSS.n5778 VSS.n5777 9.3
R22061 VSS.n3586 VSS.n3584 9.3
R22062 VSS.n5785 VSS.n5784 9.3
R22063 VSS.n5784 VSS.n5783 9.3
R22064 VSS.n3628 VSS.n3625 9.3
R22065 VSS.n3616 VSS.n3612 9.3
R22066 VSS.n3604 VSS.n3601 9.3
R22067 VSS.n3592 VSS.n3589 9.3
R22068 VSS.n5736 VSS.n3629 9.3
R22069 VSS.n5736 VSS.n5735 9.3
R22070 VSS.n3634 VSS.n3632 9.3
R22071 VSS.n2887 VSS.n2886 9.3
R22072 VSS.n2887 VSS.n2867 9.3
R22073 VSS.n2867 VSS.n2866 9.3
R22074 VSS.n2871 VSS.n2870 9.3
R22075 VSS.n2895 VSS.n2894 9.3
R22076 VSS.n2894 VSS.n2893 9.3
R22077 VSS.n2893 VSS.n2892 9.3
R22078 VSS.n2899 VSS.n2853 9.3
R22079 VSS.n2900 VSS.n2899 9.3
R22080 VSS.n2901 VSS.n2900 9.3
R22081 VSS.n2907 VSS.n2906 9.3
R22082 VSS.n2910 VSS.n2909 9.3
R22083 VSS.n2910 VSS.n2848 9.3
R22084 VSS.n2848 VSS.n2847 9.3
R22085 VSS.n2917 sky130_asc_pnp_05v5_W3p40L3p40_7_0/xm1/Collector 9.3
R22086 sky130_asc_pnp_05v5_W3p40L3p40_7_0/xm1/Collector VSS.n2916 9.3
R22087 VSS.n2916 VSS.n2915 9.3
R22088 VSS.n2918 VSS.n2839 9.3
R22089 VSS.n2921 VSS.n2834 9.3
R22090 VSS.n2922 VSS.n2921 9.3
R22091 VSS.n2923 VSS.n2922 9.3
R22092 VSS.n2932 VSS.n2931 9.3
R22093 VSS.n2932 VSS.n2829 9.3
R22094 VSS.n2829 VSS.n2828 9.3
R22095 VSS.n2833 VSS.n2832 9.3
R22096 VSS.n2940 VSS.n2939 9.3
R22097 VSS.n2939 VSS.n2938 9.3
R22098 VSS.n2938 VSS.n2937 9.3
R22099 VSS.n2944 VSS.n2815 9.3
R22100 VSS.n2945 VSS.n2944 9.3
R22101 VSS.n2946 VSS.n2945 9.3
R22102 VSS.n2952 VSS.n2951 9.3
R22103 VSS.n2955 VSS.n2954 9.3
R22104 VSS.n2955 VSS.n2810 9.3
R22105 VSS.n2810 VSS.n2809 9.3
R22106 VSS.n2963 VSS.n2962 9.3
R22107 VSS.n2962 VSS.n2961 9.3
R22108 VSS.n2961 VSS.n2960 9.3
R22109 VSS.n2884 VSS.n2883 9.3
R22110 VSS.n2896 VSS.n2858 9.3
R22111 VSS.n2852 VSS.n2851 9.3
R22112 VSS.n2929 VSS.n2928 9.3
R22113 VSS.n2941 VSS.n2820 9.3
R22114 VSS.n2814 VSS.n2813 9.3
R22115 VSS.n2800 VSS.n1313 9.3
R22116 VSS.n2797 VSS.n1314 9.3
R22117 VSS.n2797 VSS.n2796 9.3
R22118 VSS.n2796 VSS.n2795 9.3
R22119 VSS.n2790 VSS.n2789 9.3
R22120 VSS.n2787 VSS.n2786 9.3
R22121 VSS.n2786 VSS.n1318 9.3
R22122 VSS.n1318 VSS.n1317 9.3
R22123 VSS.n1326 VSS.n1320 9.3
R22124 VSS.n2779 VSS.n2778 9.3
R22125 VSS.n2780 VSS.n2779 9.3
R22126 VSS.n2781 VSS.n2780 9.3
R22127 VSS.n2776 VSS.n2775 9.3
R22128 VSS.n2767 VSS.n2766 9.3
R22129 VSS.n2767 VSS.n1330 9.3
R22130 VSS.n2771 VSS.n1330 9.3
R22131 VSS.n2765 VSS.n2764 9.3
R22132 VSS.n2762 VSS.n1336 9.3
R22133 VSS.n2762 VSS.n2761 9.3
R22134 VSS.n2761 VSS.n2760 9.3
R22135 VSS.n2755 VSS.n2754 9.3
R22136 VSS.n2752 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector 9.3
R22137 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector VSS.n1339 9.3
R22138 VSS.n1339 VSS.n1338 9.3
R22139 VSS.n1347 VSS.n1341 9.3
R22140 VSS.n2745 VSS.n2744 9.3
R22141 VSS.n2746 VSS.n2745 9.3
R22142 VSS.n2747 VSS.n2746 9.3
R22143 VSS.n2742 VSS.n2741 9.3
R22144 VSS.n2733 VSS.n2732 9.3
R22145 VSS.n2733 VSS.n1351 9.3
R22146 VSS.n2737 VSS.n1351 9.3
R22147 VSS.n2731 VSS.n2730 9.3
R22148 VSS.n2728 VSS.n1357 9.3
R22149 VSS.n2728 VSS.n2727 9.3
R22150 VSS.n2727 VSS.n2726 9.3
R22151 VSS.n2721 VSS.n2720 9.3
R22152 VSS.n2718 VSS.n2717 9.3
R22153 VSS.n2717 VSS.n1360 9.3
R22154 VSS.n1360 VSS.n1359 9.3
R22155 VSS.n1368 VSS.n1362 9.3
R22156 VSS.n2710 VSS.n2709 9.3
R22157 VSS.n2711 VSS.n2710 9.3
R22158 VSS.n2712 VSS.n2711 9.3
R22159 VSS.n2707 VSS.n2706 9.3
R22160 VSS.n2698 VSS.n2697 9.3
R22161 VSS.n2698 VSS.n1372 9.3
R22162 VSS.n2702 VSS.n1372 9.3
R22163 VSS.n2694 VSS.n1376 9.3
R22164 VSS.n2691 VSS.n1378 9.3
R22165 VSS.n2683 VSS.n1378 9.3
R22166 VSS.n2684 VSS.n2683 9.3
R22167 VSS.n2690 VSS.n2689 9.3
R22168 VSS.n2395 VSS.n2394 9.3
R22169 VSS.n2395 VSS.n1382 9.3
R22170 VSS.n1384 VSS.n1382 9.3
R22171 VSS.n2393 VSS.n2392 9.3
R22172 VSS.n2403 VSS.n2402 9.3
R22173 VSS.n2402 VSS.n2401 9.3
R22174 VSS.n2401 VSS.n2400 9.3
R22175 VSS.n2404 VSS.n2383 9.3
R22176 VSS.n2407 VSS.n2378 9.3
R22177 VSS.n2408 VSS.n2407 9.3
R22178 VSS.n2409 VSS.n2408 9.3
R22179 VSS.n2415 VSS.n2414 9.3
R22180 VSS.n2418 VSS.n2417 9.3
R22181 VSS.n2418 VSS.n2373 9.3
R22182 VSS.n2373 VSS.n2372 9.3
R22183 VSS.n2377 VSS.n2376 9.3
R22184 VSS.n2425 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector 9.3
R22185 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector VSS.n2424 9.3
R22186 VSS.n2424 VSS.n2423 9.3
R22187 VSS.n2426 VSS.n2364 9.3
R22188 VSS.n2429 VSS.n2359 9.3
R22189 VSS.n2430 VSS.n2429 9.3
R22190 VSS.n2431 VSS.n2430 9.3
R22191 VSS.n2437 VSS.n2436 9.3
R22192 VSS.n2440 VSS.n2439 9.3
R22193 VSS.n2440 VSS.n2354 9.3
R22194 VSS.n2354 VSS.n2353 9.3
R22195 VSS.n2358 VSS.n2357 9.3
R22196 VSS.n2448 VSS.n2447 9.3
R22197 VSS.n2447 VSS.n2446 9.3
R22198 VSS.n2446 VSS.n2445 9.3
R22199 VSS.n2449 VSS.n2345 9.3
R22200 VSS.n2452 VSS.n2340 9.3
R22201 VSS.n2453 VSS.n2452 9.3
R22202 VSS.n2454 VSS.n2453 9.3
R22203 VSS.n2460 VSS.n2459 9.3
R22204 VSS.n2463 VSS.n2462 9.3
R22205 VSS.n2463 VSS.n2335 9.3
R22206 VSS.n2335 VSS.n2334 9.3
R22207 VSS.n2339 VSS.n2338 9.3
R22208 VSS.n2471 VSS.n2470 9.3
R22209 VSS.n2470 VSS.n2469 9.3
R22210 VSS.n2469 VSS.n2468 9.3
R22211 VSS.n2473 VSS.n2290 9.3
R22212 VSS.n2476 VSS.n2285 9.3
R22213 VSS.n2477 VSS.n2476 9.3
R22214 VSS.n2478 VSS.n2477 9.3
R22215 VSS.n2484 VSS.n2483 9.3
R22216 VSS.n2487 VSS.n2486 9.3
R22217 VSS.n2487 VSS.n2280 9.3
R22218 VSS.n2280 VSS.n2279 9.3
R22219 VSS.n2284 VSS.n2283 9.3
R22220 VSS.n2495 VSS.n2494 9.3
R22221 VSS.n2494 VSS.n2493 9.3
R22222 VSS.n2493 VSS.n2492 9.3
R22223 VSS.n2496 VSS.n2271 9.3
R22224 VSS.n2499 VSS.n2266 9.3
R22225 VSS.n2500 VSS.n2499 9.3
R22226 VSS.n2501 VSS.n2500 9.3
R22227 VSS.n2507 VSS.n2506 9.3
R22228 VSS.n2510 VSS.n2509 9.3
R22229 VSS.n2510 VSS.n2261 9.3
R22230 VSS.n2261 VSS.n2260 9.3
R22231 VSS.n2265 VSS.n2264 9.3
R22232 VSS.n2517 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector 9.3
R22233 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector VSS.n2516 9.3
R22234 VSS.n2516 VSS.n2515 9.3
R22235 VSS.n2518 VSS.n2252 9.3
R22236 VSS.n2521 VSS.n2247 9.3
R22237 VSS.n2522 VSS.n2521 9.3
R22238 VSS.n2523 VSS.n2522 9.3
R22239 VSS.n2529 VSS.n2528 9.3
R22240 VSS.n2532 VSS.n2531 9.3
R22241 VSS.n2532 VSS.n2242 9.3
R22242 VSS.n2242 VSS.n2241 9.3
R22243 VSS.n2246 VSS.n2245 9.3
R22244 VSS.n2540 VSS.n2539 9.3
R22245 VSS.n2539 VSS.n2538 9.3
R22246 VSS.n2538 VSS.n2537 9.3
R22247 VSS.n2541 VSS.n2233 9.3
R22248 VSS.n2544 VSS.n2228 9.3
R22249 VSS.n2545 VSS.n2544 9.3
R22250 VSS.n2546 VSS.n2545 9.3
R22251 VSS.n2552 VSS.n2551 9.3
R22252 VSS.n2555 VSS.n2554 9.3
R22253 VSS.n2555 VSS.n2223 9.3
R22254 VSS.n2223 VSS.n2222 9.3
R22255 VSS.n2227 VSS.n2226 9.3
R22256 VSS.n2563 VSS.n2562 9.3
R22257 VSS.n2562 VSS.n2561 9.3
R22258 VSS.n2561 VSS.n2560 9.3
R22259 VSS.n2566 VSS.n2565 9.3
R22260 VSS.n2569 VSS.n2568 9.3
R22261 VSS.n2570 VSS.n2569 9.3
R22262 VSS.n2571 VSS.n2570 9.3
R22263 VSS.n2213 VSS.n2212 9.3
R22264 VSS.n2204 VSS.n2203 9.3
R22265 VSS.n2204 VSS.n1486 9.3
R22266 VSS.n2208 VSS.n1486 9.3
R22267 VSS.n2202 VSS.n2201 9.3
R22268 VSS.n2199 VSS.n1492 9.3
R22269 VSS.n2199 VSS.n2198 9.3
R22270 VSS.n2198 VSS.n2197 9.3
R22271 VSS.n2192 VSS.n2191 9.3
R22272 VSS.n2189 VSS.n2188 9.3
R22273 VSS.n2188 VSS.n1495 9.3
R22274 VSS.n1495 VSS.n1494 9.3
R22275 VSS.n1503 VSS.n1497 9.3
R22276 VSS.n2181 VSS.n2180 9.3
R22277 VSS.n2182 VSS.n2181 9.3
R22278 VSS.n2183 VSS.n2182 9.3
R22279 VSS.n2178 VSS.n2177 9.3
R22280 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector VSS.n2169 9.3
R22281 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector VSS.n1507 9.3
R22282 VSS.n2173 VSS.n1507 9.3
R22283 VSS.n2168 VSS.n2167 9.3
R22284 VSS.n2165 VSS.n1513 9.3
R22285 VSS.n2165 VSS.n2164 9.3
R22286 VSS.n2164 VSS.n2163 9.3
R22287 VSS.n2158 VSS.n2157 9.3
R22288 VSS.n2155 VSS.n2154 9.3
R22289 VSS.n2154 VSS.n1516 9.3
R22290 VSS.n1516 VSS.n1515 9.3
R22291 VSS.n1524 VSS.n1518 9.3
R22292 VSS.n2147 VSS.n2146 9.3
R22293 VSS.n2148 VSS.n2147 9.3
R22294 VSS.n2149 VSS.n2148 9.3
R22295 VSS.n2144 VSS.n2143 9.3
R22296 VSS.n2135 VSS.n2134 9.3
R22297 VSS.n2135 VSS.n1528 9.3
R22298 VSS.n2139 VSS.n1528 9.3
R22299 VSS.n2133 VSS.n2132 9.3
R22300 VSS.n2130 VSS.n1534 9.3
R22301 VSS.n2130 VSS.n2129 9.3
R22302 VSS.n2129 VSS.n2128 9.3
R22303 VSS.n2123 VSS.n2122 9.3
R22304 VSS.n2120 VSS.n2119 9.3
R22305 VSS.n2119 VSS.n1537 9.3
R22306 VSS.n1537 VSS.n1536 9.3
R22307 VSS.n2108 VSS.n2107 9.3
R22308 VSS.n2111 VSS.n2110 9.3
R22309 VSS.n2112 VSS.n2111 9.3
R22310 VSS.n2113 VSS.n2112 9.3
R22311 VSS.n1788 VSS.n1548 9.3
R22312 VSS.n1794 VSS.n1793 9.3
R22313 VSS.n1794 VSS.n1783 9.3
R22314 VSS.n1783 VSS.n1782 9.3
R22315 VSS.n1791 VSS.n1790 9.3
R22316 VSS.n1802 VSS.n1801 9.3
R22317 VSS.n1801 VSS.n1800 9.3
R22318 VSS.n1800 VSS.n1799 9.3
R22319 VSS.n1803 VSS.n1774 9.3
R22320 VSS.n1806 VSS.n1769 9.3
R22321 VSS.n1807 VSS.n1806 9.3
R22322 VSS.n1808 VSS.n1807 9.3
R22323 VSS.n1814 VSS.n1813 9.3
R22324 VSS.n1817 VSS.n1816 9.3
R22325 VSS.n1817 VSS.n1764 9.3
R22326 VSS.n1764 VSS.n1763 9.3
R22327 VSS.n1768 VSS.n1767 9.3
R22328 VSS.n1824 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector 9.3
R22329 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector VSS.n1823 9.3
R22330 VSS.n1823 VSS.n1822 9.3
R22331 VSS.n1825 VSS.n1755 9.3
R22332 VSS.n1828 VSS.n1750 9.3
R22333 VSS.n1829 VSS.n1828 9.3
R22334 VSS.n1830 VSS.n1829 9.3
R22335 VSS.n1836 VSS.n1835 9.3
R22336 VSS.n1839 VSS.n1838 9.3
R22337 VSS.n1839 VSS.n1745 9.3
R22338 VSS.n1745 VSS.n1744 9.3
R22339 VSS.n1749 VSS.n1748 9.3
R22340 VSS.n1847 VSS.n1846 9.3
R22341 VSS.n1846 VSS.n1845 9.3
R22342 VSS.n1845 VSS.n1844 9.3
R22343 VSS.n1848 VSS.n1736 9.3
R22344 VSS.n1851 VSS.n1731 9.3
R22345 VSS.n1852 VSS.n1851 9.3
R22346 VSS.n1853 VSS.n1852 9.3
R22347 VSS.n1859 VSS.n1858 9.3
R22348 VSS.n1862 VSS.n1861 9.3
R22349 VSS.n1862 VSS.n1726 9.3
R22350 VSS.n1726 VSS.n1725 9.3
R22351 VSS.n1730 VSS.n1729 9.3
R22352 VSS.n1870 VSS.n1869 9.3
R22353 VSS.n1869 VSS.n1868 9.3
R22354 VSS.n1868 VSS.n1867 9.3
R22355 VSS.n1872 VSS.n1681 9.3
R22356 VSS.n1875 VSS.n1676 9.3
R22357 VSS.n1876 VSS.n1875 9.3
R22358 VSS.n1877 VSS.n1876 9.3
R22359 VSS.n1883 VSS.n1882 9.3
R22360 VSS.n1886 VSS.n1885 9.3
R22361 VSS.n1886 VSS.n1671 9.3
R22362 VSS.n1671 VSS.n1670 9.3
R22363 VSS.n1675 VSS.n1674 9.3
R22364 VSS.n1894 VSS.n1893 9.3
R22365 VSS.n1893 VSS.n1892 9.3
R22366 VSS.n1892 VSS.n1891 9.3
R22367 VSS.n1895 VSS.n1662 9.3
R22368 VSS.n1898 VSS.n1657 9.3
R22369 VSS.n1899 VSS.n1898 9.3
R22370 VSS.n1900 VSS.n1899 9.3
R22371 VSS.n1906 VSS.n1905 9.3
R22372 VSS.n1909 VSS.n1908 9.3
R22373 VSS.n1909 VSS.n1652 9.3
R22374 VSS.n1652 VSS.n1651 9.3
R22375 VSS.n1656 VSS.n1655 9.3
R22376 VSS.n1916 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector 9.3
R22377 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector VSS.n1915 9.3
R22378 VSS.n1915 VSS.n1914 9.3
R22379 VSS.n1917 VSS.n1643 9.3
R22380 VSS.n1920 VSS.n1638 9.3
R22381 VSS.n1921 VSS.n1920 9.3
R22382 VSS.n1922 VSS.n1921 9.3
R22383 VSS.n1928 VSS.n1927 9.3
R22384 VSS.n1931 VSS.n1930 9.3
R22385 VSS.n1931 VSS.n1633 9.3
R22386 VSS.n1633 VSS.n1632 9.3
R22387 VSS.n1637 VSS.n1636 9.3
R22388 VSS.n1939 VSS.n1938 9.3
R22389 VSS.n1938 VSS.n1937 9.3
R22390 VSS.n1937 VSS.n1936 9.3
R22391 VSS.n1940 VSS.n1624 9.3
R22392 VSS.n1943 VSS.n1619 9.3
R22393 VSS.n1944 VSS.n1943 9.3
R22394 VSS.n1945 VSS.n1944 9.3
R22395 VSS.n1951 VSS.n1950 9.3
R22396 VSS.n1954 VSS.n1953 9.3
R22397 VSS.n1954 VSS.n1613 9.3
R22398 VSS.n1613 VSS.n1612 9.3
R22399 VSS.n1618 VSS.n1617 9.3
R22400 VSS.n1961 VSS.n1610 9.3
R22401 VSS.n1961 VSS.n1960 9.3
R22402 VSS.n1960 VSS.n1959 9.3
R22403 VSS.n2876 VSS.n2872 9.3
R22404 VSS.n2876 VSS.n1270 9.3
R22405 VSS.n1272 VSS.n1270 9.3
R22406 VSS.n2873 VSS.n1269 9.3
R22407 VSS.n674 VSS.n673 9.3
R22408 VSS.n673 VSS.n573 9.3
R22409 VSS.n676 VSS.n675 9.3
R22410 VSS.n680 VSS.n679 9.3
R22411 VSS.n679 VSS.n678 9.3
R22412 VSS.n686 VSS.n685 9.3
R22413 VSS.n685 VSS.n684 9.3
R22414 VSS.n688 VSS.n687 9.3
R22415 VSS.n692 VSS.n691 9.3
R22416 VSS.n691 VSS.n690 9.3
R22417 VSS.n698 VSS.n697 9.3
R22418 VSS.n697 VSS.n696 9.3
R22419 VSS.n699 VSS.n644 9.3
R22420 VSS.n703 VSS.n643 9.3
R22421 VSS.n703 VSS.n702 9.3
R22422 VSS.n712 VSS.n710 9.3
R22423 VSS.n712 VSS.n711 9.3
R22424 VSS.n642 VSS.n584 9.3
R22425 VSS.n639 VSS.n586 9.3
R22426 VSS.n639 VSS.n583 9.3
R22427 VSS.n671 VSS.n670 9.3
R22428 VSS.n682 VSS.n681 9.3
R22429 VSS.n694 VSS.n693 9.3
R22430 VSS.n708 VSS.n707 9.3
R22431 VSS.n669 VSS.n668 9.3
R22432 VSS.n668 VSS.n548 9.3
R22433 VSS.n546 VSS.n545 9.3
R22434 VSS.n764 VSS.n763 9.3
R22435 VSS.n763 VSS.n483 9.3
R22436 VSS.n766 VSS.n765 9.3
R22437 VSS.n770 VSS.n769 9.3
R22438 VSS.n769 VSS.n768 9.3
R22439 VSS.n776 VSS.n775 9.3
R22440 VSS.n775 VSS.n774 9.3
R22441 VSS.n778 VSS.n777 9.3
R22442 VSS.n782 VSS.n781 9.3
R22443 VSS.n781 VSS.n780 9.3
R22444 VSS.n788 VSS.n787 9.3
R22445 VSS.n787 VSS.n786 9.3
R22446 VSS.n789 VSS.n734 9.3
R22447 VSS.n793 VSS.n733 9.3
R22448 VSS.n793 VSS.n792 9.3
R22449 VSS.n802 VSS.n800 9.3
R22450 VSS.n802 VSS.n801 9.3
R22451 VSS.n732 VSS.n494 9.3
R22452 VSS.n729 VSS.n496 9.3
R22453 VSS.n729 VSS.n493 9.3
R22454 VSS.n761 VSS.n760 9.3
R22455 VSS.n772 VSS.n771 9.3
R22456 VSS.n784 VSS.n783 9.3
R22457 VSS.n798 VSS.n797 9.3
R22458 VSS.n759 VSS.n758 9.3
R22459 VSS.n758 VSS.n458 9.3
R22460 VSS.n456 VSS.n455 9.3
R22461 VSS.n854 VSS.n853 9.3
R22462 VSS.n853 VSS.n393 9.3
R22463 VSS.n856 VSS.n855 9.3
R22464 VSS.n860 VSS.n859 9.3
R22465 VSS.n859 VSS.n858 9.3
R22466 VSS.n866 VSS.n865 9.3
R22467 VSS.n865 VSS.n864 9.3
R22468 VSS.n868 VSS.n867 9.3
R22469 VSS.n872 VSS.n871 9.3
R22470 VSS.n871 VSS.n870 9.3
R22471 VSS.n878 VSS.n877 9.3
R22472 VSS.n877 VSS.n876 9.3
R22473 VSS.n879 VSS.n824 9.3
R22474 VSS.n883 VSS.n823 9.3
R22475 VSS.n883 VSS.n882 9.3
R22476 VSS.n892 VSS.n890 9.3
R22477 VSS.n892 VSS.n891 9.3
R22478 VSS.n822 VSS.n404 9.3
R22479 VSS.n819 VSS.n406 9.3
R22480 VSS.n819 VSS.n403 9.3
R22481 VSS.n851 VSS.n850 9.3
R22482 VSS.n862 VSS.n861 9.3
R22483 VSS.n874 VSS.n873 9.3
R22484 VSS.n888 VSS.n887 9.3
R22485 VSS.n849 VSS.n848 9.3
R22486 VSS.n848 VSS.n368 9.3
R22487 VSS.n366 VSS.n365 9.3
R22488 VSS.n944 VSS.n943 9.3
R22489 VSS.n943 VSS.n303 9.3
R22490 VSS.n946 VSS.n945 9.3
R22491 VSS.n950 VSS.n949 9.3
R22492 VSS.n949 VSS.n948 9.3
R22493 VSS.n956 VSS.n955 9.3
R22494 VSS.n955 VSS.n954 9.3
R22495 VSS.n958 VSS.n957 9.3
R22496 VSS.n962 VSS.n961 9.3
R22497 VSS.n961 VSS.n960 9.3
R22498 VSS.n968 VSS.n967 9.3
R22499 VSS.n967 VSS.n966 9.3
R22500 VSS.n969 VSS.n914 9.3
R22501 VSS.n973 VSS.n913 9.3
R22502 VSS.n973 VSS.n972 9.3
R22503 VSS.n982 VSS.n980 9.3
R22504 VSS.n982 VSS.n981 9.3
R22505 VSS.n912 VSS.n314 9.3
R22506 VSS.n909 VSS.n316 9.3
R22507 VSS.n909 VSS.n313 9.3
R22508 VSS.n941 VSS.n940 9.3
R22509 VSS.n952 VSS.n951 9.3
R22510 VSS.n964 VSS.n963 9.3
R22511 VSS.n978 VSS.n977 9.3
R22512 VSS.n939 VSS.n938 9.3
R22513 VSS.n938 VSS.n278 9.3
R22514 VSS.n276 VSS.n275 9.3
R22515 VSS.n1034 VSS.n1033 9.3
R22516 VSS.n1033 VSS.n213 9.3
R22517 VSS.n1036 VSS.n1035 9.3
R22518 VSS.n1040 VSS.n1039 9.3
R22519 VSS.n1039 VSS.n1038 9.3
R22520 VSS.n1046 VSS.n1045 9.3
R22521 VSS.n1045 VSS.n1044 9.3
R22522 VSS.n1048 VSS.n1047 9.3
R22523 VSS.n1052 VSS.n1051 9.3
R22524 VSS.n1051 VSS.n1050 9.3
R22525 VSS.n1058 VSS.n1057 9.3
R22526 VSS.n1057 VSS.n1056 9.3
R22527 VSS.n1059 VSS.n1004 9.3
R22528 VSS.n1063 VSS.n1003 9.3
R22529 VSS.n1063 VSS.n1062 9.3
R22530 VSS.n1072 VSS.n1070 9.3
R22531 VSS.n1072 VSS.n1071 9.3
R22532 VSS.n1002 VSS.n224 9.3
R22533 VSS.n999 VSS.n226 9.3
R22534 VSS.n999 VSS.n223 9.3
R22535 VSS.n1031 VSS.n1030 9.3
R22536 VSS.n1042 VSS.n1041 9.3
R22537 VSS.n1054 VSS.n1053 9.3
R22538 VSS.n1068 VSS.n1067 9.3
R22539 VSS.n1029 VSS.n1028 9.3
R22540 VSS.n1028 VSS.n188 9.3
R22541 VSS.n186 VSS.n185 9.3
R22542 VSS.n1124 VSS.n1123 9.3
R22543 VSS.n1123 VSS.n123 9.3
R22544 VSS.n1126 VSS.n1125 9.3
R22545 VSS.n1130 VSS.n1129 9.3
R22546 VSS.n1129 VSS.n1128 9.3
R22547 VSS.n1136 VSS.n1135 9.3
R22548 VSS.n1135 VSS.n1134 9.3
R22549 VSS.n1138 VSS.n1137 9.3
R22550 VSS.n1142 VSS.n1141 9.3
R22551 VSS.n1141 VSS.n1140 9.3
R22552 VSS.n1148 VSS.n1147 9.3
R22553 VSS.n1147 VSS.n1146 9.3
R22554 VSS.n1149 VSS.n1094 9.3
R22555 VSS.n1153 VSS.n1093 9.3
R22556 VSS.n1153 VSS.n1152 9.3
R22557 VSS.n1162 VSS.n1160 9.3
R22558 VSS.n1162 VSS.n1161 9.3
R22559 VSS.n1092 VSS.n134 9.3
R22560 VSS.n1089 VSS.n136 9.3
R22561 VSS.n1089 VSS.n133 9.3
R22562 VSS.n1121 VSS.n1120 9.3
R22563 VSS.n1132 VSS.n1131 9.3
R22564 VSS.n1144 VSS.n1143 9.3
R22565 VSS.n1158 VSS.n1157 9.3
R22566 VSS.n1119 VSS.n1118 9.3
R22567 VSS.n1118 VSS.n98 9.3
R22568 VSS.n96 VSS.n95 9.3
R22569 VSS.n1209 VSS.n1208 9.3
R22570 VSS.n1208 VSS.n32 9.3
R22571 VSS.n1211 VSS.n1210 9.3
R22572 VSS.n1215 VSS.n1214 9.3
R22573 VSS.n1214 VSS.n1213 9.3
R22574 VSS.n1221 VSS.n1220 9.3
R22575 VSS.n1220 VSS.n1219 9.3
R22576 VSS.n1223 VSS.n1222 9.3
R22577 VSS.n1227 VSS.n1226 9.3
R22578 VSS.n1226 VSS.n1225 9.3
R22579 VSS.n1233 VSS.n1232 9.3
R22580 VSS.n1232 VSS.n1231 9.3
R22581 VSS.n1234 VSS.n1184 9.3
R22582 VSS.n1238 VSS.n1183 9.3
R22583 VSS.n1238 VSS.n1237 9.3
R22584 VSS.n1247 VSS.n1245 9.3
R22585 VSS.n1247 VSS.n1246 9.3
R22586 VSS.n1182 VSS.n43 9.3
R22587 VSS.n1179 VSS.n45 9.3
R22588 VSS.n1179 VSS.n42 9.3
R22589 VSS.n1206 VSS.n1205 9.3
R22590 VSS.n1217 VSS.n1216 9.3
R22591 VSS.n1229 VSS.n1228 9.3
R22592 VSS.n1243 VSS.n1242 9.3
R22593 VSS.n1256 VSS.n5 9.3
R22594 VSS.n1256 VSS.n1255 9.3
R22595 VSS.n1259 VSS.n4 9.3
R22596 VSS.n1261 VSS.n1260 9.3
R22597 VSS.n17663 VSS.n17662 9.3
R22598 VSS.n17666 VSS.n17654 9.3
R22599 VSS.n17671 VSS.n17652 9.3
R22600 VSS.n17677 VSS.n17676 9.3
R22601 VSS.n17684 VSS.n17683 9.3
R22602 VSS.n17689 VSS.n17646 9.3
R22603 VSS.n17694 VSS.n17644 9.3
R22604 VSS.n17700 VSS.n17699 9.3
R22605 VSS.n17701 VSS.n17641 9.3
R22606 VSS.n17698 VSS.n17643 9.3
R22607 VSS.n17697 VSS.n17696 9.3
R22608 VSS.n17693 VSS.n17645 9.3
R22609 VSS.n17691 VSS.n17690 9.3
R22610 VSS.n17688 VSS.n17687 9.3
R22611 VSS.n17685 VSS.n17647 9.3
R22612 VSS.n17682 VSS.n17648 9.3
R22613 VSS.n17678 VSS.n17649 9.3
R22614 VSS.n17675 VSS.n17651 9.3
R22615 VSS.n17674 VSS.n17673 9.3
R22616 VSS.n17670 VSS.n17669 9.3
R22617 VSS.n17668 VSS.n17667 9.3
R22618 VSS.n17665 VSS.n17664 9.3
R22619 VSS.n17661 VSS.n17656 9.3
R22620 VSS.n17660 VSS.n17659 9.3
R22621 VSS.n17329 VSS.n17328 9.066
R22622 VSS.n17223 VSS.n17222 9.066
R22623 VSS.n17133 VSS.n17132 9.066
R22624 VSS.n17043 VSS.n17042 9.066
R22625 VSS.n16953 VSS.n16952 9.066
R22626 VSS.n16863 VSS.n16862 9.066
R22627 VSS.n16773 VSS.n16772 9.066
R22628 VSS.n16683 VSS.n16682 9.066
R22629 VSS.n11151 VSS.n11149 9.066
R22630 VSS.n11241 VSS.n11239 9.066
R22631 VSS.n11331 VSS.n11329 9.066
R22632 VSS.n11421 VSS.n11419 9.066
R22633 VSS.n13541 VSS.n13539 9.066
R22634 VSS.n13631 VSS.n13629 9.066
R22635 VSS.n13721 VSS.n13719 9.066
R22636 VSS.n13826 VSS.n13825 9.066
R22637 VSS.n9159 VSS.n9158 9.066
R22638 VSS.n10178 VSS.n10177 9.066
R22639 VSS.n10088 VSS.n10087 9.066
R22640 VSS.n9998 VSS.n9997 9.066
R22641 VSS.n9908 VSS.n9907 9.066
R22642 VSS.n9818 VSS.n9817 9.066
R22643 VSS.n9728 VSS.n9727 9.066
R22644 VSS.n10317 VSS.n9181 9.066
R22645 VSS.n5668 VSS.n3577 9.066
R22646 VSS.n5790 VSS.n3519 9.066
R22647 VSS.n5912 VSS.n3461 9.066
R22648 VSS.n6034 VSS.n3403 9.066
R22649 VSS.n6156 VSS.n3345 9.066
R22650 VSS.n6278 VSS.n3287 9.066
R22651 VSS.n6400 VSS.n3229 9.066
R22652 VSS.n6538 VSS.n6537 9.066
R22653 VSS.n1176 VSS.n1175 9.066
R22654 VSS.n1086 VSS.n1085 9.066
R22655 VSS.n996 VSS.n995 9.066
R22656 VSS.n906 VSS.n905 9.066
R22657 VSS.n816 VSS.n815 9.066
R22658 VSS.n726 VSS.n725 9.066
R22659 VSS.n636 VSS.n635 9.066
R22660 VSS.n14014 VSS.n14013 8.921
R22661 VSS.n12063 VSS.n12062 8.921
R22662 VSS.n7175 VSS.n7005 8.921
R22663 VSS.n3645 VSS.n3644 8.921
R22664 VSS.n3044 VSS.n1269 8.921
R22665 VSS.n6801 VSS.n6800 8.791
R22666 VSS.n17551 sky130_asc_res_xhigh_po_2p85_1_15/VGND 8.691
R22667 VSS.n6880 VSS.n6729 8.662
R22668 VSS.n17526 sky130_asc_res_xhigh_po_2p85_1_12/VGND 8.593
R22669 VSS.n14728 VSS.n14362 8.533
R22670 VSS.n15998 VSS.n15997 8.533
R22671 VSS.n12791 VSS.n12789 8.533
R22672 VSS.n12213 VSS.n12212 8.533
R22673 VSS.n7842 VSS.n7841 8.533
R22674 VSS.n7179 VSS.n7178 8.533
R22675 VSS.n6831 VSS.n6756 8.533
R22676 VSS.n4244 VSS.n4242 8.533
R22677 VSS.n5655 VSS.n3648 8.533
R22678 VSS.n1969 VSS.n1603 8.533
R22679 VSS.n3045 VSS.n1268 8.533
R22680 VSS sky130_asc_cap_mim_m3_1_4/VGND 8.443
R22681 VSS.n6880 VSS.n6879 8.403
R22682 VSS.n16765 VSS.n16764 8.156
R22683 VSS.n16855 VSS.n16854 8.156
R22684 VSS.n16945 VSS.n16944 8.156
R22685 VSS.n17035 VSS.n17034 8.156
R22686 VSS.n17125 VSS.n17124 8.156
R22687 VSS.n17215 VSS.n17214 8.156
R22688 VSS.n17305 VSS.n17304 8.156
R22689 VSS.n9810 VSS.n9809 8.156
R22690 VSS.n9900 VSS.n9899 8.156
R22691 VSS.n9990 VSS.n9989 8.156
R22692 VSS.n10080 VSS.n10079 8.156
R22693 VSS.n10170 VSS.n10169 8.156
R22694 VSS.n10260 VSS.n10259 8.156
R22695 VSS.n8977 VSS.n8935 8.156
R22696 VSS.n6598 VSS.n6597 8.156
R22697 VSS.n3282 VSS.n3234 8.156
R22698 VSS.n3340 VSS.n3292 8.156
R22699 VSS.n3398 VSS.n3350 8.156
R22700 VSS.n3456 VSS.n3408 8.156
R22701 VSS.n3514 VSS.n3466 8.156
R22702 VSS.n3572 VSS.n3524 8.156
R22703 VSS.n3630 VSS.n3582 8.156
R22704 VSS.n718 VSS.n717 8.156
R22705 VSS.n808 VSS.n807 8.156
R22706 VSS.n898 VSS.n897 8.156
R22707 VSS.n988 VSS.n987 8.156
R22708 VSS.n1078 VSS.n1077 8.156
R22709 VSS.n1168 VSS.n1167 8.156
R22710 VSS.n1252 VSS.n7 8.156
R22711 VSS.n10463 VSS.n10462 8.153
R22712 VSS.n17650 VSS.n17642 8.152
R22713 VSS.n14722 VSS.n14367 8.145
R22714 VSS.n12793 VSS.n12792 8.145
R22715 VSS.n7836 VSS.n7671 8.145
R22716 VSS.n4246 VSS.n4245 8.145
R22717 VSS.n1963 VSS.n1608 8.145
R22718 VSS.n10462 VSS.n10429 8.125
R22719 VSS.n10462 VSS.n10424 8.125
R22720 VSS.n17672 VSS.n17642 8.125
R22721 VSS.n17686 VSS.n17642 8.124
R22722 VSS.n10462 VSS.n10430 8.097
R22723 VSS.n10462 VSS.n10422 8.097
R22724 VSS.n17653 VSS.n17642 8.097
R22725 VSS.n17692 VSS.n17642 8.096
R22726 VSS.n10462 VSS.n10431 8.069
R22727 VSS.n10462 VSS.n10420 8.069
R22728 VSS.n17655 VSS.n17642 8.069
R22729 VSS.n17695 VSS.n17642 8.069
R22730 VSS.n6606 VSS.n6605 8.069
R22731 VSS.n10462 VSS.n10461 8.043
R22732 VSS.n10462 VSS.n10418 8.043
R22733 VSS.n17702 VSS.n17642 8.043
R22734 VSS.n17657 VSS.n17642 8.043
R22735 sky130_asc_cap_mim_m3_1_0/VGND sky130_asc_nfet_01v8_lvt_1_1/VGND 7.799
R22736 sky130_asc_nfet_01v8_lvt_9_1/VGND VSS.n3135 7.749
R22737 sky130_asc_cap_mim_m3_1_3/VGND sky130_asc_cap_mim_m3_1_0/VGND 7.73
R22738 sky130_asc_cap_mim_m3_1_1/VGND sky130_asc_cap_mim_m3_1_3/VGND 7.73
R22739 sky130_asc_pfet_01v8_lvt_60_1/VGND sky130_asc_cap_mim_m3_1_2/VGND 7.728
R22740 VSS.n9157 VSS.n9156 7.464
R22741 VSS.t20 VSS.n9155 7.262
R22742 VSS.n15684 VSS.n15682 7.24
R22743 VSS.n15785 VSS.n15784 7.24
R22744 VSS.n15693 VSS.n15691 7.24
R22745 VSS.n15703 VSS.n15701 7.24
R22746 VSS.n15762 VSS.n15761 7.24
R22747 VSS.n15712 VSS.n15710 7.24
R22748 VSS.n15722 VSS.n15720 7.24
R22749 VSS.n15740 VSS.n15739 7.24
R22750 VSS.n15730 VSS.n15729 7.24
R22751 VSS.n14006 VSS.n14004 7.24
R22752 VSS.n16010 VSS.n16009 7.24
R22753 VSS.n15572 VSS.n15570 7.24
R22754 VSS.n15877 VSS.n15876 7.24
R22755 VSS.n15581 VSS.n15579 7.24
R22756 VSS.n15591 VSS.n15589 7.24
R22757 VSS.n15854 VSS.n15853 7.24
R22758 VSS.n15600 VSS.n15598 7.24
R22759 VSS.n15610 VSS.n15608 7.24
R22760 VSS.n15832 VSS.n15831 7.24
R22761 VSS.n15619 VSS.n15617 7.24
R22762 VSS.n15629 VSS.n15627 7.24
R22763 VSS.n15809 VSS.n15808 7.24
R22764 VSS.n15465 VSS.n15464 7.24
R22765 VSS.n14127 VSS.n14122 7.24
R22766 VSS.n15481 VSS.n15480 7.24
R22767 VSS.n15489 VSS.n14113 7.24
R22768 VSS.n15500 VSS.n15499 7.24
R22769 VSS.n14106 VSS.n14101 7.24
R22770 VSS.n15515 VSS.n15514 7.24
R22771 VSS.n15523 VSS.n14092 7.24
R22772 VSS.n15534 VSS.n15533 7.24
R22773 VSS.n14085 VSS.n14080 7.24
R22774 VSS.n15550 VSS.n15549 7.24
R22775 VSS.n15097 VSS.n15095 7.24
R22776 VSS.n15218 VSS.n15217 7.24
R22777 VSS.n15106 VSS.n15104 7.24
R22778 VSS.n15116 VSS.n15114 7.24
R22779 VSS.n15195 VSS.n15194 7.24
R22780 VSS.n15125 VSS.n15123 7.24
R22781 VSS.n15135 VSS.n15133 7.24
R22782 VSS.n15173 VSS.n15172 7.24
R22783 VSS.n15144 VSS.n15142 7.24
R22784 VSS.n15151 VSS.n15150 7.24
R22785 VSS.n15448 VSS.n15447 7.24
R22786 VSS.n14985 VSS.n14983 7.24
R22787 VSS.n15310 VSS.n15309 7.24
R22788 VSS.n14994 VSS.n14992 7.24
R22789 VSS.n15004 VSS.n15002 7.24
R22790 VSS.n15287 VSS.n15286 7.24
R22791 VSS.n15013 VSS.n15011 7.24
R22792 VSS.n15023 VSS.n15021 7.24
R22793 VSS.n15265 VSS.n15264 7.24
R22794 VSS.n15032 VSS.n15030 7.24
R22795 VSS.n15042 VSS.n15040 7.24
R22796 VSS.n15242 VSS.n15241 7.24
R22797 VSS.n14883 VSS.n14882 7.24
R22798 VSS.n14891 VSS.n14290 7.24
R22799 VSS.n14902 VSS.n14901 7.24
R22800 VSS.n14283 VSS.n14278 7.24
R22801 VSS.n14918 VSS.n14917 7.24
R22802 VSS.n14926 VSS.n14269 7.24
R22803 VSS.n14936 VSS.n14935 7.24
R22804 VSS.n14262 VSS.n14257 7.24
R22805 VSS.n14952 VSS.n14951 7.24
R22806 VSS.n14960 VSS.n14248 7.24
R22807 VSS.n14971 VSS.n14970 7.24
R22808 VSS.n14488 VSS.n14486 7.24
R22809 VSS.n14617 VSS.n14616 7.24
R22810 VSS.n14497 VSS.n14495 7.24
R22811 VSS.n14507 VSS.n14505 7.24
R22812 VSS.n14594 VSS.n14593 7.24
R22813 VSS.n14516 VSS.n14514 7.24
R22814 VSS.n14526 VSS.n14524 7.24
R22815 VSS.n14572 VSS.n14571 7.24
R22816 VSS.n14535 VSS.n14533 7.24
R22817 VSS.n14549 VSS.n14543 7.24
R22818 VSS.n14547 VSS.n14546 7.24
R22819 VSS.n14376 VSS.n14373 7.24
R22820 VSS.n14709 VSS.n14708 7.24
R22821 VSS.n14385 VSS.n14383 7.24
R22822 VSS.n14395 VSS.n14393 7.24
R22823 VSS.n14686 VSS.n14685 7.24
R22824 VSS.n14404 VSS.n14402 7.24
R22825 VSS.n14414 VSS.n14412 7.24
R22826 VSS.n14664 VSS.n14663 7.24
R22827 VSS.n14423 VSS.n14421 7.24
R22828 VSS.n14433 VSS.n14431 7.24
R22829 VSS.n14641 VSS.n14640 7.24
R22830 VSS.n11998 VSS.n11996 7.24
R22831 VSS.n12293 VSS.n12292 7.24
R22832 VSS.n12007 VSS.n12005 7.24
R22833 VSS.n12017 VSS.n12015 7.24
R22834 VSS.n12270 VSS.n12269 7.24
R22835 VSS.n12026 VSS.n12024 7.24
R22836 VSS.n12036 VSS.n12034 7.24
R22837 VSS.n12248 VSS.n12247 7.24
R22838 VSS.n12045 VSS.n12043 7.24
R22839 VSS.n12055 VSS.n12053 7.24
R22840 VSS.n12225 VSS.n12224 7.24
R22841 VSS.n11919 VSS.n11917 7.24
R22842 VSS.n12385 VSS.n12384 7.24
R22843 VSS.n11928 VSS.n11926 7.24
R22844 VSS.n11938 VSS.n11936 7.24
R22845 VSS.n12362 VSS.n12361 7.24
R22846 VSS.n11947 VSS.n11945 7.24
R22847 VSS.n11957 VSS.n11955 7.24
R22848 VSS.n12340 VSS.n12339 7.24
R22849 VSS.n11966 VSS.n11964 7.24
R22850 VSS.n11976 VSS.n11974 7.24
R22851 VSS.n12317 VSS.n12316 7.24
R22852 VSS.n11817 VSS.n11816 7.24
R22853 VSS.n11825 VSS.n11595 7.24
R22854 VSS.n11836 VSS.n11835 7.24
R22855 VSS.n11588 VSS.n11583 7.24
R22856 VSS.n11852 VSS.n11851 7.24
R22857 VSS.n11860 VSS.n11574 7.24
R22858 VSS.n11870 VSS.n11869 7.24
R22859 VSS.n11567 VSS.n11562 7.24
R22860 VSS.n11886 VSS.n11885 7.24
R22861 VSS.n11894 VSS.n11553 7.24
R22862 VSS.n11905 VSS.n11904 7.24
R22863 VSS.n11679 VSS.n11667 7.24
R22864 VSS.n11690 VSS.n11689 7.24
R22865 VSS.n11660 VSS.n11655 7.24
R22866 VSS.n11706 VSS.n11705 7.24
R22867 VSS.n11714 VSS.n11646 7.24
R22868 VSS.n11725 VSS.n11724 7.24
R22869 VSS.n11639 VSS.n11634 7.24
R22870 VSS.n11740 VSS.n11739 7.24
R22871 VSS.n11748 VSS.n11625 7.24
R22872 VSS.n11759 VSS.n11758 7.24
R22873 VSS.n11618 VSS.n11617 7.24
R22874 VSS.n13297 VSS.n13296 7.24
R22875 VSS.n13260 VSS.n13258 7.24
R22876 VSS.n13274 VSS.n13268 7.24
R22877 VSS.n13272 VSS.n13271 7.24
R22878 VSS.n11440 VSS.n11438 7.24
R22879 VSS.n13444 VSS.n13443 7.24
R22880 VSS.n11449 VSS.n11447 7.24
R22881 VSS.n11459 VSS.n11457 7.24
R22882 VSS.n13422 VSS.n13421 7.24
R22883 VSS.n11468 VSS.n11466 7.24
R22884 VSS.n11478 VSS.n11476 7.24
R22885 VSS.n13158 VSS.n12576 7.24
R22886 VSS.n13169 VSS.n13168 7.24
R22887 VSS.n12569 VSS.n12564 7.24
R22888 VSS.n13185 VSS.n13184 7.24
R22889 VSS.n13193 VSS.n12555 7.24
R22890 VSS.n13204 VSS.n13203 7.24
R22891 VSS.n12548 VSS.n12543 7.24
R22892 VSS.n13219 VSS.n13218 7.24
R22893 VSS.n13227 VSS.n12534 7.24
R22894 VSS.n13239 VSS.n13238 7.24
R22895 VSS.n13245 VSS.n13244 7.24
R22896 VSS.n13048 VSS.n13047 7.24
R22897 VSS.n12903 VSS.n12901 7.24
R22898 VSS.n12913 VSS.n12911 7.24
R22899 VSS.n13025 VSS.n13024 7.24
R22900 VSS.n12922 VSS.n12920 7.24
R22901 VSS.n12932 VSS.n12930 7.24
R22902 VSS.n13003 VSS.n13002 7.24
R22903 VSS.n12941 VSS.n12939 7.24
R22904 VSS.n12951 VSS.n12949 7.24
R22905 VSS.n12980 VSS.n12979 7.24
R22906 VSS.n12961 VSS.n12958 7.24
R22907 VSS.n12801 VSS.n12717 7.24
R22908 VSS.n12812 VSS.n12811 7.24
R22909 VSS.n12710 VSS.n12705 7.24
R22910 VSS.n12828 VSS.n12827 7.24
R22911 VSS.n12836 VSS.n12696 7.24
R22912 VSS.n12847 VSS.n12846 7.24
R22913 VSS.n12689 VSS.n12684 7.24
R22914 VSS.n12862 VSS.n12861 7.24
R22915 VSS.n12870 VSS.n12675 7.24
R22916 VSS.n12882 VSS.n12881 7.24
R22917 VSS.n12888 VSS.n12887 7.24
R22918 VSS.n7081 VSS.n7080 7.24
R22919 VSS.n7062 VSS.n7057 7.24
R22920 VSS.n7097 VSS.n7096 7.24
R22921 VSS.n7105 VSS.n7048 7.24
R22922 VSS.n7116 VSS.n7115 7.24
R22923 VSS.n7041 VSS.n7036 7.24
R22924 VSS.n7131 VSS.n7130 7.24
R22925 VSS.n7139 VSS.n7027 7.24
R22926 VSS.n7150 VSS.n7149 7.24
R22927 VSS.n7020 VSS.n7015 7.24
R22928 VSS.n7166 VSS.n7165 7.24
R22929 VSS.n8756 VSS.n8739 7.24
R22930 VSS.n8749 VSS.n8748 7.24
R22931 VSS.n6912 VSS.n6910 7.24
R22932 VSS.n8916 VSS.n8915 7.24
R22933 VSS.n6921 VSS.n6919 7.24
R22934 VSS.n6931 VSS.n6929 7.24
R22935 VSS.n8894 VSS.n8893 7.24
R22936 VSS.n6940 VSS.n6938 7.24
R22937 VSS.n6950 VSS.n6948 7.24
R22938 VSS.n8871 VSS.n8870 7.24
R22939 VSS.n6959 VSS.n6957 7.24
R22940 VSS.n8644 VSS.n8643 7.24
R22941 VSS.n8652 VSS.n7309 7.24
R22942 VSS.n8663 VSS.n8662 7.24
R22943 VSS.n7302 VSS.n7297 7.24
R22944 VSS.n8679 VSS.n8678 7.24
R22945 VSS.n8687 VSS.n7288 7.24
R22946 VSS.n8697 VSS.n8696 7.24
R22947 VSS.n7281 VSS.n7276 7.24
R22948 VSS.n8713 VSS.n8712 7.24
R22949 VSS.n8721 VSS.n7267 7.24
R22950 VSS.n8732 VSS.n8731 7.24
R22951 VSS.n8534 VSS.n8381 7.24
R22952 VSS.n8395 VSS.n8392 7.24
R22953 VSS.n8521 VSS.n8520 7.24
R22954 VSS.n8404 VSS.n8402 7.24
R22955 VSS.n8414 VSS.n8412 7.24
R22956 VSS.n8498 VSS.n8497 7.24
R22957 VSS.n8423 VSS.n8421 7.24
R22958 VSS.n8433 VSS.n8431 7.24
R22959 VSS.n8476 VSS.n8475 7.24
R22960 VSS.n8442 VSS.n8440 7.24
R22961 VSS.n8451 VSS.n8449 7.24
R22962 VSS.n8286 VSS.n8285 7.24
R22963 VSS.n8294 VSS.n7449 7.24
R22964 VSS.n8305 VSS.n8304 7.24
R22965 VSS.n7442 VSS.n7437 7.24
R22966 VSS.n8321 VSS.n8320 7.24
R22967 VSS.n8329 VSS.n7428 7.24
R22968 VSS.n8339 VSS.n8338 7.24
R22969 VSS.n7421 VSS.n7416 7.24
R22970 VSS.n8355 VSS.n8354 7.24
R22971 VSS.n8363 VSS.n7407 7.24
R22972 VSS.n8374 VSS.n8373 7.24
R22973 VSS.n8176 VSS.n8023 7.24
R22974 VSS.n8037 VSS.n8034 7.24
R22975 VSS.n8163 VSS.n8162 7.24
R22976 VSS.n8046 VSS.n8044 7.24
R22977 VSS.n8056 VSS.n8054 7.24
R22978 VSS.n8140 VSS.n8139 7.24
R22979 VSS.n8065 VSS.n8063 7.24
R22980 VSS.n8075 VSS.n8073 7.24
R22981 VSS.n8118 VSS.n8117 7.24
R22982 VSS.n8084 VSS.n8082 7.24
R22983 VSS.n8093 VSS.n8091 7.24
R22984 VSS.n7928 VSS.n7927 7.24
R22985 VSS.n7936 VSS.n7589 7.24
R22986 VSS.n7947 VSS.n7946 7.24
R22987 VSS.n7582 VSS.n7577 7.24
R22988 VSS.n7963 VSS.n7962 7.24
R22989 VSS.n7971 VSS.n7568 7.24
R22990 VSS.n7981 VSS.n7980 7.24
R22991 VSS.n7561 VSS.n7556 7.24
R22992 VSS.n7997 VSS.n7996 7.24
R22993 VSS.n8005 VSS.n7547 7.24
R22994 VSS.n8016 VSS.n8015 7.24
R22995 VSS.n7683 VSS.n7680 7.24
R22996 VSS.n7823 VSS.n7822 7.24
R22997 VSS.n7692 VSS.n7690 7.24
R22998 VSS.n7702 VSS.n7700 7.24
R22999 VSS.n7800 VSS.n7799 7.24
R23000 VSS.n7711 VSS.n7709 7.24
R23001 VSS.n7721 VSS.n7719 7.24
R23002 VSS.n7778 VSS.n7777 7.24
R23003 VSS.n7730 VSS.n7728 7.24
R23004 VSS.n7740 VSS.n7738 7.24
R23005 VSS.n7755 VSS.n7754 7.24
R23006 VSS.n5561 VSS.n5560 7.24
R23007 VSS.n5427 VSS.n5425 7.24
R23008 VSS.n5437 VSS.n5435 7.24
R23009 VSS.n5538 VSS.n5537 7.24
R23010 VSS.n5446 VSS.n5444 7.24
R23011 VSS.n5456 VSS.n5454 7.24
R23012 VSS.n5516 VSS.n5515 7.24
R23013 VSS.n5465 VSS.n5463 7.24
R23014 VSS.n5475 VSS.n5473 7.24
R23015 VSS.n5493 VSS.n5492 7.24
R23016 VSS.n5483 VSS.n5482 7.24
R23017 VSS.n5325 VSS.n3747 7.24
R23018 VSS.n5336 VSS.n5335 7.24
R23019 VSS.n3740 VSS.n3735 7.24
R23020 VSS.n5352 VSS.n5351 7.24
R23021 VSS.n5360 VSS.n3726 7.24
R23022 VSS.n5371 VSS.n5370 7.24
R23023 VSS.n3719 VSS.n3714 7.24
R23024 VSS.n5386 VSS.n5385 7.24
R23025 VSS.n5394 VSS.n3705 7.24
R23026 VSS.n5406 VSS.n5405 7.24
R23027 VSS.n5412 VSS.n5411 7.24
R23028 VSS.n5215 VSS.n5214 7.24
R23029 VSS.n5070 VSS.n5068 7.24
R23030 VSS.n5080 VSS.n5078 7.24
R23031 VSS.n5192 VSS.n5191 7.24
R23032 VSS.n5089 VSS.n5087 7.24
R23033 VSS.n5099 VSS.n5097 7.24
R23034 VSS.n5170 VSS.n5169 7.24
R23035 VSS.n5108 VSS.n5106 7.24
R23036 VSS.n5118 VSS.n5116 7.24
R23037 VSS.n5147 VSS.n5146 7.24
R23038 VSS.n5128 VSS.n5125 7.24
R23039 VSS.n4968 VSS.n3888 7.24
R23040 VSS.n4979 VSS.n4978 7.24
R23041 VSS.n3881 VSS.n3876 7.24
R23042 VSS.n4995 VSS.n4994 7.24
R23043 VSS.n5003 VSS.n3867 7.24
R23044 VSS.n5014 VSS.n5013 7.24
R23045 VSS.n3860 VSS.n3855 7.24
R23046 VSS.n5029 VSS.n5028 7.24
R23047 VSS.n5037 VSS.n3846 7.24
R23048 VSS.n5049 VSS.n5048 7.24
R23049 VSS.n5055 VSS.n5054 7.24
R23050 VSS.n4858 VSS.n4857 7.24
R23051 VSS.n4713 VSS.n4711 7.24
R23052 VSS.n4723 VSS.n4721 7.24
R23053 VSS.n4835 VSS.n4834 7.24
R23054 VSS.n4732 VSS.n4730 7.24
R23055 VSS.n4742 VSS.n4740 7.24
R23056 VSS.n4813 VSS.n4812 7.24
R23057 VSS.n4751 VSS.n4749 7.24
R23058 VSS.n4761 VSS.n4759 7.24
R23059 VSS.n4790 VSS.n4789 7.24
R23060 VSS.n4771 VSS.n4768 7.24
R23061 VSS.n4611 VSS.n4029 7.24
R23062 VSS.n4622 VSS.n4621 7.24
R23063 VSS.n4022 VSS.n4017 7.24
R23064 VSS.n4638 VSS.n4637 7.24
R23065 VSS.n4646 VSS.n4008 7.24
R23066 VSS.n4657 VSS.n4656 7.24
R23067 VSS.n4001 VSS.n3996 7.24
R23068 VSS.n4672 VSS.n4671 7.24
R23069 VSS.n4680 VSS.n3987 7.24
R23070 VSS.n4692 VSS.n4691 7.24
R23071 VSS.n4698 VSS.n4697 7.24
R23072 VSS.n4501 VSS.n4500 7.24
R23073 VSS.n4356 VSS.n4354 7.24
R23074 VSS.n4366 VSS.n4364 7.24
R23075 VSS.n4478 VSS.n4477 7.24
R23076 VSS.n4375 VSS.n4373 7.24
R23077 VSS.n4385 VSS.n4383 7.24
R23078 VSS.n4456 VSS.n4455 7.24
R23079 VSS.n4394 VSS.n4392 7.24
R23080 VSS.n4404 VSS.n4402 7.24
R23081 VSS.n4433 VSS.n4432 7.24
R23082 VSS.n4414 VSS.n4411 7.24
R23083 VSS.n4254 VSS.n4170 7.24
R23084 VSS.n4265 VSS.n4264 7.24
R23085 VSS.n4163 VSS.n4158 7.24
R23086 VSS.n4281 VSS.n4280 7.24
R23087 VSS.n4289 VSS.n4149 7.24
R23088 VSS.n4300 VSS.n4299 7.24
R23089 VSS.n4142 VSS.n4137 7.24
R23090 VSS.n4315 VSS.n4314 7.24
R23091 VSS.n4323 VSS.n4128 7.24
R23092 VSS.n4335 VSS.n4334 7.24
R23093 VSS.n4341 VSS.n4340 7.24
R23094 VSS.n2813 VSS.n2811 7.24
R23095 VSS.n2951 VSS.n2950 7.24
R23096 VSS.n2822 VSS.n2820 7.24
R23097 VSS.n2832 VSS.n2830 7.24
R23098 VSS.n2928 VSS.n2927 7.24
R23099 VSS.n2841 VSS.n2839 7.24
R23100 VSS.n2851 VSS.n2849 7.24
R23101 VSS.n2906 VSS.n2905 7.24
R23102 VSS.n2860 VSS.n2858 7.24
R23103 VSS.n2870 VSS.n2868 7.24
R23104 VSS.n2883 VSS.n2882 7.24
R23105 VSS.n2706 VSS.n2705 7.24
R23106 VSS.n1368 VSS.n1363 7.24
R23107 VSS.n2722 VSS.n2721 7.24
R23108 VSS.n2730 VSS.n1354 7.24
R23109 VSS.n2741 VSS.n2740 7.24
R23110 VSS.n1347 VSS.n1342 7.24
R23111 VSS.n2756 VSS.n2755 7.24
R23112 VSS.n2764 VSS.n1333 7.24
R23113 VSS.n2775 VSS.n2774 7.24
R23114 VSS.n1326 VSS.n1321 7.24
R23115 VSS.n2791 VSS.n2790 7.24
R23116 VSS.n2338 VSS.n2336 7.24
R23117 VSS.n2459 VSS.n2458 7.24
R23118 VSS.n2347 VSS.n2345 7.24
R23119 VSS.n2357 VSS.n2355 7.24
R23120 VSS.n2436 VSS.n2435 7.24
R23121 VSS.n2366 VSS.n2364 7.24
R23122 VSS.n2376 VSS.n2374 7.24
R23123 VSS.n2414 VSS.n2413 7.24
R23124 VSS.n2385 VSS.n2383 7.24
R23125 VSS.n2392 VSS.n2391 7.24
R23126 VSS.n2689 VSS.n2688 7.24
R23127 VSS.n2226 VSS.n2224 7.24
R23128 VSS.n2551 VSS.n2550 7.24
R23129 VSS.n2235 VSS.n2233 7.24
R23130 VSS.n2245 VSS.n2243 7.24
R23131 VSS.n2528 VSS.n2527 7.24
R23132 VSS.n2254 VSS.n2252 7.24
R23133 VSS.n2264 VSS.n2262 7.24
R23134 VSS.n2506 VSS.n2505 7.24
R23135 VSS.n2273 VSS.n2271 7.24
R23136 VSS.n2283 VSS.n2281 7.24
R23137 VSS.n2483 VSS.n2482 7.24
R23138 VSS.n2124 VSS.n2123 7.24
R23139 VSS.n2132 VSS.n1531 7.24
R23140 VSS.n2143 VSS.n2142 7.24
R23141 VSS.n1524 VSS.n1519 7.24
R23142 VSS.n2159 VSS.n2158 7.24
R23143 VSS.n2167 VSS.n1510 7.24
R23144 VSS.n2177 VSS.n2176 7.24
R23145 VSS.n1503 VSS.n1498 7.24
R23146 VSS.n2193 VSS.n2192 7.24
R23147 VSS.n2201 VSS.n1489 7.24
R23148 VSS.n2212 VSS.n2211 7.24
R23149 VSS.n1729 VSS.n1727 7.24
R23150 VSS.n1858 VSS.n1857 7.24
R23151 VSS.n1738 VSS.n1736 7.24
R23152 VSS.n1748 VSS.n1746 7.24
R23153 VSS.n1835 VSS.n1834 7.24
R23154 VSS.n1757 VSS.n1755 7.24
R23155 VSS.n1767 VSS.n1765 7.24
R23156 VSS.n1813 VSS.n1812 7.24
R23157 VSS.n1776 VSS.n1774 7.24
R23158 VSS.n1790 VSS.n1784 7.24
R23159 VSS.n1788 VSS.n1787 7.24
R23160 VSS.n1617 VSS.n1614 7.24
R23161 VSS.n1950 VSS.n1949 7.24
R23162 VSS.n1626 VSS.n1624 7.24
R23163 VSS.n1636 VSS.n1634 7.24
R23164 VSS.n1927 VSS.n1926 7.24
R23165 VSS.n1645 VSS.n1643 7.24
R23166 VSS.n1655 VSS.n1653 7.24
R23167 VSS.n1905 VSS.n1904 7.24
R23168 VSS.n1664 VSS.n1662 7.24
R23169 VSS.n1674 VSS.n1672 7.24
R23170 VSS.n1882 VSS.n1881 7.24
R23171 VSS.n17486 sky130_asc_res_xhigh_po_2p85_1_16/VGND 7.16
R23172 VSS.n13966 sky130_asc_res_xhigh_po_2p85_1_17/VGND 7.159
R23173 VSS.n17330 VSS.n17329 7.111
R23174 VSS.n17222 VSS.n16141 7.111
R23175 VSS.n17132 VSS.n16231 7.111
R23176 VSS.n17042 VSS.n16321 7.111
R23177 VSS.n16952 VSS.n16411 7.111
R23178 VSS.n16862 VSS.n16501 7.111
R23179 VSS.n16772 VSS.n16591 7.111
R23180 VSS.n16682 VSS.n16681 7.111
R23181 VSS.n11149 VSS.n11148 7.111
R23182 VSS.n11239 VSS.n11058 7.111
R23183 VSS.n11329 VSS.n10968 7.111
R23184 VSS.n11419 VSS.n10878 7.111
R23185 VSS.n13539 VSS.n10788 7.111
R23186 VSS.n13629 VSS.n10698 7.111
R23187 VSS.n13719 VSS.n10608 7.111
R23188 VSS.n13827 VSS.n13826 7.111
R23189 VSS.n9159 VSS.n8982 7.111
R23190 VSS.n10177 VSS.n9276 7.111
R23191 VSS.n10087 VSS.n9366 7.111
R23192 VSS.n9997 VSS.n9456 7.111
R23193 VSS.n9907 VSS.n9546 7.111
R23194 VSS.n9817 VSS.n9636 7.111
R23195 VSS.n9727 VSS.n9726 7.111
R23196 VSS.n10317 VSS.n10316 7.111
R23197 VSS.n5684 VSS.n3577 7.111
R23198 VSS.n5806 VSS.n3519 7.111
R23199 VSS.n5928 VSS.n3461 7.111
R23200 VSS.n6050 VSS.n3403 7.111
R23201 VSS.n6172 VSS.n3345 7.111
R23202 VSS.n6294 VSS.n3287 7.111
R23203 VSS.n6416 VSS.n3229 7.111
R23204 VSS.n6539 VSS.n6538 7.111
R23205 VSS.n1175 VSS.n94 7.111
R23206 VSS.n1085 VSS.n184 7.111
R23207 VSS.n995 VSS.n274 7.111
R23208 VSS.n905 VSS.n364 7.111
R23209 VSS.n815 VSS.n454 7.111
R23210 VSS.n725 VSS.n544 7.111
R23211 VSS.n635 VSS.n634 7.111
R23212 sky130_asc_pnp_05v5_W3p40L3p40_1_0/VGND VSS.n6899 7.109
R23213 VSS.n16682 VSS.n16633 6.925
R23214 VSS.n11149 VSS.n11100 6.925
R23215 VSS.n9727 VSS.n9678 6.925
R23216 VSS.n6538 VSS.n3136 6.925
R23217 VSS.n635 VSS.n586 6.925
R23218 VSS.n17329 VSS.n17311 6.783
R23219 VSS.n17222 VSS.n17221 6.783
R23220 VSS.n17132 VSS.n17131 6.783
R23221 VSS.n17042 VSS.n17041 6.783
R23222 VSS.n16952 VSS.n16951 6.783
R23223 VSS.n16862 VSS.n16861 6.783
R23224 VSS.n16772 VSS.n16771 6.783
R23225 VSS.n11239 VSS.n11238 6.783
R23226 VSS.n11329 VSS.n11328 6.783
R23227 VSS.n11419 VSS.n11418 6.783
R23228 VSS.n13539 VSS.n13538 6.783
R23229 VSS.n13629 VSS.n13628 6.783
R23230 VSS.n13719 VSS.n13718 6.783
R23231 VSS.n13826 VSS.n13808 6.783
R23232 VSS.n9160 VSS.n9159 6.783
R23233 VSS.n10177 VSS.n10176 6.783
R23234 VSS.n10087 VSS.n10086 6.783
R23235 VSS.n9997 VSS.n9996 6.783
R23236 VSS.n9907 VSS.n9906 6.783
R23237 VSS.n9817 VSS.n9816 6.783
R23238 VSS.n10318 VSS.n10317 6.783
R23239 VSS.n5786 VSS.n3577 6.783
R23240 VSS.n5908 VSS.n3519 6.783
R23241 VSS.n6030 VSS.n3461 6.783
R23242 VSS.n6152 VSS.n3403 6.783
R23243 VSS.n6274 VSS.n3345 6.783
R23244 VSS.n6396 VSS.n3287 6.783
R23245 VSS.n6518 VSS.n3229 6.783
R23246 VSS.n1175 VSS.n1174 6.783
R23247 VSS.n1085 VSS.n1084 6.783
R23248 VSS.n995 VSS.n994 6.783
R23249 VSS.n905 VSS.n904 6.783
R23250 VSS.n815 VSS.n814 6.783
R23251 VSS.n725 VSS.n724 6.783
R23252 VSS.n17600 VSS.n3051 6.743
R23253 VSS.n15950 VSS.n15949 6.723
R23254 VSS.n15922 VSS.n14054 6.723
R23255 VSS.n14191 VSS.n14157 6.723
R23256 VSS.n15385 VSS.n14204 6.723
R23257 VSS.n15360 VSS.n15359 6.723
R23258 VSS.n14839 VSS.n14321 6.723
R23259 VSS.n14780 VSS.n14779 6.723
R23260 VSS.n12165 VSS.n12164 6.723
R23261 VSS.n12434 VSS.n11528 6.723
R23262 VSS.n12459 VSS.n12458 6.723
R23263 VSS.n12485 VSS.n11496 6.723
R23264 VSS.n13341 VSS.n12498 6.723
R23265 VSS.n12626 VSS.n12597 6.723
R23266 VSS.n13092 VSS.n12639 6.723
R23267 VSS.n8828 VSS.n7226 6.723
R23268 VSS.n8804 VSS.n8803 6.723
R23269 VSS.n8606 VSS.n7366 6.723
R23270 VSS.n8582 VSS.n8581 6.723
R23271 VSS.n8248 VSS.n7506 6.723
R23272 VSS.n8224 VSS.n8223 6.723
R23273 VSS.n7890 VSS.n7646 6.723
R23274 VSS.n5605 VSS.n3669 6.723
R23275 VSS.n3797 VSS.n3768 6.723
R23276 VSS.n5259 VSS.n3810 6.723
R23277 VSS.n3938 VSS.n3909 6.723
R23278 VSS.n4902 VSS.n3951 6.723
R23279 VSS.n4079 VSS.n4050 6.723
R23280 VSS.n4545 VSS.n4092 6.723
R23281 VSS.n2996 VSS.n1295 6.723
R23282 VSS.n1432 VSS.n1398 6.723
R23283 VSS.n2626 VSS.n1445 6.723
R23284 VSS.n2601 VSS.n2600 6.723
R23285 VSS.n2080 VSS.n1562 6.723
R23286 VSS.n2021 VSS.n2020 6.723
R23287 sky130_asc_res_xhigh_po_2p85_2_0/VGND VSS.n17524 6.663
R23288 sky130_asc_res_xhigh_po_2p85_1_22/VGND VSS.n17480 6.66
R23289 sky130_asc_pfet_01v8_lvt_6_0/VGND VSS.n10488 6.659
R23290 VSS.n10373 sky130_asc_res_xhigh_po_2p85_1_8/VGND 6.654
R23291 sky130_asc_res_xhigh_po_2p85_1_19/VGND VSS.n17599 6.654
R23292 sky130_asc_res_xhigh_po_2p85_1_1/VGND sky130_asc_res_xhigh_po_2p85_2_1/VGND 6.609
R23293 VSS.n17480 VSS.n17479 6.532
R23294 VSS.n1267 sky130_asc_nfet_01v8_lvt_1_1/SOURCE 6.4
R23295 VSS.n17524 VSS.n17523 6.345
R23296 VSS.n6608 VSS.n6607 6.316
R23297 VSS.n3085 sky130_asc_res_xhigh_po_2p85_1_18/VGND 6.245
R23298 sky130_asc_cap_mim_m3_1_5/VGND sky130_asc_pfet_01v8_lvt_12_0/VGND 6.208
R23299 sky130_asc_cap_mim_m3_1_9/VGND sky130_asc_pfet_01v8_lvt_12_1/VGND 6.207
R23300 VSS.n15949 VSS.n14039 6.206
R23301 VSS.n14169 VSS.n14054 6.206
R23302 VSS.n15411 VSS.n14157 6.206
R23303 VSS.n15385 VSS.n15384 6.206
R23304 VSS.n15359 VSS.n14223 6.206
R23305 VSS.n14839 VSS.n14838 6.206
R23306 VSS.n14779 VSS.n14335 6.206
R23307 VSS.n12164 VSS.n12088 6.206
R23308 VSS.n12435 VSS.n12434 6.206
R23309 VSS.n12459 VSS.n11508 6.206
R23310 VSS.n13367 VSS.n11496 6.206
R23311 VSS.n13342 VSS.n13341 6.206
R23312 VSS.n13118 VSS.n12597 6.206
R23313 VSS.n13093 VSS.n13092 6.206
R23314 VSS.n8828 VSS.n8827 6.206
R23315 VSS.n8803 VSS.n8802 6.206
R23316 VSS.n8606 VSS.n8605 6.206
R23317 VSS.n8581 VSS.n8580 6.206
R23318 VSS.n8248 VSS.n8247 6.206
R23319 VSS.n8223 VSS.n8222 6.206
R23320 VSS.n7890 VSS.n7889 6.206
R23321 VSS.n5606 VSS.n5605 6.206
R23322 VSS.n5285 VSS.n3768 6.206
R23323 VSS.n5260 VSS.n5259 6.206
R23324 VSS.n4928 VSS.n3909 6.206
R23325 VSS.n4903 VSS.n4902 6.206
R23326 VSS.n4571 VSS.n4050 6.206
R23327 VSS.n4546 VSS.n4545 6.206
R23328 VSS.n1410 VSS.n1295 6.206
R23329 VSS.n2652 VSS.n1398 6.206
R23330 VSS.n2626 VSS.n2625 6.206
R23331 VSS.n2600 VSS.n1464 6.206
R23332 VSS.n2080 VSS.n2079 6.206
R23333 VSS.n2020 VSS.n1576 6.206
R23334 VSS.n15999 VSS.n15998 6.201
R23335 VSS.n12214 VSS.n12213 6.201
R23336 VSS.n7178 VSS.n7177 6.201
R23337 VSS.n3648 VSS.n3647 6.201
R23338 VSS.n3046 VSS.n3045 6.201
R23339 VSS.n13961 VSS.n13960 6.137
R23340 VSS.n1264 VSS.n1263 5.922
R23341 VSS.n17467 VSS.n17466 5.903
R23342 VSS.n15676 VSS.n15670 5.818
R23343 VSS.n15891 VSS.n14071 5.818
R23344 VSS.n15454 VSS.n14134 5.818
R23345 VSS.n15089 VSS.n15083 5.818
R23346 VSS.n14976 VSS.n14236 5.818
R23347 VSS.n14865 VSS.n14299 5.818
R23348 VSS.n14480 VSS.n14474 5.818
R23349 VSS.n11990 VSS.n11984 5.818
R23350 VSS.n11910 VSS.n11541 5.818
R23351 VSS.n11775 VSS.n11604 5.818
R23352 VSS.n13398 VSS.n11481 5.818
R23353 VSS.n13314 VSS.n12517 5.818
R23354 VSS.n13150 VSS.n13149 5.818
R23355 VSS.n13065 VSS.n12658 5.818
R23356 VSS.n7068 VSS.n6968 5.818
R23357 VSS.n8764 VSS.n8763 5.818
R23358 VSS.n7324 VSS.n7318 5.818
R23359 VSS.n8542 VSS.n8541 5.818
R23360 VSS.n7464 VSS.n7458 5.818
R23361 VSS.n8184 VSS.n8183 5.818
R23362 VSS.n7604 VSS.n7598 5.818
R23363 VSS.n5578 VSS.n3688 5.818
R23364 VSS.n5317 VSS.n5316 5.818
R23365 VSS.n5232 VSS.n3829 5.818
R23366 VSS.n4960 VSS.n4959 5.818
R23367 VSS.n4875 VSS.n3970 5.818
R23368 VSS.n4603 VSS.n4602 5.818
R23369 VSS.n4518 VSS.n4111 5.818
R23370 VSS.n2965 VSS.n1312 5.818
R23371 VSS.n2695 VSS.n1375 5.818
R23372 VSS.n2330 VSS.n2324 5.818
R23373 VSS.n2217 VSS.n1477 5.818
R23374 VSS.n2106 VSS.n1540 5.818
R23375 VSS.n1721 VSS.n1715 5.818
R23376 VSS.n17721 sky130_asc_res_xhigh_po_2p85_1_3/VGND 5.76
R23377 VSS.n17720 sky130_asc_res_xhigh_po_2p85_1_4/VGND 5.76
R23378 sky130_asc_res_xhigh_po_2p85_1_1/VGND VSS.n17722 5.75
R23379 VSS.n17385 VSS.n16036 5.655
R23380 VSS.n17327 VSS.n16036 5.655
R23381 VSS.n11089 VSS.n11083 5.655
R23382 VSS.n11150 VSS.n11089 5.655
R23383 VSS.n10999 VSS.n10993 5.655
R23384 VSS.n11240 VSS.n10999 5.655
R23385 VSS.n10909 VSS.n10903 5.655
R23386 VSS.n11330 VSS.n10909 5.655
R23387 VSS.n10819 VSS.n10813 5.655
R23388 VSS.n11420 VSS.n10819 5.655
R23389 VSS.n10729 VSS.n10723 5.655
R23390 VSS.n13540 VSS.n10729 5.655
R23391 VSS.n10639 VSS.n10633 5.655
R23392 VSS.n13630 VSS.n10639 5.655
R23393 VSS.n10549 VSS.n10543 5.655
R23394 VSS.n13720 VSS.n10549 5.655
R23395 VSS.n13885 VSS.n10504 5.655
R23396 VSS.n13824 VSS.n10504 5.655
R23397 VSS.n10323 VSS.n9179 5.655
R23398 VSS.n10314 VSS.n9179 5.655
R23399 VSS.n10444 VSS.n10443 5.647
R23400 VSS.n10469 VSS.n10468 5.647
R23401 VSS.n17677 VSS.n17651 5.647
R23402 VSS.n17685 VSS.n17684 5.647
R23403 sky130_asc_pnp_05v5_W3p40L3p40_8_2/VGND sky130_asc_nfet_01v8_lvt_9_1/VGND 5.497
R23404 sky130_asc_pnp_05v5_W3p40L3p40_8_1/VGND sky130_asc_nfet_01v8_lvt_9_2/VGND 5.497
R23405 VSS.n17460 VSS.n16044 5.446
R23406 VSS.n17460 VSS.n16045 5.446
R23407 VSS.n17460 VSS.n16043 5.446
R23408 VSS.n17460 VSS.n16046 5.446
R23409 VSS.n17460 VSS.n16042 5.446
R23410 VSS.n17460 VSS.n17459 5.446
R23411 VSS.n17460 VSS.n16041 5.446
R23412 VSS.n17460 VSS.n16040 5.446
R23413 VSS.n17305 VSS.n16086 5.446
R23414 VSS.n17305 VSS.n16087 5.446
R23415 VSS.n17305 VSS.n16085 5.446
R23416 VSS.n17305 VSS.n16088 5.446
R23417 VSS.n17305 VSS.n16084 5.446
R23418 VSS.n17305 VSS.n16089 5.446
R23419 VSS.n17305 VSS.n16083 5.446
R23420 VSS.n17305 VSS.n17303 5.446
R23421 VSS.n17215 VSS.n16176 5.446
R23422 VSS.n17215 VSS.n16177 5.446
R23423 VSS.n17215 VSS.n16175 5.446
R23424 VSS.n17215 VSS.n16178 5.446
R23425 VSS.n17215 VSS.n16174 5.446
R23426 VSS.n17215 VSS.n16179 5.446
R23427 VSS.n17215 VSS.n16173 5.446
R23428 VSS.n17215 VSS.n17213 5.446
R23429 VSS.n17125 VSS.n16266 5.446
R23430 VSS.n17125 VSS.n16267 5.446
R23431 VSS.n17125 VSS.n16265 5.446
R23432 VSS.n17125 VSS.n16268 5.446
R23433 VSS.n17125 VSS.n16264 5.446
R23434 VSS.n17125 VSS.n16269 5.446
R23435 VSS.n17125 VSS.n16263 5.446
R23436 VSS.n17125 VSS.n17123 5.446
R23437 VSS.n17035 VSS.n16356 5.446
R23438 VSS.n17035 VSS.n16357 5.446
R23439 VSS.n17035 VSS.n16355 5.446
R23440 VSS.n17035 VSS.n16358 5.446
R23441 VSS.n17035 VSS.n16354 5.446
R23442 VSS.n17035 VSS.n16359 5.446
R23443 VSS.n17035 VSS.n16353 5.446
R23444 VSS.n17035 VSS.n17033 5.446
R23445 VSS.n16945 VSS.n16446 5.446
R23446 VSS.n16945 VSS.n16447 5.446
R23447 VSS.n16945 VSS.n16445 5.446
R23448 VSS.n16945 VSS.n16448 5.446
R23449 VSS.n16945 VSS.n16444 5.446
R23450 VSS.n16945 VSS.n16449 5.446
R23451 VSS.n16945 VSS.n16443 5.446
R23452 VSS.n16945 VSS.n16943 5.446
R23453 VSS.n16855 VSS.n16536 5.446
R23454 VSS.n16855 VSS.n16537 5.446
R23455 VSS.n16855 VSS.n16535 5.446
R23456 VSS.n16855 VSS.n16538 5.446
R23457 VSS.n16855 VSS.n16534 5.446
R23458 VSS.n16855 VSS.n16539 5.446
R23459 VSS.n16855 VSS.n16533 5.446
R23460 VSS.n16855 VSS.n16853 5.446
R23461 VSS.n16765 VSS.n16626 5.446
R23462 VSS.n16765 VSS.n16627 5.446
R23463 VSS.n16765 VSS.n16625 5.446
R23464 VSS.n16765 VSS.n16628 5.446
R23465 VSS.n16765 VSS.n16624 5.446
R23466 VSS.n16765 VSS.n16629 5.446
R23467 VSS.n16765 VSS.n16623 5.446
R23468 VSS.n16765 VSS.n16763 5.446
R23469 VSS.n11232 VSS.n11093 5.446
R23470 VSS.n11232 VSS.n11094 5.446
R23471 VSS.n11232 VSS.n11092 5.446
R23472 VSS.n11232 VSS.n11095 5.446
R23473 VSS.n11232 VSS.n11091 5.446
R23474 VSS.n11232 VSS.n11096 5.446
R23475 VSS.n11232 VSS.n11090 5.446
R23476 VSS.n11232 VSS.n11231 5.446
R23477 VSS.n11322 VSS.n11003 5.446
R23478 VSS.n11322 VSS.n11004 5.446
R23479 VSS.n11322 VSS.n11002 5.446
R23480 VSS.n11322 VSS.n11005 5.446
R23481 VSS.n11322 VSS.n11001 5.446
R23482 VSS.n11322 VSS.n11006 5.446
R23483 VSS.n11322 VSS.n11000 5.446
R23484 VSS.n11322 VSS.n11321 5.446
R23485 VSS.n11412 VSS.n10913 5.446
R23486 VSS.n11412 VSS.n10914 5.446
R23487 VSS.n11412 VSS.n10912 5.446
R23488 VSS.n11412 VSS.n10915 5.446
R23489 VSS.n11412 VSS.n10911 5.446
R23490 VSS.n11412 VSS.n10916 5.446
R23491 VSS.n11412 VSS.n10910 5.446
R23492 VSS.n11412 VSS.n11411 5.446
R23493 VSS.n13532 VSS.n10823 5.446
R23494 VSS.n13532 VSS.n10824 5.446
R23495 VSS.n13532 VSS.n10822 5.446
R23496 VSS.n13532 VSS.n10825 5.446
R23497 VSS.n13532 VSS.n10821 5.446
R23498 VSS.n13532 VSS.n10826 5.446
R23499 VSS.n13532 VSS.n10820 5.446
R23500 VSS.n13532 VSS.n13531 5.446
R23501 VSS.n13622 VSS.n10733 5.446
R23502 VSS.n13622 VSS.n10734 5.446
R23503 VSS.n13622 VSS.n10732 5.446
R23504 VSS.n13622 VSS.n10735 5.446
R23505 VSS.n13622 VSS.n10731 5.446
R23506 VSS.n13622 VSS.n10736 5.446
R23507 VSS.n13622 VSS.n10730 5.446
R23508 VSS.n13622 VSS.n13621 5.446
R23509 VSS.n13712 VSS.n10643 5.446
R23510 VSS.n13712 VSS.n10644 5.446
R23511 VSS.n13712 VSS.n10642 5.446
R23512 VSS.n13712 VSS.n10645 5.446
R23513 VSS.n13712 VSS.n10641 5.446
R23514 VSS.n13712 VSS.n10646 5.446
R23515 VSS.n13712 VSS.n10640 5.446
R23516 VSS.n13712 VSS.n13711 5.446
R23517 VSS.n13802 VSS.n10553 5.446
R23518 VSS.n13802 VSS.n10554 5.446
R23519 VSS.n13802 VSS.n10552 5.446
R23520 VSS.n13802 VSS.n10555 5.446
R23521 VSS.n13802 VSS.n10551 5.446
R23522 VSS.n13802 VSS.n10556 5.446
R23523 VSS.n13802 VSS.n10550 5.446
R23524 VSS.n13802 VSS.n13801 5.446
R23525 VSS.n13952 VSS.n10511 5.446
R23526 VSS.n13952 VSS.n10512 5.446
R23527 VSS.n13952 VSS.n10510 5.446
R23528 VSS.n13952 VSS.n10513 5.446
R23529 VSS.n13952 VSS.n10509 5.446
R23530 VSS.n13952 VSS.n13951 5.446
R23531 VSS.n13952 VSS.n10508 5.446
R23532 VSS.n13952 VSS.n10495 5.446
R23533 VSS.t20 VSS.n9010 5.446
R23534 VSS.t20 VSS.n9011 5.446
R23535 VSS.t20 VSS.n9009 5.446
R23536 VSS.t20 VSS.n9012 5.446
R23537 VSS.t20 VSS.n9013 5.446
R23538 VSS.t20 VSS.n9008 5.446
R23539 VSS.t20 VSS.n9014 5.446
R23540 VSS.t20 VSS.n9007 5.446
R23541 VSS.n10260 VSS.n9221 5.446
R23542 VSS.n10260 VSS.n9222 5.446
R23543 VSS.n10260 VSS.n9220 5.446
R23544 VSS.n10260 VSS.n9223 5.446
R23545 VSS.n10260 VSS.n9219 5.446
R23546 VSS.n10260 VSS.n9224 5.446
R23547 VSS.n10260 VSS.n9218 5.446
R23548 VSS.n10260 VSS.n10258 5.446
R23549 VSS.n10170 VSS.n9311 5.446
R23550 VSS.n10170 VSS.n9312 5.446
R23551 VSS.n10170 VSS.n9310 5.446
R23552 VSS.n10170 VSS.n9313 5.446
R23553 VSS.n10170 VSS.n9309 5.446
R23554 VSS.n10170 VSS.n9314 5.446
R23555 VSS.n10170 VSS.n9308 5.446
R23556 VSS.n10170 VSS.n10168 5.446
R23557 VSS.n10080 VSS.n9401 5.446
R23558 VSS.n10080 VSS.n9402 5.446
R23559 VSS.n10080 VSS.n9400 5.446
R23560 VSS.n10080 VSS.n9403 5.446
R23561 VSS.n10080 VSS.n9399 5.446
R23562 VSS.n10080 VSS.n9404 5.446
R23563 VSS.n10080 VSS.n9398 5.446
R23564 VSS.n10080 VSS.n10078 5.446
R23565 VSS.n9990 VSS.n9491 5.446
R23566 VSS.n9990 VSS.n9492 5.446
R23567 VSS.n9990 VSS.n9490 5.446
R23568 VSS.n9990 VSS.n9493 5.446
R23569 VSS.n9990 VSS.n9489 5.446
R23570 VSS.n9990 VSS.n9494 5.446
R23571 VSS.n9990 VSS.n9488 5.446
R23572 VSS.n9990 VSS.n9988 5.446
R23573 VSS.n9900 VSS.n9581 5.446
R23574 VSS.n9900 VSS.n9582 5.446
R23575 VSS.n9900 VSS.n9580 5.446
R23576 VSS.n9900 VSS.n9583 5.446
R23577 VSS.n9900 VSS.n9579 5.446
R23578 VSS.n9900 VSS.n9584 5.446
R23579 VSS.n9900 VSS.n9578 5.446
R23580 VSS.n9900 VSS.n9898 5.446
R23581 VSS.n9810 VSS.n9671 5.446
R23582 VSS.n9810 VSS.n9672 5.446
R23583 VSS.n9810 VSS.n9670 5.446
R23584 VSS.n9810 VSS.n9673 5.446
R23585 VSS.n9810 VSS.n9669 5.446
R23586 VSS.n9810 VSS.n9674 5.446
R23587 VSS.n9810 VSS.n9668 5.446
R23588 VSS.n9810 VSS.n9808 5.446
R23589 VSS.n10331 VSS.n8935 5.446
R23590 VSS.n10337 VSS.n8935 5.446
R23591 VSS.n10343 VSS.n8935 5.446
R23592 VSS.n10349 VSS.n8935 5.446
R23593 VSS.n10355 VSS.n8935 5.446
R23594 VSS.n10361 VSS.n8935 5.446
R23595 VSS.n10367 VSS.n8935 5.446
R23596 VSS.n9182 VSS.n8935 5.446
R23597 VSS.n5740 VSS.n3582 5.446
R23598 VSS.n5746 VSS.n3582 5.446
R23599 VSS.n5752 VSS.n3582 5.446
R23600 VSS.n5758 VSS.n3582 5.446
R23601 VSS.n5764 VSS.n3582 5.446
R23602 VSS.n5770 VSS.n3582 5.446
R23603 VSS.n5776 VSS.n3582 5.446
R23604 VSS.n5782 VSS.n3582 5.446
R23605 VSS.n5862 VSS.n3524 5.446
R23606 VSS.n5868 VSS.n3524 5.446
R23607 VSS.n5874 VSS.n3524 5.446
R23608 VSS.n5880 VSS.n3524 5.446
R23609 VSS.n5886 VSS.n3524 5.446
R23610 VSS.n5892 VSS.n3524 5.446
R23611 VSS.n5898 VSS.n3524 5.446
R23612 VSS.n5904 VSS.n3524 5.446
R23613 VSS.n5984 VSS.n3466 5.446
R23614 VSS.n5990 VSS.n3466 5.446
R23615 VSS.n5996 VSS.n3466 5.446
R23616 VSS.n6002 VSS.n3466 5.446
R23617 VSS.n6008 VSS.n3466 5.446
R23618 VSS.n6014 VSS.n3466 5.446
R23619 VSS.n6020 VSS.n3466 5.446
R23620 VSS.n6026 VSS.n3466 5.446
R23621 VSS.n6106 VSS.n3408 5.446
R23622 VSS.n6112 VSS.n3408 5.446
R23623 VSS.n6118 VSS.n3408 5.446
R23624 VSS.n6124 VSS.n3408 5.446
R23625 VSS.n6130 VSS.n3408 5.446
R23626 VSS.n6136 VSS.n3408 5.446
R23627 VSS.n6142 VSS.n3408 5.446
R23628 VSS.n6148 VSS.n3408 5.446
R23629 VSS.n6228 VSS.n3350 5.446
R23630 VSS.n6234 VSS.n3350 5.446
R23631 VSS.n6240 VSS.n3350 5.446
R23632 VSS.n6246 VSS.n3350 5.446
R23633 VSS.n6252 VSS.n3350 5.446
R23634 VSS.n6258 VSS.n3350 5.446
R23635 VSS.n6264 VSS.n3350 5.446
R23636 VSS.n6270 VSS.n3350 5.446
R23637 VSS.n6350 VSS.n3292 5.446
R23638 VSS.n6356 VSS.n3292 5.446
R23639 VSS.n6362 VSS.n3292 5.446
R23640 VSS.n6368 VSS.n3292 5.446
R23641 VSS.n6374 VSS.n3292 5.446
R23642 VSS.n6380 VSS.n3292 5.446
R23643 VSS.n6386 VSS.n3292 5.446
R23644 VSS.n6392 VSS.n3292 5.446
R23645 VSS.n6472 VSS.n3234 5.446
R23646 VSS.n6478 VSS.n3234 5.446
R23647 VSS.n6484 VSS.n3234 5.446
R23648 VSS.n6490 VSS.n3234 5.446
R23649 VSS.n6496 VSS.n3234 5.446
R23650 VSS.n6502 VSS.n3234 5.446
R23651 VSS.n6508 VSS.n3234 5.446
R23652 VSS.n6514 VSS.n3234 5.446
R23653 VSS.n6598 VSS.n3153 5.446
R23654 VSS.n6598 VSS.n3154 5.446
R23655 VSS.n6598 VSS.n3152 5.446
R23656 VSS.n6598 VSS.n3155 5.446
R23657 VSS.n6598 VSS.n3151 5.446
R23658 VSS.n6598 VSS.n3156 5.446
R23659 VSS.n6598 VSS.n3150 5.446
R23660 VSS.n6598 VSS.n3140 5.446
R23661 VSS.n1252 VSS.n38 5.446
R23662 VSS.n1252 VSS.n39 5.446
R23663 VSS.n1252 VSS.n37 5.446
R23664 VSS.n1252 VSS.n40 5.446
R23665 VSS.n1252 VSS.n36 5.446
R23666 VSS.n1252 VSS.n41 5.446
R23667 VSS.n1252 VSS.n35 5.446
R23668 VSS.n1252 VSS.n1251 5.446
R23669 VSS.n1168 VSS.n129 5.446
R23670 VSS.n1168 VSS.n130 5.446
R23671 VSS.n1168 VSS.n128 5.446
R23672 VSS.n1168 VSS.n131 5.446
R23673 VSS.n1168 VSS.n127 5.446
R23674 VSS.n1168 VSS.n132 5.446
R23675 VSS.n1168 VSS.n126 5.446
R23676 VSS.n1168 VSS.n1166 5.446
R23677 VSS.n1078 VSS.n219 5.446
R23678 VSS.n1078 VSS.n220 5.446
R23679 VSS.n1078 VSS.n218 5.446
R23680 VSS.n1078 VSS.n221 5.446
R23681 VSS.n1078 VSS.n217 5.446
R23682 VSS.n1078 VSS.n222 5.446
R23683 VSS.n1078 VSS.n216 5.446
R23684 VSS.n1078 VSS.n1076 5.446
R23685 VSS.n988 VSS.n309 5.446
R23686 VSS.n988 VSS.n310 5.446
R23687 VSS.n988 VSS.n308 5.446
R23688 VSS.n988 VSS.n311 5.446
R23689 VSS.n988 VSS.n307 5.446
R23690 VSS.n988 VSS.n312 5.446
R23691 VSS.n988 VSS.n306 5.446
R23692 VSS.n988 VSS.n986 5.446
R23693 VSS.n898 VSS.n399 5.446
R23694 VSS.n898 VSS.n400 5.446
R23695 VSS.n898 VSS.n398 5.446
R23696 VSS.n898 VSS.n401 5.446
R23697 VSS.n898 VSS.n397 5.446
R23698 VSS.n898 VSS.n402 5.446
R23699 VSS.n898 VSS.n396 5.446
R23700 VSS.n898 VSS.n896 5.446
R23701 VSS.n808 VSS.n489 5.446
R23702 VSS.n808 VSS.n490 5.446
R23703 VSS.n808 VSS.n488 5.446
R23704 VSS.n808 VSS.n491 5.446
R23705 VSS.n808 VSS.n487 5.446
R23706 VSS.n808 VSS.n492 5.446
R23707 VSS.n808 VSS.n486 5.446
R23708 VSS.n808 VSS.n806 5.446
R23709 VSS.n718 VSS.n579 5.446
R23710 VSS.n718 VSS.n580 5.446
R23711 VSS.n718 VSS.n578 5.446
R23712 VSS.n718 VSS.n581 5.446
R23713 VSS.n718 VSS.n577 5.446
R23714 VSS.n718 VSS.n582 5.446
R23715 VSS.n718 VSS.n576 5.446
R23716 VSS.n718 VSS.n716 5.446
R23717 VSS.n17718 sky130_asc_pfet_01v8_lvt_12_0/VGND 5.433
R23718 VSS.n10464 VSS.n10426 5.341
R23719 VSS.n17680 VSS.n17679 5.341
R23720 VSS.n10467 VSS.n10426 5.233
R23721 VSS.n17679 VSS.n17678 5.233
R23722 VSS.n17703 VSS.n17702 5.079
R23723 VSS.n10486 VSS.n10418 5.007
R23724 VSS.n10449 VSS.n10448 4.894
R23725 VSS.n10474 VSS.n10473 4.894
R23726 VSS.n17671 VSS.n17670 4.894
R23727 VSS.n17691 VSS.n17646 4.894
R23728 sky130_asc_res_xhigh_po_2p85_2_0/Rout VSS.t4 4.868
R23729 sky130_asc_res_xhigh_po_2p85_2_1/Rout VSS.t7 4.868
R23730 VSS.n6606 VSS.t10 4.85
R23731 sky130_asc_pnp_05v5_W3p40L3p40_8_3/VGND sky130_asc_res_xhigh_po_2p85_1_22/VGND 4.846
R23732 VSS.n14369 VSS.n14367 4.792
R23733 VSS.n12792 VSS.n12720 4.792
R23734 VSS.n7676 VSS.n7671 4.792
R23735 VSS.n4245 VSS.n4173 4.792
R23736 VSS.n1610 VSS.n1608 4.792
R23737 VSS.n16002 VSS.n16001 4.65
R23738 VSS.n14375 VSS.n14368 4.65
R23739 VSS.n14711 VSS.n14374 4.65
R23740 VSS.n14701 VSS.n14700 4.65
R23741 VSS.n14387 VSS.n14384 4.65
R23742 VSS.n14688 VSS.n14394 4.65
R23743 VSS.n14678 VSS.n14677 4.65
R23744 VSS.n14406 VSS.n14403 4.65
R23745 VSS.n14666 VSS.n14413 4.65
R23746 VSS.n14656 VSS.n14655 4.65
R23747 VSS.n14425 VSS.n14422 4.65
R23748 VSS.n14643 VSS.n14432 4.65
R23749 VSS.n14633 VSS.n14632 4.65
R23750 VSS.n14477 VSS.n14475 4.65
R23751 VSS.n14619 VSS.n14487 4.65
R23752 VSS.n14609 VSS.n14608 4.65
R23753 VSS.n14499 VSS.n14496 4.65
R23754 VSS.n14596 VSS.n14506 4.65
R23755 VSS.n14586 VSS.n14585 4.65
R23756 VSS.n14518 VSS.n14515 4.65
R23757 VSS.n14574 VSS.n14525 4.65
R23758 VSS.n14564 VSS.n14563 4.65
R23759 VSS.n14537 VSS.n14534 4.65
R23760 VSS.n14551 VSS.n14548 4.65
R23761 VSS.n14868 VSS.n14306 4.65
R23762 VSS.n14880 VSS.n14297 4.65
R23763 VSS.n14890 VSS.n14291 4.65
R23764 VSS.n14286 VSS.n14285 4.65
R23765 VSS.n14904 VSS.n14284 4.65
R23766 VSS.n14915 VSS.n14276 4.65
R23767 VSS.n14925 VSS.n14270 4.65
R23768 VSS.n14265 VSS.n14264 4.65
R23769 VSS.n14938 VSS.n14263 4.65
R23770 VSS.n14949 VSS.n14255 4.65
R23771 VSS.n14959 VSS.n14249 4.65
R23772 VSS.n14244 VSS.n14243 4.65
R23773 VSS.n15326 VSS.n14242 4.65
R23774 VSS.n14975 VSS.n14973 4.65
R23775 VSS.n15312 VSS.n14984 4.65
R23776 VSS.n15302 VSS.n15301 4.65
R23777 VSS.n14996 VSS.n14993 4.65
R23778 VSS.n15289 VSS.n15003 4.65
R23779 VSS.n15279 VSS.n15278 4.65
R23780 VSS.n15015 VSS.n15012 4.65
R23781 VSS.n15267 VSS.n15022 4.65
R23782 VSS.n15257 VSS.n15256 4.65
R23783 VSS.n15034 VSS.n15031 4.65
R23784 VSS.n15244 VSS.n15041 4.65
R23785 VSS.n15234 VSS.n15233 4.65
R23786 VSS.n15086 VSS.n15084 4.65
R23787 VSS.n15220 VSS.n15096 4.65
R23788 VSS.n15210 VSS.n15209 4.65
R23789 VSS.n15108 VSS.n15105 4.65
R23790 VSS.n15197 VSS.n15115 4.65
R23791 VSS.n15187 VSS.n15186 4.65
R23792 VSS.n15127 VSS.n15124 4.65
R23793 VSS.n15175 VSS.n15134 4.65
R23794 VSS.n15165 VSS.n15164 4.65
R23795 VSS.n15146 VSS.n15143 4.65
R23796 VSS.n14139 VSS.n14138 4.65
R23797 VSS.n15452 VSS.n15451 4.65
R23798 VSS.n14130 VSS.n14129 4.65
R23799 VSS.n15467 VSS.n14128 4.65
R23800 VSS.n15478 VSS.n14120 4.65
R23801 VSS.n15488 VSS.n14114 4.65
R23802 VSS.n14109 VSS.n14108 4.65
R23803 VSS.n15502 VSS.n14107 4.65
R23804 VSS.n15512 VSS.n14099 4.65
R23805 VSS.n15522 VSS.n14093 4.65
R23806 VSS.n14088 VSS.n14087 4.65
R23807 VSS.n15536 VSS.n14086 4.65
R23808 VSS.n15547 VSS.n14078 4.65
R23809 VSS.n15558 VSS.n15557 4.65
R23810 VSS.n15562 VSS.n15560 4.65
R23811 VSS.n15879 VSS.n15571 4.65
R23812 VSS.n15869 VSS.n15868 4.65
R23813 VSS.n15583 VSS.n15580 4.65
R23814 VSS.n15856 VSS.n15590 4.65
R23815 VSS.n15846 VSS.n15845 4.65
R23816 VSS.n15602 VSS.n15599 4.65
R23817 VSS.n15834 VSS.n15609 4.65
R23818 VSS.n15824 VSS.n15823 4.65
R23819 VSS.n15621 VSS.n15618 4.65
R23820 VSS.n15811 VSS.n15628 4.65
R23821 VSS.n15801 VSS.n15800 4.65
R23822 VSS.n16012 VSS.n14005 4.65
R23823 VSS.n13998 VSS.n13996 4.65
R23824 VSS.n15732 VSS.n15731 4.65
R23825 VSS.n15742 VSS.n15721 4.65
R23826 VSS.n15714 VSS.n15711 4.65
R23827 VSS.n15754 VSS.n15753 4.65
R23828 VSS.n15764 VSS.n15702 4.65
R23829 VSS.n15695 VSS.n15692 4.65
R23830 VSS.n15777 VSS.n15776 4.65
R23831 VSS.n15787 VSS.n15683 4.65
R23832 VSS.n15673 VSS.n15671 4.65
R23833 VSS.n16714 VSS.n16712 4.65
R23834 VSS.n16719 VSS.n16709 4.65
R23835 VSS.n16724 VSS.n16706 4.65
R23836 VSS.n16730 VSS.n16702 4.65
R23837 VSS.n16736 VSS.n16698 4.65
R23838 VSS.n16742 VSS.n16692 4.65
R23839 VSS.n16748 VSS.n16747 4.65
R23840 VSS.n16756 VSS.n16632 4.65
R23841 VSS.n16688 VSS.n16687 4.65
R23842 VSS.n16770 VSS.n16769 4.65
R23843 VSS.n16804 VSS.n16802 4.65
R23844 VSS.n16809 VSS.n16799 4.65
R23845 VSS.n16814 VSS.n16796 4.65
R23846 VSS.n16820 VSS.n16792 4.65
R23847 VSS.n16826 VSS.n16788 4.65
R23848 VSS.n16832 VSS.n16782 4.65
R23849 VSS.n16838 VSS.n16837 4.65
R23850 VSS.n16846 VSS.n16542 4.65
R23851 VSS.n16778 VSS.n16777 4.65
R23852 VSS.n16860 VSS.n16859 4.65
R23853 VSS.n16894 VSS.n16892 4.65
R23854 VSS.n16899 VSS.n16889 4.65
R23855 VSS.n16904 VSS.n16886 4.65
R23856 VSS.n16910 VSS.n16882 4.65
R23857 VSS.n16916 VSS.n16878 4.65
R23858 VSS.n16922 VSS.n16872 4.65
R23859 VSS.n16928 VSS.n16927 4.65
R23860 VSS.n16936 VSS.n16452 4.65
R23861 VSS.n16868 VSS.n16867 4.65
R23862 VSS.n16950 VSS.n16949 4.65
R23863 VSS.n16984 VSS.n16982 4.65
R23864 VSS.n16989 VSS.n16979 4.65
R23865 VSS.n16994 VSS.n16976 4.65
R23866 VSS.n17000 VSS.n16972 4.65
R23867 VSS.n17006 VSS.n16968 4.65
R23868 VSS.n17012 VSS.n16962 4.65
R23869 VSS.n17018 VSS.n17017 4.65
R23870 VSS.n17026 VSS.n16362 4.65
R23871 VSS.n16958 VSS.n16957 4.65
R23872 VSS.n17040 VSS.n17039 4.65
R23873 VSS.n17074 VSS.n17072 4.65
R23874 VSS.n17079 VSS.n17069 4.65
R23875 VSS.n17084 VSS.n17066 4.65
R23876 VSS.n17090 VSS.n17062 4.65
R23877 VSS.n17096 VSS.n17058 4.65
R23878 VSS.n17102 VSS.n17052 4.65
R23879 VSS.n17108 VSS.n17107 4.65
R23880 VSS.n17116 VSS.n16272 4.65
R23881 VSS.n17048 VSS.n17047 4.65
R23882 VSS.n17130 VSS.n17129 4.65
R23883 VSS.n17164 VSS.n17162 4.65
R23884 VSS.n17169 VSS.n17159 4.65
R23885 VSS.n17174 VSS.n17156 4.65
R23886 VSS.n17180 VSS.n17152 4.65
R23887 VSS.n17186 VSS.n17148 4.65
R23888 VSS.n17192 VSS.n17142 4.65
R23889 VSS.n17198 VSS.n17197 4.65
R23890 VSS.n17206 VSS.n16182 4.65
R23891 VSS.n17138 VSS.n17137 4.65
R23892 VSS.n17220 VSS.n17219 4.65
R23893 VSS.n17254 VSS.n17252 4.65
R23894 VSS.n17259 VSS.n17249 4.65
R23895 VSS.n17264 VSS.n17246 4.65
R23896 VSS.n17270 VSS.n17242 4.65
R23897 VSS.n17276 VSS.n17238 4.65
R23898 VSS.n17282 VSS.n17232 4.65
R23899 VSS.n17288 VSS.n17287 4.65
R23900 VSS.n17296 VSS.n16092 4.65
R23901 VSS.n17228 VSS.n17227 4.65
R23902 VSS.n17310 VSS.n17309 4.65
R23903 VSS.n17334 VSS.n17333 4.65
R23904 VSS.n16028 VSS.n16026 4.65
R23905 VSS.n17426 VSS.n17411 4.65
R23906 VSS.n17432 VSS.n17407 4.65
R23907 VSS.n17438 VSS.n17401 4.65
R23908 VSS.n17444 VSS.n17443 4.65
R23909 VSS.n17452 VSS.n16049 4.65
R23910 VSS.n17397 VSS.n17396 4.65
R23911 VSS.n17389 VSS.n16051 4.65
R23912 VSS.n12217 VSS.n12216 4.65
R23913 VSS.n12800 VSS.n12718 4.65
R23914 VSS.n12713 VSS.n12712 4.65
R23915 VSS.n12814 VSS.n12711 4.65
R23916 VSS.n12825 VSS.n12703 4.65
R23917 VSS.n12835 VSS.n12697 4.65
R23918 VSS.n12692 VSS.n12691 4.65
R23919 VSS.n12849 VSS.n12690 4.65
R23920 VSS.n12859 VSS.n12682 4.65
R23921 VSS.n12869 VSS.n12676 4.65
R23922 VSS.n12669 VSS.n12668 4.65
R23923 VSS.n12886 VSS.n12885 4.65
R23924 VSS.n13062 VSS.n12660 4.65
R23925 VSS.n13050 VSS.n12894 4.65
R23926 VSS.n13040 VSS.n13039 4.65
R23927 VSS.n12905 VSS.n12902 4.65
R23928 VSS.n13027 VSS.n12912 4.65
R23929 VSS.n13017 VSS.n13016 4.65
R23930 VSS.n12924 VSS.n12921 4.65
R23931 VSS.n13005 VSS.n12931 4.65
R23932 VSS.n12995 VSS.n12994 4.65
R23933 VSS.n12943 VSS.n12940 4.65
R23934 VSS.n12982 VSS.n12950 4.65
R23935 VSS.n12972 VSS.n12971 4.65
R23936 VSS.n12963 VSS.n12960 4.65
R23937 VSS.n13157 VSS.n12577 4.65
R23938 VSS.n12572 VSS.n12571 4.65
R23939 VSS.n13171 VSS.n12570 4.65
R23940 VSS.n13182 VSS.n12562 4.65
R23941 VSS.n13192 VSS.n12556 4.65
R23942 VSS.n12551 VSS.n12550 4.65
R23943 VSS.n13206 VSS.n12549 4.65
R23944 VSS.n13216 VSS.n12541 4.65
R23945 VSS.n13226 VSS.n12535 4.65
R23946 VSS.n12528 VSS.n12527 4.65
R23947 VSS.n13243 VSS.n13242 4.65
R23948 VSS.n13311 VSS.n12519 4.65
R23949 VSS.n13299 VSS.n13251 4.65
R23950 VSS.n13289 VSS.n13288 4.65
R23951 VSS.n13262 VSS.n13259 4.65
R23952 VSS.n13276 VSS.n13273 4.65
R23953 VSS.n11432 VSS.n11430 4.65
R23954 VSS.n13446 VSS.n11439 4.65
R23955 VSS.n13437 VSS.n13436 4.65
R23956 VSS.n11451 VSS.n11448 4.65
R23957 VSS.n13424 VSS.n11458 4.65
R23958 VSS.n13414 VSS.n13413 4.65
R23959 VSS.n11470 VSS.n11467 4.65
R23960 VSS.n13401 VSS.n11477 4.65
R23961 VSS.n11678 VSS.n11668 4.65
R23962 VSS.n11663 VSS.n11662 4.65
R23963 VSS.n11692 VSS.n11661 4.65
R23964 VSS.n11703 VSS.n11653 4.65
R23965 VSS.n11713 VSS.n11647 4.65
R23966 VSS.n11642 VSS.n11641 4.65
R23967 VSS.n11727 VSS.n11640 4.65
R23968 VSS.n11737 VSS.n11632 4.65
R23969 VSS.n11747 VSS.n11626 4.65
R23970 VSS.n11621 VSS.n11620 4.65
R23971 VSS.n11761 VSS.n11619 4.65
R23972 VSS.n11772 VSS.n11610 4.65
R23973 VSS.n11814 VSS.n11602 4.65
R23974 VSS.n11824 VSS.n11596 4.65
R23975 VSS.n11591 VSS.n11590 4.65
R23976 VSS.n11838 VSS.n11589 4.65
R23977 VSS.n11849 VSS.n11581 4.65
R23978 VSS.n11859 VSS.n11575 4.65
R23979 VSS.n11570 VSS.n11569 4.65
R23980 VSS.n11872 VSS.n11568 4.65
R23981 VSS.n11883 VSS.n11560 4.65
R23982 VSS.n11893 VSS.n11554 4.65
R23983 VSS.n11549 VSS.n11548 4.65
R23984 VSS.n12401 VSS.n11547 4.65
R23985 VSS.n11909 VSS.n11907 4.65
R23986 VSS.n12387 VSS.n11918 4.65
R23987 VSS.n12377 VSS.n12376 4.65
R23988 VSS.n11930 VSS.n11927 4.65
R23989 VSS.n12364 VSS.n11937 4.65
R23990 VSS.n12354 VSS.n12353 4.65
R23991 VSS.n11949 VSS.n11946 4.65
R23992 VSS.n12342 VSS.n11956 4.65
R23993 VSS.n12332 VSS.n12331 4.65
R23994 VSS.n11968 VSS.n11965 4.65
R23995 VSS.n12319 VSS.n11975 4.65
R23996 VSS.n12309 VSS.n12308 4.65
R23997 VSS.n12227 VSS.n12054 4.65
R23998 VSS.n12047 VSS.n12044 4.65
R23999 VSS.n12240 VSS.n12239 4.65
R24000 VSS.n12250 VSS.n12035 4.65
R24001 VSS.n12028 VSS.n12025 4.65
R24002 VSS.n12262 VSS.n12261 4.65
R24003 VSS.n12272 VSS.n12016 4.65
R24004 VSS.n12009 VSS.n12006 4.65
R24005 VSS.n12285 VSS.n12284 4.65
R24006 VSS.n12295 VSS.n11997 4.65
R24007 VSS.n11987 VSS.n11985 4.65
R24008 VSS.n13897 VSS.n13896 4.65
R24009 VSS.n13944 VSS.n10516 4.65
R24010 VSS.n13936 VSS.n13935 4.65
R24011 VSS.n13930 VSS.n13901 4.65
R24012 VSS.n13924 VSS.n13907 4.65
R24013 VSS.n13918 VSS.n13911 4.65
R24014 VSS.n13831 VSS.n13830 4.65
R24015 VSS.n13834 VSS.n13833 4.65
R24016 VSS.n13752 VSS.n13748 4.65
R24017 VSS.n13763 VSS.n13742 4.65
R24018 VSS.n13768 VSS.n13739 4.65
R24019 VSS.n13774 VSS.n13735 4.65
R24020 VSS.n13780 VSS.n13729 4.65
R24021 VSS.n13786 VSS.n13785 4.65
R24022 VSS.n13794 VSS.n10559 4.65
R24023 VSS.n13662 VSS.n13658 4.65
R24024 VSS.n13673 VSS.n13652 4.65
R24025 VSS.n13678 VSS.n13649 4.65
R24026 VSS.n13684 VSS.n13645 4.65
R24027 VSS.n13690 VSS.n13639 4.65
R24028 VSS.n13696 VSS.n13695 4.65
R24029 VSS.n13704 VSS.n10649 4.65
R24030 VSS.n13572 VSS.n13568 4.65
R24031 VSS.n13583 VSS.n13562 4.65
R24032 VSS.n13588 VSS.n13559 4.65
R24033 VSS.n13594 VSS.n13555 4.65
R24034 VSS.n13600 VSS.n13549 4.65
R24035 VSS.n13606 VSS.n13605 4.65
R24036 VSS.n13614 VSS.n10739 4.65
R24037 VSS.n13481 VSS.n13477 4.65
R24038 VSS.n13492 VSS.n13471 4.65
R24039 VSS.n13497 VSS.n13468 4.65
R24040 VSS.n13503 VSS.n13464 4.65
R24041 VSS.n13509 VSS.n13458 4.65
R24042 VSS.n13516 VSS.n13515 4.65
R24043 VSS.n13524 VSS.n10829 4.65
R24044 VSS.n11362 VSS.n11358 4.65
R24045 VSS.n11373 VSS.n11352 4.65
R24046 VSS.n11378 VSS.n11349 4.65
R24047 VSS.n11384 VSS.n11345 4.65
R24048 VSS.n11390 VSS.n11339 4.65
R24049 VSS.n11396 VSS.n11395 4.65
R24050 VSS.n11404 VSS.n10919 4.65
R24051 VSS.n11272 VSS.n11268 4.65
R24052 VSS.n11283 VSS.n11262 4.65
R24053 VSS.n11288 VSS.n11259 4.65
R24054 VSS.n11294 VSS.n11255 4.65
R24055 VSS.n11300 VSS.n11249 4.65
R24056 VSS.n11306 VSS.n11305 4.65
R24057 VSS.n11314 VSS.n11009 4.65
R24058 VSS.n11182 VSS.n11178 4.65
R24059 VSS.n11193 VSS.n11172 4.65
R24060 VSS.n11198 VSS.n11169 4.65
R24061 VSS.n11204 VSS.n11165 4.65
R24062 VSS.n11210 VSS.n11159 4.65
R24063 VSS.n11216 VSS.n11215 4.65
R24064 VSS.n11224 VSS.n11099 4.65
R24065 VSS.n11155 VSS.n11154 4.65
R24066 VSS.n11187 VSS.n11175 4.65
R24067 VSS.n11237 VSS.n11236 4.65
R24068 VSS.n11245 VSS.n11244 4.65
R24069 VSS.n11277 VSS.n11265 4.65
R24070 VSS.n11327 VSS.n11326 4.65
R24071 VSS.n11335 VSS.n11334 4.65
R24072 VSS.n11367 VSS.n11355 4.65
R24073 VSS.n11417 VSS.n11416 4.65
R24074 VSS.n11425 VSS.n11424 4.65
R24075 VSS.n13486 VSS.n13474 4.65
R24076 VSS.n13537 VSS.n13536 4.65
R24077 VSS.n13545 VSS.n13544 4.65
R24078 VSS.n13577 VSS.n13565 4.65
R24079 VSS.n13627 VSS.n13626 4.65
R24080 VSS.n13635 VSS.n13634 4.65
R24081 VSS.n13667 VSS.n13655 4.65
R24082 VSS.n13717 VSS.n13716 4.65
R24083 VSS.n13725 VSS.n13724 4.65
R24084 VSS.n13757 VSS.n13745 4.65
R24085 VSS.n13807 VSS.n13806 4.65
R24086 VSS.n13889 VSS.n10518 4.65
R24087 VSS.n10465 VSS.n10464 4.65
R24088 VSS.n7174 VSS.n7006 4.65
R24089 VSS.n7682 VSS.n7675 4.65
R24090 VSS.n7825 VSS.n7681 4.65
R24091 VSS.n7815 VSS.n7814 4.65
R24092 VSS.n7694 VSS.n7691 4.65
R24093 VSS.n7802 VSS.n7701 4.65
R24094 VSS.n7792 VSS.n7791 4.65
R24095 VSS.n7713 VSS.n7710 4.65
R24096 VSS.n7780 VSS.n7720 4.65
R24097 VSS.n7770 VSS.n7769 4.65
R24098 VSS.n7732 VSS.n7729 4.65
R24099 VSS.n7757 VSS.n7739 4.65
R24100 VSS.n7747 VSS.n7746 4.65
R24101 VSS.n7925 VSS.n7596 4.65
R24102 VSS.n7935 VSS.n7590 4.65
R24103 VSS.n7585 VSS.n7584 4.65
R24104 VSS.n7949 VSS.n7583 4.65
R24105 VSS.n7960 VSS.n7575 4.65
R24106 VSS.n7970 VSS.n7569 4.65
R24107 VSS.n7564 VSS.n7563 4.65
R24108 VSS.n7983 VSS.n7562 4.65
R24109 VSS.n7994 VSS.n7554 4.65
R24110 VSS.n8004 VSS.n7548 4.65
R24111 VSS.n7543 VSS.n7542 4.65
R24112 VSS.n8187 VSS.n7541 4.65
R24113 VSS.n8028 VSS.n8027 4.65
R24114 VSS.n8036 VSS.n8024 4.65
R24115 VSS.n8165 VSS.n8035 4.65
R24116 VSS.n8155 VSS.n8154 4.65
R24117 VSS.n8048 VSS.n8045 4.65
R24118 VSS.n8142 VSS.n8055 4.65
R24119 VSS.n8133 VSS.n8132 4.65
R24120 VSS.n8067 VSS.n8064 4.65
R24121 VSS.n8120 VSS.n8074 4.65
R24122 VSS.n8110 VSS.n8109 4.65
R24123 VSS.n8086 VSS.n8083 4.65
R24124 VSS.n8097 VSS.n8092 4.65
R24125 VSS.n8283 VSS.n7456 4.65
R24126 VSS.n8293 VSS.n7450 4.65
R24127 VSS.n7445 VSS.n7444 4.65
R24128 VSS.n8307 VSS.n7443 4.65
R24129 VSS.n8318 VSS.n7435 4.65
R24130 VSS.n8328 VSS.n7429 4.65
R24131 VSS.n7424 VSS.n7423 4.65
R24132 VSS.n8341 VSS.n7422 4.65
R24133 VSS.n8352 VSS.n7414 4.65
R24134 VSS.n8362 VSS.n7408 4.65
R24135 VSS.n7403 VSS.n7402 4.65
R24136 VSS.n8545 VSS.n7401 4.65
R24137 VSS.n8386 VSS.n8385 4.65
R24138 VSS.n8394 VSS.n8382 4.65
R24139 VSS.n8523 VSS.n8393 4.65
R24140 VSS.n8513 VSS.n8512 4.65
R24141 VSS.n8406 VSS.n8403 4.65
R24142 VSS.n8500 VSS.n8413 4.65
R24143 VSS.n8491 VSS.n8490 4.65
R24144 VSS.n8425 VSS.n8422 4.65
R24145 VSS.n8478 VSS.n8432 4.65
R24146 VSS.n8468 VSS.n8467 4.65
R24147 VSS.n8444 VSS.n8441 4.65
R24148 VSS.n8455 VSS.n8450 4.65
R24149 VSS.n8641 VSS.n7316 4.65
R24150 VSS.n8651 VSS.n7310 4.65
R24151 VSS.n7305 VSS.n7304 4.65
R24152 VSS.n8665 VSS.n7303 4.65
R24153 VSS.n8676 VSS.n7295 4.65
R24154 VSS.n8686 VSS.n7289 4.65
R24155 VSS.n7284 VSS.n7283 4.65
R24156 VSS.n8699 VSS.n7282 4.65
R24157 VSS.n8710 VSS.n7274 4.65
R24158 VSS.n8720 VSS.n7268 4.65
R24159 VSS.n7263 VSS.n7262 4.65
R24160 VSS.n8767 VSS.n7261 4.65
R24161 VSS.n8744 VSS.n8743 4.65
R24162 VSS.n8746 VSS.n8740 4.65
R24163 VSS.n6904 VSS.n6902 4.65
R24164 VSS.n8918 VSS.n6911 4.65
R24165 VSS.n8908 VSS.n8907 4.65
R24166 VSS.n6923 VSS.n6920 4.65
R24167 VSS.n8896 VSS.n6930 4.65
R24168 VSS.n8886 VSS.n8885 4.65
R24169 VSS.n6942 VSS.n6939 4.65
R24170 VSS.n8873 VSS.n6949 4.65
R24171 VSS.n8863 VSS.n8862 4.65
R24172 VSS.n6961 VSS.n6958 4.65
R24173 VSS.n7163 VSS.n7013 4.65
R24174 VSS.n7152 VSS.n7021 4.65
R24175 VSS.n7023 VSS.n7022 4.65
R24176 VSS.n7138 VSS.n7028 4.65
R24177 VSS.n7128 VSS.n7034 4.65
R24178 VSS.n7118 VSS.n7042 4.65
R24179 VSS.n7044 VSS.n7043 4.65
R24180 VSS.n7104 VSS.n7049 4.65
R24181 VSS.n7094 VSS.n7055 4.65
R24182 VSS.n7083 VSS.n7063 4.65
R24183 VSS.n7065 VSS.n7064 4.65
R24184 VSS.n8933 VSS.n8931 4.65
R24185 VSS.n9759 VSS.n9757 4.65
R24186 VSS.n9764 VSS.n9754 4.65
R24187 VSS.n9769 VSS.n9751 4.65
R24188 VSS.n9775 VSS.n9747 4.65
R24189 VSS.n9781 VSS.n9743 4.65
R24190 VSS.n9787 VSS.n9737 4.65
R24191 VSS.n9793 VSS.n9792 4.65
R24192 VSS.n9801 VSS.n9677 4.65
R24193 VSS.n9733 VSS.n9732 4.65
R24194 VSS.n9815 VSS.n9814 4.65
R24195 VSS.n9849 VSS.n9847 4.65
R24196 VSS.n9854 VSS.n9844 4.65
R24197 VSS.n9859 VSS.n9841 4.65
R24198 VSS.n9865 VSS.n9837 4.65
R24199 VSS.n9871 VSS.n9833 4.65
R24200 VSS.n9877 VSS.n9827 4.65
R24201 VSS.n9883 VSS.n9882 4.65
R24202 VSS.n9891 VSS.n9587 4.65
R24203 VSS.n9823 VSS.n9822 4.65
R24204 VSS.n9905 VSS.n9904 4.65
R24205 VSS.n9939 VSS.n9937 4.65
R24206 VSS.n9944 VSS.n9934 4.65
R24207 VSS.n9949 VSS.n9931 4.65
R24208 VSS.n9955 VSS.n9927 4.65
R24209 VSS.n9961 VSS.n9923 4.65
R24210 VSS.n9967 VSS.n9917 4.65
R24211 VSS.n9973 VSS.n9972 4.65
R24212 VSS.n9981 VSS.n9497 4.65
R24213 VSS.n9913 VSS.n9912 4.65
R24214 VSS.n9995 VSS.n9994 4.65
R24215 VSS.n10029 VSS.n10027 4.65
R24216 VSS.n10034 VSS.n10024 4.65
R24217 VSS.n10039 VSS.n10021 4.65
R24218 VSS.n10045 VSS.n10017 4.65
R24219 VSS.n10051 VSS.n10013 4.65
R24220 VSS.n10057 VSS.n10007 4.65
R24221 VSS.n10063 VSS.n10062 4.65
R24222 VSS.n10071 VSS.n9407 4.65
R24223 VSS.n10003 VSS.n10002 4.65
R24224 VSS.n10085 VSS.n10084 4.65
R24225 VSS.n10119 VSS.n10117 4.65
R24226 VSS.n10124 VSS.n10114 4.65
R24227 VSS.n10129 VSS.n10111 4.65
R24228 VSS.n10135 VSS.n10107 4.65
R24229 VSS.n10141 VSS.n10103 4.65
R24230 VSS.n10147 VSS.n10097 4.65
R24231 VSS.n10153 VSS.n10152 4.65
R24232 VSS.n10161 VSS.n9317 4.65
R24233 VSS.n10093 VSS.n10092 4.65
R24234 VSS.n10175 VSS.n10174 4.65
R24235 VSS.n10209 VSS.n10207 4.65
R24236 VSS.n10214 VSS.n10204 4.65
R24237 VSS.n10219 VSS.n10201 4.65
R24238 VSS.n10225 VSS.n10197 4.65
R24239 VSS.n10231 VSS.n10193 4.65
R24240 VSS.n10237 VSS.n10187 4.65
R24241 VSS.n10243 VSS.n10242 4.65
R24242 VSS.n10251 VSS.n9227 4.65
R24243 VSS.n10183 VSS.n10182 4.65
R24244 VSS.n10265 VSS.n10264 4.65
R24245 VSS.n9036 VSS.n9033 4.65
R24246 VSS.n9044 VSS.n9031 4.65
R24247 VSS.n9052 VSS.n9029 4.65
R24248 VSS.n9060 VSS.n9027 4.65
R24249 VSS.n9068 VSS.n9025 4.65
R24250 VSS.n9076 VSS.n9023 4.65
R24251 VSS.n9084 VSS.n9021 4.65
R24252 VSS.n9092 VSS.n9019 4.65
R24253 VSS.n9151 VSS.n9018 4.65
R24254 VSS.n9148 VSS.n9097 4.65
R24255 VSS.n9162 VSS.n9161 4.65
R24256 VSS.n8979 VSS.n8973 4.65
R24257 VSS.n8974 VSS.n8967 4.65
R24258 VSS.n8968 VSS.n8960 4.65
R24259 VSS.n8962 VSS.n8961 4.65
R24260 VSS.n8955 VSS.n8949 4.65
R24261 VSS.n8950 VSS.n8943 4.65
R24262 VSS.n8944 VSS.n8938 4.65
R24263 VSS.n10319 VSS.n9186 4.65
R24264 VSS.n6881 VSS.n6880 4.65
R24265 VSS.n3638 VSS.n3636 4.65
R24266 VSS.n4253 VSS.n4171 4.65
R24267 VSS.n4166 VSS.n4165 4.65
R24268 VSS.n4267 VSS.n4164 4.65
R24269 VSS.n4278 VSS.n4156 4.65
R24270 VSS.n4288 VSS.n4150 4.65
R24271 VSS.n4145 VSS.n4144 4.65
R24272 VSS.n4302 VSS.n4143 4.65
R24273 VSS.n4312 VSS.n4135 4.65
R24274 VSS.n4322 VSS.n4129 4.65
R24275 VSS.n4122 VSS.n4121 4.65
R24276 VSS.n4339 VSS.n4338 4.65
R24277 VSS.n4515 VSS.n4113 4.65
R24278 VSS.n4503 VSS.n4347 4.65
R24279 VSS.n4493 VSS.n4492 4.65
R24280 VSS.n4358 VSS.n4355 4.65
R24281 VSS.n4480 VSS.n4365 4.65
R24282 VSS.n4470 VSS.n4469 4.65
R24283 VSS.n4377 VSS.n4374 4.65
R24284 VSS.n4458 VSS.n4384 4.65
R24285 VSS.n4448 VSS.n4447 4.65
R24286 VSS.n4396 VSS.n4393 4.65
R24287 VSS.n4435 VSS.n4403 4.65
R24288 VSS.n4425 VSS.n4424 4.65
R24289 VSS.n4416 VSS.n4413 4.65
R24290 VSS.n4610 VSS.n4030 4.65
R24291 VSS.n4025 VSS.n4024 4.65
R24292 VSS.n4624 VSS.n4023 4.65
R24293 VSS.n4635 VSS.n4015 4.65
R24294 VSS.n4645 VSS.n4009 4.65
R24295 VSS.n4004 VSS.n4003 4.65
R24296 VSS.n4659 VSS.n4002 4.65
R24297 VSS.n4669 VSS.n3994 4.65
R24298 VSS.n4679 VSS.n3988 4.65
R24299 VSS.n3981 VSS.n3980 4.65
R24300 VSS.n4696 VSS.n4695 4.65
R24301 VSS.n4872 VSS.n3972 4.65
R24302 VSS.n4860 VSS.n4704 4.65
R24303 VSS.n4850 VSS.n4849 4.65
R24304 VSS.n4715 VSS.n4712 4.65
R24305 VSS.n4837 VSS.n4722 4.65
R24306 VSS.n4827 VSS.n4826 4.65
R24307 VSS.n4734 VSS.n4731 4.65
R24308 VSS.n4815 VSS.n4741 4.65
R24309 VSS.n4805 VSS.n4804 4.65
R24310 VSS.n4753 VSS.n4750 4.65
R24311 VSS.n4792 VSS.n4760 4.65
R24312 VSS.n4782 VSS.n4781 4.65
R24313 VSS.n4773 VSS.n4770 4.65
R24314 VSS.n4967 VSS.n3889 4.65
R24315 VSS.n3884 VSS.n3883 4.65
R24316 VSS.n4981 VSS.n3882 4.65
R24317 VSS.n4992 VSS.n3874 4.65
R24318 VSS.n5002 VSS.n3868 4.65
R24319 VSS.n3863 VSS.n3862 4.65
R24320 VSS.n5016 VSS.n3861 4.65
R24321 VSS.n5026 VSS.n3853 4.65
R24322 VSS.n5036 VSS.n3847 4.65
R24323 VSS.n3840 VSS.n3839 4.65
R24324 VSS.n5053 VSS.n5052 4.65
R24325 VSS.n5229 VSS.n3831 4.65
R24326 VSS.n5217 VSS.n5061 4.65
R24327 VSS.n5207 VSS.n5206 4.65
R24328 VSS.n5072 VSS.n5069 4.65
R24329 VSS.n5194 VSS.n5079 4.65
R24330 VSS.n5184 VSS.n5183 4.65
R24331 VSS.n5091 VSS.n5088 4.65
R24332 VSS.n5172 VSS.n5098 4.65
R24333 VSS.n5162 VSS.n5161 4.65
R24334 VSS.n5110 VSS.n5107 4.65
R24335 VSS.n5149 VSS.n5117 4.65
R24336 VSS.n5139 VSS.n5138 4.65
R24337 VSS.n5130 VSS.n5127 4.65
R24338 VSS.n5324 VSS.n3748 4.65
R24339 VSS.n3743 VSS.n3742 4.65
R24340 VSS.n5338 VSS.n3741 4.65
R24341 VSS.n5349 VSS.n3733 4.65
R24342 VSS.n5359 VSS.n3727 4.65
R24343 VSS.n3722 VSS.n3721 4.65
R24344 VSS.n5373 VSS.n3720 4.65
R24345 VSS.n5383 VSS.n3712 4.65
R24346 VSS.n5393 VSS.n3706 4.65
R24347 VSS.n3699 VSS.n3698 4.65
R24348 VSS.n5410 VSS.n5409 4.65
R24349 VSS.n5575 VSS.n3690 4.65
R24350 VSS.n5485 VSS.n5484 4.65
R24351 VSS.n5495 VSS.n5474 4.65
R24352 VSS.n5467 VSS.n5464 4.65
R24353 VSS.n5508 VSS.n5507 4.65
R24354 VSS.n5518 VSS.n5455 4.65
R24355 VSS.n5448 VSS.n5445 4.65
R24356 VSS.n5530 VSS.n5529 4.65
R24357 VSS.n5540 VSS.n5436 4.65
R24358 VSS.n5429 VSS.n5426 4.65
R24359 VSS.n5553 VSS.n5552 4.65
R24360 VSS.n5563 VSS.n5418 4.65
R24361 VSS.n6593 VSS.n3160 4.65
R24362 VSS.n3224 VSS.n3161 4.65
R24363 VSS.n3216 VSS.n3163 4.65
R24364 VSS.n3208 VSS.n3165 4.65
R24365 VSS.n3200 VSS.n3167 4.65
R24366 VSS.n3192 VSS.n3169 4.65
R24367 VSS.n3184 VSS.n3171 4.65
R24368 VSS.n3176 VSS.n3173 4.65
R24369 VSS.n6604 VSS.n6603 4.65
R24370 VSS.n6590 VSS.n6519 4.65
R24371 VSS.n3285 VSS.n3278 4.65
R24372 VSS.n3279 VSS.n3272 4.65
R24373 VSS.n3273 VSS.n3265 4.65
R24374 VSS.n3267 VSS.n3266 4.65
R24375 VSS.n3260 VSS.n3254 4.65
R24376 VSS.n3255 VSS.n3248 4.65
R24377 VSS.n3249 VSS.n3242 4.65
R24378 VSS.n3243 VSS.n3237 4.65
R24379 VSS.n3232 VSS.n3230 4.65
R24380 VSS.n6398 VSS.n6397 4.65
R24381 VSS.n3343 VSS.n3336 4.65
R24382 VSS.n3337 VSS.n3330 4.65
R24383 VSS.n3331 VSS.n3323 4.65
R24384 VSS.n3325 VSS.n3324 4.65
R24385 VSS.n3318 VSS.n3312 4.65
R24386 VSS.n3313 VSS.n3306 4.65
R24387 VSS.n3307 VSS.n3300 4.65
R24388 VSS.n3301 VSS.n3295 4.65
R24389 VSS.n3290 VSS.n3288 4.65
R24390 VSS.n6276 VSS.n6275 4.65
R24391 VSS.n3401 VSS.n3394 4.65
R24392 VSS.n3395 VSS.n3388 4.65
R24393 VSS.n3389 VSS.n3381 4.65
R24394 VSS.n3383 VSS.n3382 4.65
R24395 VSS.n3376 VSS.n3370 4.65
R24396 VSS.n3371 VSS.n3364 4.65
R24397 VSS.n3365 VSS.n3358 4.65
R24398 VSS.n3359 VSS.n3353 4.65
R24399 VSS.n3348 VSS.n3346 4.65
R24400 VSS.n6154 VSS.n6153 4.65
R24401 VSS.n3459 VSS.n3452 4.65
R24402 VSS.n3453 VSS.n3446 4.65
R24403 VSS.n3447 VSS.n3439 4.65
R24404 VSS.n3441 VSS.n3440 4.65
R24405 VSS.n3434 VSS.n3428 4.65
R24406 VSS.n3429 VSS.n3422 4.65
R24407 VSS.n3423 VSS.n3416 4.65
R24408 VSS.n3417 VSS.n3411 4.65
R24409 VSS.n3406 VSS.n3404 4.65
R24410 VSS.n6032 VSS.n6031 4.65
R24411 VSS.n3517 VSS.n3510 4.65
R24412 VSS.n3511 VSS.n3504 4.65
R24413 VSS.n3505 VSS.n3497 4.65
R24414 VSS.n3499 VSS.n3498 4.65
R24415 VSS.n3492 VSS.n3486 4.65
R24416 VSS.n3487 VSS.n3480 4.65
R24417 VSS.n3481 VSS.n3474 4.65
R24418 VSS.n3475 VSS.n3469 4.65
R24419 VSS.n3464 VSS.n3462 4.65
R24420 VSS.n5910 VSS.n5909 4.65
R24421 VSS.n3575 VSS.n3568 4.65
R24422 VSS.n3569 VSS.n3562 4.65
R24423 VSS.n3563 VSS.n3555 4.65
R24424 VSS.n3557 VSS.n3556 4.65
R24425 VSS.n3550 VSS.n3544 4.65
R24426 VSS.n3545 VSS.n3538 4.65
R24427 VSS.n3539 VSS.n3532 4.65
R24428 VSS.n3533 VSS.n3527 4.65
R24429 VSS.n3522 VSS.n3520 4.65
R24430 VSS.n5788 VSS.n5787 4.65
R24431 VSS.n3633 VSS.n3626 4.65
R24432 VSS.n3627 VSS.n3620 4.65
R24433 VSS.n3621 VSS.n3613 4.65
R24434 VSS.n3615 VSS.n3614 4.65
R24435 VSS.n3608 VSS.n3602 4.65
R24436 VSS.n3603 VSS.n3596 4.65
R24437 VSS.n3597 VSS.n3590 4.65
R24438 VSS.n3591 VSS.n3585 4.65
R24439 VSS.n3580 VSS.n3578 4.65
R24440 VSS.n5666 VSS.n5665 4.65
R24441 VSS.n2875 VSS.n2874 4.65
R24442 VSS.n1616 VSS.n1609 4.65
R24443 VSS.n1952 VSS.n1615 4.65
R24444 VSS.n1942 VSS.n1941 4.65
R24445 VSS.n1628 VSS.n1625 4.65
R24446 VSS.n1929 VSS.n1635 4.65
R24447 VSS.n1919 VSS.n1918 4.65
R24448 VSS.n1647 VSS.n1644 4.65
R24449 VSS.n1907 VSS.n1654 4.65
R24450 VSS.n1897 VSS.n1896 4.65
R24451 VSS.n1666 VSS.n1663 4.65
R24452 VSS.n1884 VSS.n1673 4.65
R24453 VSS.n1874 VSS.n1873 4.65
R24454 VSS.n1718 VSS.n1716 4.65
R24455 VSS.n1860 VSS.n1728 4.65
R24456 VSS.n1850 VSS.n1849 4.65
R24457 VSS.n1740 VSS.n1737 4.65
R24458 VSS.n1837 VSS.n1747 4.65
R24459 VSS.n1827 VSS.n1826 4.65
R24460 VSS.n1759 VSS.n1756 4.65
R24461 VSS.n1815 VSS.n1766 4.65
R24462 VSS.n1805 VSS.n1804 4.65
R24463 VSS.n1778 VSS.n1775 4.65
R24464 VSS.n1792 VSS.n1789 4.65
R24465 VSS.n2109 VSS.n1547 4.65
R24466 VSS.n2121 VSS.n1538 4.65
R24467 VSS.n2131 VSS.n1532 4.65
R24468 VSS.n1527 VSS.n1526 4.65
R24469 VSS.n2145 VSS.n1525 4.65
R24470 VSS.n2156 VSS.n1517 4.65
R24471 VSS.n2166 VSS.n1511 4.65
R24472 VSS.n1506 VSS.n1505 4.65
R24473 VSS.n2179 VSS.n1504 4.65
R24474 VSS.n2190 VSS.n1496 4.65
R24475 VSS.n2200 VSS.n1490 4.65
R24476 VSS.n1485 VSS.n1484 4.65
R24477 VSS.n2567 VSS.n1483 4.65
R24478 VSS.n2216 VSS.n2214 4.65
R24479 VSS.n2553 VSS.n2225 4.65
R24480 VSS.n2543 VSS.n2542 4.65
R24481 VSS.n2237 VSS.n2234 4.65
R24482 VSS.n2530 VSS.n2244 4.65
R24483 VSS.n2520 VSS.n2519 4.65
R24484 VSS.n2256 VSS.n2253 4.65
R24485 VSS.n2508 VSS.n2263 4.65
R24486 VSS.n2498 VSS.n2497 4.65
R24487 VSS.n2275 VSS.n2272 4.65
R24488 VSS.n2485 VSS.n2282 4.65
R24489 VSS.n2475 VSS.n2474 4.65
R24490 VSS.n2327 VSS.n2325 4.65
R24491 VSS.n2461 VSS.n2337 4.65
R24492 VSS.n2451 VSS.n2450 4.65
R24493 VSS.n2349 VSS.n2346 4.65
R24494 VSS.n2438 VSS.n2356 4.65
R24495 VSS.n2428 VSS.n2427 4.65
R24496 VSS.n2368 VSS.n2365 4.65
R24497 VSS.n2416 VSS.n2375 4.65
R24498 VSS.n2406 VSS.n2405 4.65
R24499 VSS.n2387 VSS.n2384 4.65
R24500 VSS.n1380 VSS.n1379 4.65
R24501 VSS.n2693 VSS.n2692 4.65
R24502 VSS.n1371 VSS.n1370 4.65
R24503 VSS.n2708 VSS.n1369 4.65
R24504 VSS.n2719 VSS.n1361 4.65
R24505 VSS.n2729 VSS.n1355 4.65
R24506 VSS.n1350 VSS.n1349 4.65
R24507 VSS.n2743 VSS.n1348 4.65
R24508 VSS.n2753 VSS.n1340 4.65
R24509 VSS.n2763 VSS.n1334 4.65
R24510 VSS.n1329 VSS.n1328 4.65
R24511 VSS.n2777 VSS.n1327 4.65
R24512 VSS.n2788 VSS.n1319 4.65
R24513 VSS.n2799 VSS.n2798 4.65
R24514 VSS.n2885 VSS.n2869 4.65
R24515 VSS.n2862 VSS.n2859 4.65
R24516 VSS.n2898 VSS.n2897 4.65
R24517 VSS.n2908 VSS.n2850 4.65
R24518 VSS.n2843 VSS.n2840 4.65
R24519 VSS.n2920 VSS.n2919 4.65
R24520 VSS.n2930 VSS.n2831 4.65
R24521 VSS.n2824 VSS.n2821 4.65
R24522 VSS.n2943 VSS.n2942 4.65
R24523 VSS.n2953 VSS.n2812 4.65
R24524 VSS.n2803 VSS.n2801 4.65
R24525 VSS.n667 VSS.n665 4.65
R24526 VSS.n672 VSS.n662 4.65
R24527 VSS.n677 VSS.n659 4.65
R24528 VSS.n683 VSS.n655 4.65
R24529 VSS.n689 VSS.n651 4.65
R24530 VSS.n695 VSS.n645 4.65
R24531 VSS.n701 VSS.n700 4.65
R24532 VSS.n709 VSS.n585 4.65
R24533 VSS.n641 VSS.n640 4.65
R24534 VSS.n723 VSS.n722 4.65
R24535 VSS.n757 VSS.n755 4.65
R24536 VSS.n762 VSS.n752 4.65
R24537 VSS.n767 VSS.n749 4.65
R24538 VSS.n773 VSS.n745 4.65
R24539 VSS.n779 VSS.n741 4.65
R24540 VSS.n785 VSS.n735 4.65
R24541 VSS.n791 VSS.n790 4.65
R24542 VSS.n799 VSS.n495 4.65
R24543 VSS.n731 VSS.n730 4.65
R24544 VSS.n813 VSS.n812 4.65
R24545 VSS.n847 VSS.n845 4.65
R24546 VSS.n852 VSS.n842 4.65
R24547 VSS.n857 VSS.n839 4.65
R24548 VSS.n863 VSS.n835 4.65
R24549 VSS.n869 VSS.n831 4.65
R24550 VSS.n875 VSS.n825 4.65
R24551 VSS.n881 VSS.n880 4.65
R24552 VSS.n889 VSS.n405 4.65
R24553 VSS.n821 VSS.n820 4.65
R24554 VSS.n903 VSS.n902 4.65
R24555 VSS.n937 VSS.n935 4.65
R24556 VSS.n942 VSS.n932 4.65
R24557 VSS.n947 VSS.n929 4.65
R24558 VSS.n953 VSS.n925 4.65
R24559 VSS.n959 VSS.n921 4.65
R24560 VSS.n965 VSS.n915 4.65
R24561 VSS.n971 VSS.n970 4.65
R24562 VSS.n979 VSS.n315 4.65
R24563 VSS.n911 VSS.n910 4.65
R24564 VSS.n993 VSS.n992 4.65
R24565 VSS.n1027 VSS.n1025 4.65
R24566 VSS.n1032 VSS.n1022 4.65
R24567 VSS.n1037 VSS.n1019 4.65
R24568 VSS.n1043 VSS.n1015 4.65
R24569 VSS.n1049 VSS.n1011 4.65
R24570 VSS.n1055 VSS.n1005 4.65
R24571 VSS.n1061 VSS.n1060 4.65
R24572 VSS.n1069 VSS.n225 4.65
R24573 VSS.n1001 VSS.n1000 4.65
R24574 VSS.n1083 VSS.n1082 4.65
R24575 VSS.n1117 VSS.n1115 4.65
R24576 VSS.n1122 VSS.n1112 4.65
R24577 VSS.n1127 VSS.n1109 4.65
R24578 VSS.n1133 VSS.n1105 4.65
R24579 VSS.n1139 VSS.n1101 4.65
R24580 VSS.n1145 VSS.n1095 4.65
R24581 VSS.n1151 VSS.n1150 4.65
R24582 VSS.n1159 VSS.n135 4.65
R24583 VSS.n1091 VSS.n1090 4.65
R24584 VSS.n1173 VSS.n1172 4.65
R24585 VSS.n1258 VSS.n1257 4.65
R24586 VSS.n1207 VSS.n1202 4.65
R24587 VSS.n1212 VSS.n1199 4.65
R24588 VSS.n1218 VSS.n1195 4.65
R24589 VSS.n1224 VSS.n1191 4.65
R24590 VSS.n1230 VSS.n1185 4.65
R24591 VSS.n1236 VSS.n1235 4.65
R24592 VSS.n1244 VSS.n44 4.65
R24593 VSS.n1181 VSS.n1180 4.65
R24594 VSS.n1262 VSS.n2 4.65
R24595 VSS.n17681 VSS.n17680 4.65
R24596 VSS.n15669 VSS.n15637 4.608
R24597 VSS.n15663 VSS.n15637 4.608
R24598 VSS.n15663 VSS.n15662 4.608
R24599 VSS.n15662 VSS.n15661 4.608
R24600 VSS.n15661 VSS.n15641 4.608
R24601 VSS.n15655 VSS.n15641 4.608
R24602 VSS.n15655 VSS.n15654 4.608
R24603 VSS.n15654 VSS.n15653 4.608
R24604 VSS.n15653 VSS.n15645 4.608
R24605 VSS.n15647 VSS.n15645 4.608
R24606 VSS.n15647 VSS.n14040 4.608
R24607 VSS.n15948 VSS.n14040 4.608
R24608 VSS.n15892 VSS.n14067 4.608
R24609 VSS.n15898 VSS.n14067 4.608
R24610 VSS.n15899 VSS.n15898 4.608
R24611 VSS.n15900 VSS.n15899 4.608
R24612 VSS.n15900 VSS.n14063 4.608
R24613 VSS.n15906 VSS.n14063 4.608
R24614 VSS.n15907 VSS.n15906 4.608
R24615 VSS.n15908 VSS.n15907 4.608
R24616 VSS.n15908 VSS.n14059 4.608
R24617 VSS.n15914 VSS.n14059 4.608
R24618 VSS.n15915 VSS.n15914 4.608
R24619 VSS.n15916 VSS.n15915 4.608
R24620 VSS.n14148 VSS.n14136 4.608
R24621 VSS.n15435 VSS.n14148 4.608
R24622 VSS.n15435 VSS.n15434 4.608
R24623 VSS.n15434 VSS.n15433 4.608
R24624 VSS.n15433 VSS.n14149 4.608
R24625 VSS.n15427 VSS.n14149 4.608
R24626 VSS.n15427 VSS.n15426 4.608
R24627 VSS.n15426 VSS.n15425 4.608
R24628 VSS.n15425 VSS.n14153 4.608
R24629 VSS.n15419 VSS.n14153 4.608
R24630 VSS.n15419 VSS.n15418 4.608
R24631 VSS.n15418 VSS.n15417 4.608
R24632 VSS.n15082 VSS.n15050 4.608
R24633 VSS.n15076 VSS.n15050 4.608
R24634 VSS.n15076 VSS.n15075 4.608
R24635 VSS.n15075 VSS.n15074 4.608
R24636 VSS.n15074 VSS.n15054 4.608
R24637 VSS.n15068 VSS.n15054 4.608
R24638 VSS.n15068 VSS.n15067 4.608
R24639 VSS.n15067 VSS.n15066 4.608
R24640 VSS.n15066 VSS.n15058 4.608
R24641 VSS.n15060 VSS.n15058 4.608
R24642 VSS.n15060 VSS.n14210 4.608
R24643 VSS.n15386 VSS.n14210 4.608
R24644 VSS.n15335 VSS.n15334 4.608
R24645 VSS.n15336 VSS.n15335 4.608
R24646 VSS.n15336 VSS.n14232 4.608
R24647 VSS.n15342 VSS.n14232 4.608
R24648 VSS.n15343 VSS.n15342 4.608
R24649 VSS.n15344 VSS.n15343 4.608
R24650 VSS.n15344 VSS.n14228 4.608
R24651 VSS.n15350 VSS.n14228 4.608
R24652 VSS.n15351 VSS.n15350 4.608
R24653 VSS.n15352 VSS.n15351 4.608
R24654 VSS.n15352 VSS.n14224 4.608
R24655 VSS.n15358 VSS.n14224 4.608
R24656 VSS.n14864 VSS.n14308 4.608
R24657 VSS.n14312 VSS.n14308 4.608
R24658 VSS.n14857 VSS.n14312 4.608
R24659 VSS.n14857 VSS.n14856 4.608
R24660 VSS.n14856 VSS.n14855 4.608
R24661 VSS.n14855 VSS.n14313 4.608
R24662 VSS.n14849 VSS.n14313 4.608
R24663 VSS.n14849 VSS.n14848 4.608
R24664 VSS.n14848 VSS.n14847 4.608
R24665 VSS.n14847 VSS.n14317 4.608
R24666 VSS.n14841 VSS.n14317 4.608
R24667 VSS.n14841 VSS.n14840 4.608
R24668 VSS.n14473 VSS.n14441 4.608
R24669 VSS.n14467 VSS.n14441 4.608
R24670 VSS.n14467 VSS.n14466 4.608
R24671 VSS.n14466 VSS.n14465 4.608
R24672 VSS.n14465 VSS.n14445 4.608
R24673 VSS.n14459 VSS.n14445 4.608
R24674 VSS.n14459 VSS.n14458 4.608
R24675 VSS.n14458 VSS.n14457 4.608
R24676 VSS.n14457 VSS.n14449 4.608
R24677 VSS.n14451 VSS.n14449 4.608
R24678 VSS.n14451 VSS.n14336 4.608
R24679 VSS.n14778 VSS.n14336 4.608
R24680 VSS.n12105 VSS.n12104 4.608
R24681 VSS.n12106 VSS.n12105 4.608
R24682 VSS.n12106 VSS.n12098 4.608
R24683 VSS.n12112 VSS.n12098 4.608
R24684 VSS.n12113 VSS.n12112 4.608
R24685 VSS.n12114 VSS.n12113 4.608
R24686 VSS.n12114 VSS.n12094 4.608
R24687 VSS.n12120 VSS.n12094 4.608
R24688 VSS.n12121 VSS.n12120 4.608
R24689 VSS.n12122 VSS.n12121 4.608
R24690 VSS.n12122 VSS.n12089 4.608
R24691 VSS.n12163 VSS.n12089 4.608
R24692 VSS.n12410 VSS.n12409 4.608
R24693 VSS.n12411 VSS.n12410 4.608
R24694 VSS.n12411 VSS.n11537 4.608
R24695 VSS.n12417 VSS.n11537 4.608
R24696 VSS.n12418 VSS.n12417 4.608
R24697 VSS.n12419 VSS.n12418 4.608
R24698 VSS.n12419 VSS.n11533 4.608
R24699 VSS.n12425 VSS.n11533 4.608
R24700 VSS.n12426 VSS.n12425 4.608
R24701 VSS.n12427 VSS.n12426 4.608
R24702 VSS.n12427 VSS.n11529 4.608
R24703 VSS.n12433 VSS.n11529 4.608
R24704 VSS.n11804 VSS.n11803 4.608
R24705 VSS.n11803 VSS.n11802 4.608
R24706 VSS.n11802 VSS.n11776 4.608
R24707 VSS.n11796 VSS.n11776 4.608
R24708 VSS.n11796 VSS.n11795 4.608
R24709 VSS.n11795 VSS.n11794 4.608
R24710 VSS.n11794 VSS.n11780 4.608
R24711 VSS.n11788 VSS.n11780 4.608
R24712 VSS.n11788 VSS.n11787 4.608
R24713 VSS.n11787 VSS.n11786 4.608
R24714 VSS.n11786 VSS.n11514 4.608
R24715 VSS.n12460 VSS.n11514 4.608
R24716 VSS.n13397 VSS.n11482 4.608
R24717 VSS.n13391 VSS.n11482 4.608
R24718 VSS.n13391 VSS.n13390 4.608
R24719 VSS.n13390 VSS.n13389 4.608
R24720 VSS.n13389 VSS.n11488 4.608
R24721 VSS.n13383 VSS.n11488 4.608
R24722 VSS.n13383 VSS.n13382 4.608
R24723 VSS.n13382 VSS.n13381 4.608
R24724 VSS.n13381 VSS.n11492 4.608
R24725 VSS.n13375 VSS.n11492 4.608
R24726 VSS.n13375 VSS.n13374 4.608
R24727 VSS.n13374 VSS.n13373 4.608
R24728 VSS.n13316 VSS.n13315 4.608
R24729 VSS.n13316 VSS.n12513 4.608
R24730 VSS.n13322 VSS.n12513 4.608
R24731 VSS.n13323 VSS.n13322 4.608
R24732 VSS.n13324 VSS.n13323 4.608
R24733 VSS.n13324 VSS.n12509 4.608
R24734 VSS.n13330 VSS.n12509 4.608
R24735 VSS.n13331 VSS.n13330 4.608
R24736 VSS.n13333 VSS.n13331 4.608
R24737 VSS.n13333 VSS.n13332 4.608
R24738 VSS.n13332 VSS.n12505 4.608
R24739 VSS.n13340 VSS.n12505 4.608
R24740 VSS.n13148 VSS.n12585 4.608
R24741 VSS.n13142 VSS.n12585 4.608
R24742 VSS.n13142 VSS.n13141 4.608
R24743 VSS.n13141 VSS.n13140 4.608
R24744 VSS.n13140 VSS.n12589 4.608
R24745 VSS.n13134 VSS.n12589 4.608
R24746 VSS.n13134 VSS.n13133 4.608
R24747 VSS.n13133 VSS.n13132 4.608
R24748 VSS.n13132 VSS.n12593 4.608
R24749 VSS.n13126 VSS.n12593 4.608
R24750 VSS.n13126 VSS.n13125 4.608
R24751 VSS.n13125 VSS.n13124 4.608
R24752 VSS.n13067 VSS.n13066 4.608
R24753 VSS.n13067 VSS.n12654 4.608
R24754 VSS.n13073 VSS.n12654 4.608
R24755 VSS.n13074 VSS.n13073 4.608
R24756 VSS.n13075 VSS.n13074 4.608
R24757 VSS.n13075 VSS.n12650 4.608
R24758 VSS.n13081 VSS.n12650 4.608
R24759 VSS.n13082 VSS.n13081 4.608
R24760 VSS.n13084 VSS.n13082 4.608
R24761 VSS.n13084 VSS.n13083 4.608
R24762 VSS.n13083 VSS.n12646 4.608
R24763 VSS.n13091 VSS.n12646 4.608
R24764 VSS.n8853 VSS.n8852 4.608
R24765 VSS.n8852 VSS.n8851 4.608
R24766 VSS.n8851 VSS.n6969 4.608
R24767 VSS.n8845 VSS.n6969 4.608
R24768 VSS.n8845 VSS.n8844 4.608
R24769 VSS.n8844 VSS.n8843 4.608
R24770 VSS.n8843 VSS.n6973 4.608
R24771 VSS.n8837 VSS.n6973 4.608
R24772 VSS.n8837 VSS.n8836 4.608
R24773 VSS.n8836 VSS.n8835 4.608
R24774 VSS.n8835 VSS.n6977 4.608
R24775 VSS.n8829 VSS.n6977 4.608
R24776 VSS.n8776 VSS.n7254 4.608
R24777 VSS.n8777 VSS.n8776 4.608
R24778 VSS.n8778 VSS.n8777 4.608
R24779 VSS.n8778 VSS.n7250 4.608
R24780 VSS.n8784 VSS.n7250 4.608
R24781 VSS.n8785 VSS.n8784 4.608
R24782 VSS.n8786 VSS.n8785 4.608
R24783 VSS.n8786 VSS.n7246 4.608
R24784 VSS.n8793 VSS.n7246 4.608
R24785 VSS.n8794 VSS.n8793 4.608
R24786 VSS.n8795 VSS.n8794 4.608
R24787 VSS.n8795 VSS.n7239 4.608
R24788 VSS.n8631 VSS.n8630 4.608
R24789 VSS.n8630 VSS.n8629 4.608
R24790 VSS.n8629 VSS.n7325 4.608
R24791 VSS.n8623 VSS.n7325 4.608
R24792 VSS.n8623 VSS.n8622 4.608
R24793 VSS.n8622 VSS.n8621 4.608
R24794 VSS.n8621 VSS.n7329 4.608
R24795 VSS.n8615 VSS.n7329 4.608
R24796 VSS.n8615 VSS.n8614 4.608
R24797 VSS.n8614 VSS.n8613 4.608
R24798 VSS.n8613 VSS.n7333 4.608
R24799 VSS.n8607 VSS.n7333 4.608
R24800 VSS.n8554 VSS.n7394 4.608
R24801 VSS.n8555 VSS.n8554 4.608
R24802 VSS.n8556 VSS.n8555 4.608
R24803 VSS.n8556 VSS.n7390 4.608
R24804 VSS.n8562 VSS.n7390 4.608
R24805 VSS.n8563 VSS.n8562 4.608
R24806 VSS.n8564 VSS.n8563 4.608
R24807 VSS.n8564 VSS.n7386 4.608
R24808 VSS.n8571 VSS.n7386 4.608
R24809 VSS.n8572 VSS.n8571 4.608
R24810 VSS.n8573 VSS.n8572 4.608
R24811 VSS.n8573 VSS.n7379 4.608
R24812 VSS.n8273 VSS.n8272 4.608
R24813 VSS.n8272 VSS.n8271 4.608
R24814 VSS.n8271 VSS.n7465 4.608
R24815 VSS.n8265 VSS.n7465 4.608
R24816 VSS.n8265 VSS.n8264 4.608
R24817 VSS.n8264 VSS.n8263 4.608
R24818 VSS.n8263 VSS.n7469 4.608
R24819 VSS.n8257 VSS.n7469 4.608
R24820 VSS.n8257 VSS.n8256 4.608
R24821 VSS.n8256 VSS.n8255 4.608
R24822 VSS.n8255 VSS.n7473 4.608
R24823 VSS.n8249 VSS.n7473 4.608
R24824 VSS.n8196 VSS.n7534 4.608
R24825 VSS.n8197 VSS.n8196 4.608
R24826 VSS.n8198 VSS.n8197 4.608
R24827 VSS.n8198 VSS.n7530 4.608
R24828 VSS.n8204 VSS.n7530 4.608
R24829 VSS.n8205 VSS.n8204 4.608
R24830 VSS.n8206 VSS.n8205 4.608
R24831 VSS.n8206 VSS.n7526 4.608
R24832 VSS.n8213 VSS.n7526 4.608
R24833 VSS.n8214 VSS.n8213 4.608
R24834 VSS.n8215 VSS.n8214 4.608
R24835 VSS.n8215 VSS.n7519 4.608
R24836 VSS.n7915 VSS.n7914 4.608
R24837 VSS.n7914 VSS.n7913 4.608
R24838 VSS.n7913 VSS.n7605 4.608
R24839 VSS.n7907 VSS.n7605 4.608
R24840 VSS.n7907 VSS.n7906 4.608
R24841 VSS.n7906 VSS.n7905 4.608
R24842 VSS.n7905 VSS.n7609 4.608
R24843 VSS.n7899 VSS.n7609 4.608
R24844 VSS.n7899 VSS.n7898 4.608
R24845 VSS.n7898 VSS.n7897 4.608
R24846 VSS.n7897 VSS.n7613 4.608
R24847 VSS.n7891 VSS.n7613 4.608
R24848 VSS.n5580 VSS.n5579 4.608
R24849 VSS.n5580 VSS.n3684 4.608
R24850 VSS.n5586 VSS.n3684 4.608
R24851 VSS.n5587 VSS.n5586 4.608
R24852 VSS.n5588 VSS.n5587 4.608
R24853 VSS.n5588 VSS.n3680 4.608
R24854 VSS.n5594 VSS.n3680 4.608
R24855 VSS.n5595 VSS.n5594 4.608
R24856 VSS.n5597 VSS.n5595 4.608
R24857 VSS.n5597 VSS.n5596 4.608
R24858 VSS.n5596 VSS.n3676 4.608
R24859 VSS.n5604 VSS.n3676 4.608
R24860 VSS.n5315 VSS.n3756 4.608
R24861 VSS.n5309 VSS.n3756 4.608
R24862 VSS.n5309 VSS.n5308 4.608
R24863 VSS.n5308 VSS.n5307 4.608
R24864 VSS.n5307 VSS.n3760 4.608
R24865 VSS.n5301 VSS.n3760 4.608
R24866 VSS.n5301 VSS.n5300 4.608
R24867 VSS.n5300 VSS.n5299 4.608
R24868 VSS.n5299 VSS.n3764 4.608
R24869 VSS.n5293 VSS.n3764 4.608
R24870 VSS.n5293 VSS.n5292 4.608
R24871 VSS.n5292 VSS.n5291 4.608
R24872 VSS.n5234 VSS.n5233 4.608
R24873 VSS.n5234 VSS.n3825 4.608
R24874 VSS.n5240 VSS.n3825 4.608
R24875 VSS.n5241 VSS.n5240 4.608
R24876 VSS.n5242 VSS.n5241 4.608
R24877 VSS.n5242 VSS.n3821 4.608
R24878 VSS.n5248 VSS.n3821 4.608
R24879 VSS.n5249 VSS.n5248 4.608
R24880 VSS.n5251 VSS.n5249 4.608
R24881 VSS.n5251 VSS.n5250 4.608
R24882 VSS.n5250 VSS.n3817 4.608
R24883 VSS.n5258 VSS.n3817 4.608
R24884 VSS.n4958 VSS.n3897 4.608
R24885 VSS.n4952 VSS.n3897 4.608
R24886 VSS.n4952 VSS.n4951 4.608
R24887 VSS.n4951 VSS.n4950 4.608
R24888 VSS.n4950 VSS.n3901 4.608
R24889 VSS.n4944 VSS.n3901 4.608
R24890 VSS.n4944 VSS.n4943 4.608
R24891 VSS.n4943 VSS.n4942 4.608
R24892 VSS.n4942 VSS.n3905 4.608
R24893 VSS.n4936 VSS.n3905 4.608
R24894 VSS.n4936 VSS.n4935 4.608
R24895 VSS.n4935 VSS.n4934 4.608
R24896 VSS.n4877 VSS.n4876 4.608
R24897 VSS.n4877 VSS.n3966 4.608
R24898 VSS.n4883 VSS.n3966 4.608
R24899 VSS.n4884 VSS.n4883 4.608
R24900 VSS.n4885 VSS.n4884 4.608
R24901 VSS.n4885 VSS.n3962 4.608
R24902 VSS.n4891 VSS.n3962 4.608
R24903 VSS.n4892 VSS.n4891 4.608
R24904 VSS.n4894 VSS.n4892 4.608
R24905 VSS.n4894 VSS.n4893 4.608
R24906 VSS.n4893 VSS.n3958 4.608
R24907 VSS.n4901 VSS.n3958 4.608
R24908 VSS.n4601 VSS.n4038 4.608
R24909 VSS.n4595 VSS.n4038 4.608
R24910 VSS.n4595 VSS.n4594 4.608
R24911 VSS.n4594 VSS.n4593 4.608
R24912 VSS.n4593 VSS.n4042 4.608
R24913 VSS.n4587 VSS.n4042 4.608
R24914 VSS.n4587 VSS.n4586 4.608
R24915 VSS.n4586 VSS.n4585 4.608
R24916 VSS.n4585 VSS.n4046 4.608
R24917 VSS.n4579 VSS.n4046 4.608
R24918 VSS.n4579 VSS.n4578 4.608
R24919 VSS.n4578 VSS.n4577 4.608
R24920 VSS.n4520 VSS.n4519 4.608
R24921 VSS.n4520 VSS.n4107 4.608
R24922 VSS.n4526 VSS.n4107 4.608
R24923 VSS.n4527 VSS.n4526 4.608
R24924 VSS.n4528 VSS.n4527 4.608
R24925 VSS.n4528 VSS.n4103 4.608
R24926 VSS.n4534 VSS.n4103 4.608
R24927 VSS.n4535 VSS.n4534 4.608
R24928 VSS.n4537 VSS.n4535 4.608
R24929 VSS.n4537 VSS.n4536 4.608
R24930 VSS.n4536 VSS.n4099 4.608
R24931 VSS.n4544 VSS.n4099 4.608
R24932 VSS.n2966 VSS.n1308 4.608
R24933 VSS.n2972 VSS.n1308 4.608
R24934 VSS.n2973 VSS.n2972 4.608
R24935 VSS.n2974 VSS.n2973 4.608
R24936 VSS.n2974 VSS.n1304 4.608
R24937 VSS.n2980 VSS.n1304 4.608
R24938 VSS.n2981 VSS.n2980 4.608
R24939 VSS.n2982 VSS.n2981 4.608
R24940 VSS.n2982 VSS.n1300 4.608
R24941 VSS.n2988 VSS.n1300 4.608
R24942 VSS.n2989 VSS.n2988 4.608
R24943 VSS.n2990 VSS.n2989 4.608
R24944 VSS.n1389 VSS.n1377 4.608
R24945 VSS.n2676 VSS.n1389 4.608
R24946 VSS.n2676 VSS.n2675 4.608
R24947 VSS.n2675 VSS.n2674 4.608
R24948 VSS.n2674 VSS.n1390 4.608
R24949 VSS.n2668 VSS.n1390 4.608
R24950 VSS.n2668 VSS.n2667 4.608
R24951 VSS.n2667 VSS.n2666 4.608
R24952 VSS.n2666 VSS.n1394 4.608
R24953 VSS.n2660 VSS.n1394 4.608
R24954 VSS.n2660 VSS.n2659 4.608
R24955 VSS.n2659 VSS.n2658 4.608
R24956 VSS.n2323 VSS.n2291 4.608
R24957 VSS.n2317 VSS.n2291 4.608
R24958 VSS.n2317 VSS.n2316 4.608
R24959 VSS.n2316 VSS.n2315 4.608
R24960 VSS.n2315 VSS.n2295 4.608
R24961 VSS.n2309 VSS.n2295 4.608
R24962 VSS.n2309 VSS.n2308 4.608
R24963 VSS.n2308 VSS.n2307 4.608
R24964 VSS.n2307 VSS.n2299 4.608
R24965 VSS.n2301 VSS.n2299 4.608
R24966 VSS.n2301 VSS.n1451 4.608
R24967 VSS.n2627 VSS.n1451 4.608
R24968 VSS.n2576 VSS.n2575 4.608
R24969 VSS.n2577 VSS.n2576 4.608
R24970 VSS.n2577 VSS.n1473 4.608
R24971 VSS.n2583 VSS.n1473 4.608
R24972 VSS.n2584 VSS.n2583 4.608
R24973 VSS.n2585 VSS.n2584 4.608
R24974 VSS.n2585 VSS.n1469 4.608
R24975 VSS.n2591 VSS.n1469 4.608
R24976 VSS.n2592 VSS.n2591 4.608
R24977 VSS.n2593 VSS.n2592 4.608
R24978 VSS.n2593 VSS.n1465 4.608
R24979 VSS.n2599 VSS.n1465 4.608
R24980 VSS.n2105 VSS.n1549 4.608
R24981 VSS.n1553 VSS.n1549 4.608
R24982 VSS.n2098 VSS.n1553 4.608
R24983 VSS.n2098 VSS.n2097 4.608
R24984 VSS.n2097 VSS.n2096 4.608
R24985 VSS.n2096 VSS.n1554 4.608
R24986 VSS.n2090 VSS.n1554 4.608
R24987 VSS.n2090 VSS.n2089 4.608
R24988 VSS.n2089 VSS.n2088 4.608
R24989 VSS.n2088 VSS.n1558 4.608
R24990 VSS.n2082 VSS.n1558 4.608
R24991 VSS.n2082 VSS.n2081 4.608
R24992 VSS.n1714 VSS.n1682 4.608
R24993 VSS.n1708 VSS.n1682 4.608
R24994 VSS.n1708 VSS.n1707 4.608
R24995 VSS.n1707 VSS.n1706 4.608
R24996 VSS.n1706 VSS.n1686 4.608
R24997 VSS.n1700 VSS.n1686 4.608
R24998 VSS.n1700 VSS.n1699 4.608
R24999 VSS.n1699 VSS.n1698 4.608
R25000 VSS.n1698 VSS.n1690 4.608
R25001 VSS.n1692 VSS.n1690 4.608
R25002 VSS.n1692 VSS.n1577 4.608
R25003 VSS.n2019 VSS.n1577 4.608
R25004 sky130_asc_pnp_05v5_W3p40L3p40_8_0/VGND sky130_asc_pfet_01v8_lvt_6_0/VGND 4.583
R25005 VSS.n17717 sky130_asc_res_xhigh_po_2p85_1_7/VGND 4.535
R25006 VSS.n17465 VSS.n16025 4.5
R25007 VSS.n17465 VSS.n17464 4.5
R25008 VSS.n17483 VSS.n17482 4.5
R25009 VSS.n13960 VSS.n13959 4.5
R25010 VSS.n6897 VSS.n6896 4.5
R25011 VSS.n6898 VSS.n6897 4.5
R25012 VSS.n1264 VSS.n1 4.5
R25013 VSS.n3049 VSS.n1 4.5
R25014 VSS.n17715 sky130_asc_cap_mim_m3_1_2/VGND 4.414
R25015 VSS.n10462 VSS.t12 4.35
R25016 VSS.n10462 VSS.t2 4.35
R25017 VSS.n10435 VSS.t3 4.35
R25018 VSS.n10435 VSS.t8 4.35
R25019 VSS.n10434 VSS.t5 4.35
R25020 VSS.n10434 VSS.t6 4.35
R25021 VSS.n10432 VSS.t11 4.35
R25022 VSS.n10432 VSS.t9 4.35
R25023 VSS.n17642 VSS.t1 4.35
R25024 VSS.n15949 VSS.n15948 4.3
R25025 VSS.n15916 VSS.n14054 4.3
R25026 VSS.n15417 VSS.n14157 4.3
R25027 VSS.n15386 VSS.n15385 4.3
R25028 VSS.n15359 VSS.n15358 4.3
R25029 VSS.n14840 VSS.n14839 4.3
R25030 VSS.n14779 VSS.n14778 4.3
R25031 VSS.n12164 VSS.n12163 4.3
R25032 VSS.n12434 VSS.n12433 4.3
R25033 VSS.n12460 VSS.n12459 4.3
R25034 VSS.n13373 VSS.n11496 4.3
R25035 VSS.n13341 VSS.n13340 4.3
R25036 VSS.n13124 VSS.n12597 4.3
R25037 VSS.n13092 VSS.n13091 4.3
R25038 VSS.n8829 VSS.n8828 4.3
R25039 VSS.n8803 VSS.n7239 4.3
R25040 VSS.n8607 VSS.n8606 4.3
R25041 VSS.n8581 VSS.n7379 4.3
R25042 VSS.n8249 VSS.n8248 4.3
R25043 VSS.n8223 VSS.n7519 4.3
R25044 VSS.n7891 VSS.n7890 4.3
R25045 VSS.n5605 VSS.n5604 4.3
R25046 VSS.n5291 VSS.n3768 4.3
R25047 VSS.n5259 VSS.n5258 4.3
R25048 VSS.n4934 VSS.n3909 4.3
R25049 VSS.n4902 VSS.n4901 4.3
R25050 VSS.n4577 VSS.n4050 4.3
R25051 VSS.n4545 VSS.n4544 4.3
R25052 VSS.n2990 VSS.n1295 4.3
R25053 VSS.n2658 VSS.n1398 4.3
R25054 VSS.n2627 VSS.n2626 4.3
R25055 VSS.n2600 VSS.n2599 4.3
R25056 VSS.n2081 VSS.n2080 4.3
R25057 VSS.n2020 VSS.n2019 4.3
R25058 VSS.n10454 VSS.n10453 4.141
R25059 VSS.n10479 VSS.n10478 4.141
R25060 VSS.n17666 VSS.n17665 4.141
R25061 VSS.n17696 VSS.n17694 4.141
R25062 VSS.n17335 VSS.n17334 4.088
R25063 VSS.n17309 VSS.n17308 4.088
R25064 VSS.n17219 VSS.n17218 4.088
R25065 VSS.n17129 VSS.n17128 4.088
R25066 VSS.n17039 VSS.n17038 4.088
R25067 VSS.n16949 VSS.n16948 4.088
R25068 VSS.n16859 VSS.n16858 4.088
R25069 VSS.n16769 VSS.n16768 4.088
R25070 VSS.n11236 VSS.n11235 4.088
R25071 VSS.n11326 VSS.n11325 4.088
R25072 VSS.n11416 VSS.n11415 4.088
R25073 VSS.n13536 VSS.n13535 4.088
R25074 VSS.n13626 VSS.n13625 4.088
R25075 VSS.n13716 VSS.n13715 4.088
R25076 VSS.n13806 VSS.n13805 4.088
R25077 VSS.n13835 VSS.n13834 4.088
R25078 VSS.n9148 VSS.n9147 4.088
R25079 VSS.n10264 VSS.n10263 4.088
R25080 VSS.n10174 VSS.n10173 4.088
R25081 VSS.n10084 VSS.n10083 4.088
R25082 VSS.n9994 VSS.n9993 4.088
R25083 VSS.n9904 VSS.n9903 4.088
R25084 VSS.n9814 VSS.n9813 4.088
R25085 VSS.n9163 VSS.n9162 4.088
R25086 VSS.n5667 VSS.n5666 4.088
R25087 VSS.n5789 VSS.n5788 4.088
R25088 VSS.n5911 VSS.n5910 4.088
R25089 VSS.n6033 VSS.n6032 4.088
R25090 VSS.n6155 VSS.n6154 4.088
R25091 VSS.n6277 VSS.n6276 4.088
R25092 VSS.n6399 VSS.n6398 4.088
R25093 VSS.n6590 VSS.n6589 4.088
R25094 VSS.n1172 VSS.n1171 4.088
R25095 VSS.n1082 VSS.n1081 4.088
R25096 VSS.n992 VSS.n991 4.088
R25097 VSS.n902 VSS.n901 4.088
R25098 VSS.n812 VSS.n811 4.088
R25099 VSS.n722 VSS.n721 4.088
R25100 VSS.n14367 VSS.n14362 4.008
R25101 VSS.n12792 VSS.n12791 4.008
R25102 VSS.n7841 VSS.n7671 4.008
R25103 VSS.n4245 VSS.n4244 4.008
R25104 VSS.n1608 VSS.n1603 4.008
R25105 sky130_asc_res_xhigh_po_2p85_1_11/VGND sky130_asc_res_xhigh_po_2p85_1_13/VGND 3.953
R25106 VSS.n17719 sky130_asc_nfet_01v8_lvt_9_0/VGND 3.8
R25107 VSS.n17713 sky130_asc_nfet_01v8_lvt_1_0/VGND 3.76
R25108 VSS.n1263 VSS.n3 3.733
R25109 VSS.n9156 VSS.n8985 3.732
R25110 VSS.n17714 sky130_asc_cap_mim_m3_1_1/VGND 3.7
R25111 VSS.n17716 sky130_asc_pfet_01v8_lvt_60_2/VGND 3.698
R25112 sky130_asc_res_xhigh_po_2p85_1_20/VGND sky130_asc_pfet_01v8_lvt_6_1/VGND 3.584
R25113 VSS.n16626 VSS.n16620 3.582
R25114 VSS.n16725 VSS.n16627 3.582
R25115 VSS.n16731 VSS.n16625 3.582
R25116 VSS.n16737 VSS.n16628 3.582
R25117 VSS.n16743 VSS.n16624 3.582
R25118 VSS.n16749 VSS.n16629 3.582
R25119 VSS.n16758 VSS.n16623 3.582
R25120 VSS.n16763 VSS.n16630 3.582
R25121 VSS.n16536 VSS.n16530 3.582
R25122 VSS.n16815 VSS.n16537 3.582
R25123 VSS.n16821 VSS.n16535 3.582
R25124 VSS.n16827 VSS.n16538 3.582
R25125 VSS.n16833 VSS.n16534 3.582
R25126 VSS.n16839 VSS.n16539 3.582
R25127 VSS.n16848 VSS.n16533 3.582
R25128 VSS.n16853 VSS.n16540 3.582
R25129 VSS.n16446 VSS.n16440 3.582
R25130 VSS.n16905 VSS.n16447 3.582
R25131 VSS.n16911 VSS.n16445 3.582
R25132 VSS.n16917 VSS.n16448 3.582
R25133 VSS.n16923 VSS.n16444 3.582
R25134 VSS.n16929 VSS.n16449 3.582
R25135 VSS.n16938 VSS.n16443 3.582
R25136 VSS.n16943 VSS.n16450 3.582
R25137 VSS.n16356 VSS.n16350 3.582
R25138 VSS.n16995 VSS.n16357 3.582
R25139 VSS.n17001 VSS.n16355 3.582
R25140 VSS.n17007 VSS.n16358 3.582
R25141 VSS.n17013 VSS.n16354 3.582
R25142 VSS.n17019 VSS.n16359 3.582
R25143 VSS.n17028 VSS.n16353 3.582
R25144 VSS.n17033 VSS.n16360 3.582
R25145 VSS.n16266 VSS.n16260 3.582
R25146 VSS.n17085 VSS.n16267 3.582
R25147 VSS.n17091 VSS.n16265 3.582
R25148 VSS.n17097 VSS.n16268 3.582
R25149 VSS.n17103 VSS.n16264 3.582
R25150 VSS.n17109 VSS.n16269 3.582
R25151 VSS.n17118 VSS.n16263 3.582
R25152 VSS.n17123 VSS.n16270 3.582
R25153 VSS.n16176 VSS.n16170 3.582
R25154 VSS.n17175 VSS.n16177 3.582
R25155 VSS.n17181 VSS.n16175 3.582
R25156 VSS.n17187 VSS.n16178 3.582
R25157 VSS.n17193 VSS.n16174 3.582
R25158 VSS.n17199 VSS.n16179 3.582
R25159 VSS.n17208 VSS.n16173 3.582
R25160 VSS.n17213 VSS.n16180 3.582
R25161 VSS.n16086 VSS.n16080 3.582
R25162 VSS.n17265 VSS.n16087 3.582
R25163 VSS.n17271 VSS.n16085 3.582
R25164 VSS.n17277 VSS.n16088 3.582
R25165 VSS.n17283 VSS.n16084 3.582
R25166 VSS.n17289 VSS.n16089 3.582
R25167 VSS.n17298 VSS.n16083 3.582
R25168 VSS.n17303 VSS.n16090 3.582
R25169 VSS.n17427 VSS.n16044 3.582
R25170 VSS.n17433 VSS.n16045 3.582
R25171 VSS.n17439 VSS.n16043 3.582
R25172 VSS.n17445 VSS.n16046 3.582
R25173 VSS.n17454 VSS.n16042 3.582
R25174 VSS.n17459 VSS.n16047 3.582
R25175 VSS.n17386 VSS.n16041 3.582
R25176 VSS.n17421 VSS.n16040 3.582
R25177 VSS.n13919 VSS.n10511 3.582
R25178 VSS.n13925 VSS.n10512 3.582
R25179 VSS.n13931 VSS.n10510 3.582
R25180 VSS.n13937 VSS.n10513 3.582
R25181 VSS.n13946 VSS.n10509 3.582
R25182 VSS.n13951 VSS.n10514 3.582
R25183 VSS.n13886 VSS.n10508 3.582
R25184 VSS.n10553 VSS.n10547 3.582
R25185 VSS.n13769 VSS.n10554 3.582
R25186 VSS.n13775 VSS.n10555 3.582
R25187 VSS.n13781 VSS.n10551 3.582
R25188 VSS.n13787 VSS.n10556 3.582
R25189 VSS.n13796 VSS.n10550 3.582
R25190 VSS.n13801 VSS.n10557 3.582
R25191 VSS.n10643 VSS.n10637 3.582
R25192 VSS.n13679 VSS.n10644 3.582
R25193 VSS.n13685 VSS.n10645 3.582
R25194 VSS.n13691 VSS.n10641 3.582
R25195 VSS.n13697 VSS.n10646 3.582
R25196 VSS.n13706 VSS.n10640 3.582
R25197 VSS.n13711 VSS.n10647 3.582
R25198 VSS.n10733 VSS.n10727 3.582
R25199 VSS.n13589 VSS.n10734 3.582
R25200 VSS.n13595 VSS.n10735 3.582
R25201 VSS.n13601 VSS.n10731 3.582
R25202 VSS.n13607 VSS.n10736 3.582
R25203 VSS.n13616 VSS.n10730 3.582
R25204 VSS.n13621 VSS.n10737 3.582
R25205 VSS.n10823 VSS.n10817 3.582
R25206 VSS.n13498 VSS.n10824 3.582
R25207 VSS.n13504 VSS.n10825 3.582
R25208 VSS.n13510 VSS.n10821 3.582
R25209 VSS.n13517 VSS.n10826 3.582
R25210 VSS.n13526 VSS.n10820 3.582
R25211 VSS.n13531 VSS.n10827 3.582
R25212 VSS.n10913 VSS.n10907 3.582
R25213 VSS.n11379 VSS.n10914 3.582
R25214 VSS.n11385 VSS.n10915 3.582
R25215 VSS.n11391 VSS.n10911 3.582
R25216 VSS.n11397 VSS.n10916 3.582
R25217 VSS.n11406 VSS.n10910 3.582
R25218 VSS.n11411 VSS.n10917 3.582
R25219 VSS.n11003 VSS.n10997 3.582
R25220 VSS.n11289 VSS.n11004 3.582
R25221 VSS.n11295 VSS.n11005 3.582
R25222 VSS.n11301 VSS.n11001 3.582
R25223 VSS.n11307 VSS.n11006 3.582
R25224 VSS.n11316 VSS.n11000 3.582
R25225 VSS.n11321 VSS.n11007 3.582
R25226 VSS.n11093 VSS.n11087 3.582
R25227 VSS.n11199 VSS.n11094 3.582
R25228 VSS.n11205 VSS.n11095 3.582
R25229 VSS.n11211 VSS.n11091 3.582
R25230 VSS.n11217 VSS.n11096 3.582
R25231 VSS.n11226 VSS.n11090 3.582
R25232 VSS.n11231 VSS.n11097 3.582
R25233 VSS.n11188 VSS.n11092 3.582
R25234 VSS.n11278 VSS.n11002 3.582
R25235 VSS.n11368 VSS.n10912 3.582
R25236 VSS.n13487 VSS.n10822 3.582
R25237 VSS.n13578 VSS.n10732 3.582
R25238 VSS.n13668 VSS.n10642 3.582
R25239 VSS.n13758 VSS.n10552 3.582
R25240 VSS.n10499 VSS.n10495 3.582
R25241 VSS.n9671 VSS.n9665 3.582
R25242 VSS.n9770 VSS.n9672 3.582
R25243 VSS.n9776 VSS.n9670 3.582
R25244 VSS.n9782 VSS.n9673 3.582
R25245 VSS.n9788 VSS.n9669 3.582
R25246 VSS.n9794 VSS.n9674 3.582
R25247 VSS.n9803 VSS.n9668 3.582
R25248 VSS.n9808 VSS.n9675 3.582
R25249 VSS.n9581 VSS.n9575 3.582
R25250 VSS.n9860 VSS.n9582 3.582
R25251 VSS.n9866 VSS.n9580 3.582
R25252 VSS.n9872 VSS.n9583 3.582
R25253 VSS.n9878 VSS.n9579 3.582
R25254 VSS.n9884 VSS.n9584 3.582
R25255 VSS.n9893 VSS.n9578 3.582
R25256 VSS.n9898 VSS.n9585 3.582
R25257 VSS.n9491 VSS.n9485 3.582
R25258 VSS.n9950 VSS.n9492 3.582
R25259 VSS.n9956 VSS.n9490 3.582
R25260 VSS.n9962 VSS.n9493 3.582
R25261 VSS.n9968 VSS.n9489 3.582
R25262 VSS.n9974 VSS.n9494 3.582
R25263 VSS.n9983 VSS.n9488 3.582
R25264 VSS.n9988 VSS.n9495 3.582
R25265 VSS.n9401 VSS.n9395 3.582
R25266 VSS.n10040 VSS.n9402 3.582
R25267 VSS.n10046 VSS.n9400 3.582
R25268 VSS.n10052 VSS.n9403 3.582
R25269 VSS.n10058 VSS.n9399 3.582
R25270 VSS.n10064 VSS.n9404 3.582
R25271 VSS.n10073 VSS.n9398 3.582
R25272 VSS.n10078 VSS.n9405 3.582
R25273 VSS.n9311 VSS.n9305 3.582
R25274 VSS.n10130 VSS.n9312 3.582
R25275 VSS.n10136 VSS.n9310 3.582
R25276 VSS.n10142 VSS.n9313 3.582
R25277 VSS.n10148 VSS.n9309 3.582
R25278 VSS.n10154 VSS.n9314 3.582
R25279 VSS.n10163 VSS.n9308 3.582
R25280 VSS.n10168 VSS.n9315 3.582
R25281 VSS.n9221 VSS.n9215 3.582
R25282 VSS.n10220 VSS.n9222 3.582
R25283 VSS.n10226 VSS.n9220 3.582
R25284 VSS.n10232 VSS.n9223 3.582
R25285 VSS.n10238 VSS.n9219 3.582
R25286 VSS.n10244 VSS.n9224 3.582
R25287 VSS.n10253 VSS.n9218 3.582
R25288 VSS.n10258 VSS.n9225 3.582
R25289 VSS.n9082 VSS.n9007 3.582
R25290 VSS.n9066 VSS.n9014 3.582
R25291 VSS.n9050 VSS.n9008 3.582
R25292 VSS.n9034 VSS.n9013 3.582
R25293 VSS.n9042 VSS.n9012 3.582
R25294 VSS.n9058 VSS.n9009 3.582
R25295 VSS.n9074 VSS.n9011 3.582
R25296 VSS.n9090 VSS.n9010 3.582
R25297 VSS.n10332 VSS.n10331 3.582
R25298 VSS.n10338 VSS.n10337 3.582
R25299 VSS.n10344 VSS.n10343 3.582
R25300 VSS.n10350 VSS.n10349 3.582
R25301 VSS.n10356 VSS.n10355 3.582
R25302 VSS.n10362 VSS.n10361 3.582
R25303 VSS.n10368 VSS.n10367 3.582
R25304 VSS.n9182 VSS.n9180 3.582
R25305 VSS.n3222 VSS.n3153 3.582
R25306 VSS.n3214 VSS.n3154 3.582
R25307 VSS.n3206 VSS.n3152 3.582
R25308 VSS.n3198 VSS.n3155 3.582
R25309 VSS.n3190 VSS.n3151 3.582
R25310 VSS.n3182 VSS.n3156 3.582
R25311 VSS.n3150 VSS.n3141 3.582
R25312 VSS.n6534 VSS.n3140 3.582
R25313 VSS.n6473 VSS.n6472 3.582
R25314 VSS.n6479 VSS.n6478 3.582
R25315 VSS.n6485 VSS.n6484 3.582
R25316 VSS.n6491 VSS.n6490 3.582
R25317 VSS.n6497 VSS.n6496 3.582
R25318 VSS.n6503 VSS.n6502 3.582
R25319 VSS.n6509 VSS.n6508 3.582
R25320 VSS.n6515 VSS.n6514 3.582
R25321 VSS.n6351 VSS.n6350 3.582
R25322 VSS.n6357 VSS.n6356 3.582
R25323 VSS.n6363 VSS.n6362 3.582
R25324 VSS.n6369 VSS.n6368 3.582
R25325 VSS.n6375 VSS.n6374 3.582
R25326 VSS.n6381 VSS.n6380 3.582
R25327 VSS.n6387 VSS.n6386 3.582
R25328 VSS.n6393 VSS.n6392 3.582
R25329 VSS.n6229 VSS.n6228 3.582
R25330 VSS.n6235 VSS.n6234 3.582
R25331 VSS.n6241 VSS.n6240 3.582
R25332 VSS.n6247 VSS.n6246 3.582
R25333 VSS.n6253 VSS.n6252 3.582
R25334 VSS.n6259 VSS.n6258 3.582
R25335 VSS.n6265 VSS.n6264 3.582
R25336 VSS.n6271 VSS.n6270 3.582
R25337 VSS.n6107 VSS.n6106 3.582
R25338 VSS.n6113 VSS.n6112 3.582
R25339 VSS.n6119 VSS.n6118 3.582
R25340 VSS.n6125 VSS.n6124 3.582
R25341 VSS.n6131 VSS.n6130 3.582
R25342 VSS.n6137 VSS.n6136 3.582
R25343 VSS.n6143 VSS.n6142 3.582
R25344 VSS.n6149 VSS.n6148 3.582
R25345 VSS.n5985 VSS.n5984 3.582
R25346 VSS.n5991 VSS.n5990 3.582
R25347 VSS.n5997 VSS.n5996 3.582
R25348 VSS.n6003 VSS.n6002 3.582
R25349 VSS.n6009 VSS.n6008 3.582
R25350 VSS.n6015 VSS.n6014 3.582
R25351 VSS.n6021 VSS.n6020 3.582
R25352 VSS.n6027 VSS.n6026 3.582
R25353 VSS.n5863 VSS.n5862 3.582
R25354 VSS.n5869 VSS.n5868 3.582
R25355 VSS.n5875 VSS.n5874 3.582
R25356 VSS.n5881 VSS.n5880 3.582
R25357 VSS.n5887 VSS.n5886 3.582
R25358 VSS.n5893 VSS.n5892 3.582
R25359 VSS.n5899 VSS.n5898 3.582
R25360 VSS.n5905 VSS.n5904 3.582
R25361 VSS.n5741 VSS.n5740 3.582
R25362 VSS.n5747 VSS.n5746 3.582
R25363 VSS.n5753 VSS.n5752 3.582
R25364 VSS.n5759 VSS.n5758 3.582
R25365 VSS.n5765 VSS.n5764 3.582
R25366 VSS.n5771 VSS.n5770 3.582
R25367 VSS.n5777 VSS.n5776 3.582
R25368 VSS.n5783 VSS.n5782 3.582
R25369 VSS.n579 VSS.n573 3.582
R25370 VSS.n678 VSS.n580 3.582
R25371 VSS.n684 VSS.n578 3.582
R25372 VSS.n690 VSS.n581 3.582
R25373 VSS.n696 VSS.n577 3.582
R25374 VSS.n702 VSS.n582 3.582
R25375 VSS.n711 VSS.n576 3.582
R25376 VSS.n716 VSS.n583 3.582
R25377 VSS.n489 VSS.n483 3.582
R25378 VSS.n768 VSS.n490 3.582
R25379 VSS.n774 VSS.n488 3.582
R25380 VSS.n780 VSS.n491 3.582
R25381 VSS.n786 VSS.n487 3.582
R25382 VSS.n792 VSS.n492 3.582
R25383 VSS.n801 VSS.n486 3.582
R25384 VSS.n806 VSS.n493 3.582
R25385 VSS.n399 VSS.n393 3.582
R25386 VSS.n858 VSS.n400 3.582
R25387 VSS.n864 VSS.n398 3.582
R25388 VSS.n870 VSS.n401 3.582
R25389 VSS.n876 VSS.n397 3.582
R25390 VSS.n882 VSS.n402 3.582
R25391 VSS.n891 VSS.n396 3.582
R25392 VSS.n896 VSS.n403 3.582
R25393 VSS.n309 VSS.n303 3.582
R25394 VSS.n948 VSS.n310 3.582
R25395 VSS.n954 VSS.n308 3.582
R25396 VSS.n960 VSS.n311 3.582
R25397 VSS.n966 VSS.n307 3.582
R25398 VSS.n972 VSS.n312 3.582
R25399 VSS.n981 VSS.n306 3.582
R25400 VSS.n986 VSS.n313 3.582
R25401 VSS.n219 VSS.n213 3.582
R25402 VSS.n1038 VSS.n220 3.582
R25403 VSS.n1044 VSS.n218 3.582
R25404 VSS.n1050 VSS.n221 3.582
R25405 VSS.n1056 VSS.n217 3.582
R25406 VSS.n1062 VSS.n222 3.582
R25407 VSS.n1071 VSS.n216 3.582
R25408 VSS.n1076 VSS.n223 3.582
R25409 VSS.n129 VSS.n123 3.582
R25410 VSS.n1128 VSS.n130 3.582
R25411 VSS.n1134 VSS.n128 3.582
R25412 VSS.n1140 VSS.n131 3.582
R25413 VSS.n1146 VSS.n127 3.582
R25414 VSS.n1152 VSS.n132 3.582
R25415 VSS.n1161 VSS.n126 3.582
R25416 VSS.n1166 VSS.n133 3.582
R25417 VSS.n38 VSS.n32 3.582
R25418 VSS.n1213 VSS.n39 3.582
R25419 VSS.n1219 VSS.n37 3.582
R25420 VSS.n1225 VSS.n40 3.582
R25421 VSS.n1231 VSS.n36 3.582
R25422 VSS.n1237 VSS.n41 3.582
R25423 VSS.n1246 VSS.n35 3.582
R25424 VSS.n1251 VSS.n42 3.582
R25425 VSS.n3134 VSS.n3112 3.455
R25426 VSS.n10415 VSS.n10401 3.425
R25427 VSS.n3113 VSS.n3112 3.412
R25428 VSS.n3128 VSS.n3114 3.41
R25429 VSS.n3127 VSS.n3126 3.41
R25430 VSS.n10460 VSS.n10439 3.388
R25431 VSS.n10484 VSS.n10483 3.388
R25432 VSS.n17661 VSS.n17660 3.388
R25433 VSS.n17701 VSS.n17700 3.388
R25434 sky130_asc_res_xhigh_po_2p85_1_27/VGND VSS.n17550 3.376
R25435 VSS.n13994 VSS.n13993 3.033
R25436 sky130_asc_pnp_05v5_W3p40L3p40_1_0/xm1/Base VSS.n6703 3.022
R25437 sky130_asc_res_xhigh_po_2p85_1_29/VGND VSS.n17525 3.012
R25438 VSS.n10456 VSS.n10439 3.011
R25439 VSS.n10483 VSS.n10482 3.011
R25440 VSS.n17662 VSS.n17661 3.011
R25441 VSS.n17700 VSS.n17643 3.011
R25442 VSS.n10461 VSS.n10438 2.942
R25443 VSS.n17658 VSS.n17657 2.942
R25444 VSS.n15798 VSS.n15670 2.917
R25445 VSS.n15891 VSS.n15890 2.917
R25446 VSS.n15455 VSS.n15454 2.917
R25447 VSS.n15231 VSS.n15083 2.917
R25448 VSS.n15323 VSS.n14236 2.917
R25449 VSS.n14865 VSS.n14298 2.917
R25450 VSS.n14630 VSS.n14474 2.917
R25451 VSS.n12306 VSS.n11984 2.917
R25452 VSS.n12398 VSS.n11541 2.917
R25453 VSS.n11775 VSS.n11603 2.917
R25454 VSS.n13398 VSS.n11480 2.917
R25455 VSS.n13314 VSS.n12518 2.917
R25456 VSS.n13149 VSS.n12584 2.917
R25457 VSS.n13065 VSS.n12659 2.917
R25458 VSS.n7071 VSS.n6968 2.917
R25459 VSS.n8764 VSS.n8734 2.917
R25460 VSS.n7324 VSS.n7317 2.917
R25461 VSS.n8542 VSS.n8376 2.917
R25462 VSS.n7464 VSS.n7457 2.917
R25463 VSS.n8184 VSS.n8018 2.917
R25464 VSS.n7604 VSS.n7597 2.917
R25465 VSS.n5578 VSS.n3689 2.917
R25466 VSS.n5316 VSS.n3755 2.917
R25467 VSS.n5232 VSS.n3830 2.917
R25468 VSS.n4959 VSS.n3896 2.917
R25469 VSS.n4875 VSS.n3971 2.917
R25470 VSS.n4602 VSS.n4037 2.917
R25471 VSS.n4518 VSS.n4112 2.917
R25472 VSS.n2965 VSS.n2964 2.917
R25473 VSS.n2696 VSS.n2695 2.917
R25474 VSS.n2472 VSS.n2324 2.917
R25475 VSS.n2564 VSS.n1477 2.917
R25476 VSS.n2106 VSS.n1539 2.917
R25477 VSS.n1871 VSS.n1715 2.917
R25478 VSS.n17704 VSS.n17703 2.901
R25479 sky130_asc_res_xhigh_po_2p85_1_12/VGND sky130_asc_res_xhigh_po_2p85_1_14/VGND 2.83
R25480 sky130_asc_res_xhigh_po_2p85_1_14/VGND sky130_asc_res_xhigh_po_2p85_1_10/VGND 2.83
R25481 sky130_asc_res_xhigh_po_2p85_1_10/VGND sky130_asc_res_xhigh_po_2p85_1_30/VGND 2.83
R25482 sky130_asc_res_xhigh_po_2p85_1_30/VGND sky130_asc_res_xhigh_po_2p85_1_29/VGND 2.83
R25483 sky130_asc_res_xhigh_po_2p85_1_21/VGND sky130_asc_res_xhigh_po_2p85_1_24/VGND 2.83
R25484 sky130_asc_res_xhigh_po_2p85_1_24/VGND sky130_asc_res_xhigh_po_2p85_1_3/VGND 2.83
R25485 sky130_asc_res_xhigh_po_2p85_1_18/VGND sky130_asc_res_xhigh_po_2p85_1_20/VGND 2.83
R25486 sky130_asc_res_xhigh_po_2p85_1_15/VGND sky130_asc_res_xhigh_po_2p85_1_11/VGND 2.83
R25487 sky130_asc_res_xhigh_po_2p85_1_13/VGND sky130_asc_res_xhigh_po_2p85_1_28/VGND 2.83
R25488 sky130_asc_res_xhigh_po_2p85_1_28/VGND sky130_asc_res_xhigh_po_2p85_1_26/VGND 2.83
R25489 sky130_asc_res_xhigh_po_2p85_1_26/VGND sky130_asc_res_xhigh_po_2p85_1_23/VGND 2.83
R25490 sky130_asc_res_xhigh_po_2p85_1_23/VGND sky130_asc_res_xhigh_po_2p85_1_25/VGND 2.83
R25491 sky130_asc_res_xhigh_po_2p85_1_25/VGND sky130_asc_res_xhigh_po_2p85_1_27/VGND 2.83
R25492 sky130_asc_res_xhigh_po_2p85_1_9/VGND sky130_asc_res_xhigh_po_2p85_1_2/VGND 2.825
R25493 sky130_asc_res_xhigh_po_2p85_1_2/VGND sky130_asc_res_xhigh_po_2p85_1_4/VGND 2.825
R25494 sky130_asc_res_xhigh_po_2p85_1_6/VGND sky130_asc_res_xhigh_po_2p85_1_5/VGND 2.825
R25495 sky130_asc_cap_mim_m3_1_8/VGND sky130_asc_res_xhigh_po_2p85_1_21/VGND 2.811
R25496 sky130_asc_cap_mim_m3_1_6/VGND sky130_asc_res_xhigh_po_2p85_1_9/VGND 2.806
R25497 sky130_asc_cap_mim_m3_1_7/VGND sky130_asc_res_xhigh_po_2p85_1_6/VGND 2.806
R25498 sky130_asc_pfet_01v8_lvt_12_1/VGND sky130_asc_res_xhigh_po_2p85_1_7/VGND 2.804
R25499 VSS.n15670 VSS.n15636 2.715
R25500 VSS.n15891 VSS.n14072 2.715
R25501 VSS.n15454 VSS.n15453 2.715
R25502 VSS.n15083 VSS.n15049 2.715
R25503 VSS.n15324 VSS.n14236 2.715
R25504 VSS.n14866 VSS.n14865 2.715
R25505 VSS.n14474 VSS.n14440 2.715
R25506 VSS.n11984 VSS.n11983 2.715
R25507 VSS.n12399 VSS.n11541 2.715
R25508 VSS.n11775 VSS.n11774 2.715
R25509 VSS.n13399 VSS.n13398 2.715
R25510 VSS.n13314 VSS.n13313 2.715
R25511 VSS.n13149 VSS.n12583 2.715
R25512 VSS.n13065 VSS.n13064 2.715
R25513 VSS.n7069 VSS.n6968 2.715
R25514 VSS.n8765 VSS.n8764 2.715
R25515 VSS.n8453 VSS.n7324 2.715
R25516 VSS.n8543 VSS.n8542 2.715
R25517 VSS.n8095 VSS.n7464 2.715
R25518 VSS.n8185 VSS.n8184 2.715
R25519 VSS.n7744 VSS.n7604 2.715
R25520 VSS.n5578 VSS.n5577 2.715
R25521 VSS.n5316 VSS.n3754 2.715
R25522 VSS.n5232 VSS.n5231 2.715
R25523 VSS.n4959 VSS.n3895 2.715
R25524 VSS.n4875 VSS.n4874 2.715
R25525 VSS.n4602 VSS.n4036 2.715
R25526 VSS.n4518 VSS.n4517 2.715
R25527 VSS.n2965 VSS.n1313 2.715
R25528 VSS.n2695 VSS.n2694 2.715
R25529 VSS.n2324 VSS.n2290 2.715
R25530 VSS.n2565 VSS.n1477 2.715
R25531 VSS.n2107 VSS.n2106 2.715
R25532 VSS.n1715 VSS.n1681 2.715
R25533 VSS.n6895 VSS.n6894 2.563
R25534 VSS.n10487 VSS.n10486 2.529
R25535 VSS.n10372 sky130_asc_pnp_05v5_W3p40L3p40_8_1/VGND 2.423
R25536 sky130_asc_res_xhigh_po_2p85_1_5/VGND VSS.n10487 2.404
R25537 VSS.n10487 sky130_asc_nfet_01v8_lvt_9_0/VGND 2.398
R25538 sky130_asc_pnp_05v5_W3p40L3p40_1_0/Base VSS.n6699 2.311
R25539 VSS.n17420 VSS.n16025 2.287
R25540 VSS.n13959 VSS.n13958 2.287
R25541 VSS.n13964 VSS.n13963 2.287
R25542 VSS.n13961 VSS.n10400 2.258
R25543 VSS.n10453 VSS.n10452 2.258
R25544 VSS.n10478 VSS.n10477 2.258
R25545 VSS.n17667 VSS.n17666 2.258
R25546 VSS.n17694 VSS.n17693 2.258
R25547 VSS.n17466 VSS.n16024 2.248
R25548 VSS.n17484 VSS.n17483 2.246
R25549 VSS.n6895 VSS.n6883 2.245
R25550 VSS.n3051 VSS.n3050 2.243
R25551 VSS.n10459 VSS.n10438 2.228
R25552 VSS.n17659 VSS.n17658 2.228
R25553 VSS.n14364 VSS.n14363 1.95
R25554 VSS.n12790 VSS.n12723 1.95
R25555 VSS.n7840 VSS.n7672 1.95
R25556 VSS.n6758 VSS.n6757 1.95
R25557 VSS.n4243 VSS.n4176 1.95
R25558 VSS.n1605 VSS.n1604 1.95
R25559 sky130_asc_nfet_01v8_lvt_9_2/VGND VSS.n6900 1.929
R25560 VSS.n17387 VSS.n17312 1.777
R25561 VSS.n17387 VSS.n16051 1.777
R25562 VSS.n17395 VSS.n17394 1.777
R25563 VSS.n17396 VSS.n17395 1.777
R25564 VSS.n17456 VSS.n17455 1.777
R25565 VSS.n17455 VSS.n16049 1.777
R25566 VSS.n17447 VSS.n17446 1.777
R25567 VSS.n17446 VSS.n17444 1.777
R25568 VSS.n17440 VSS.n17404 1.777
R25569 VSS.n17440 VSS.n17438 1.777
R25570 VSS.n17434 VSS.n17408 1.777
R25571 VSS.n17428 VSS.n17412 1.777
R25572 VSS.n17428 VSS.n17426 1.777
R25573 VSS.n17422 VSS.n17415 1.777
R25574 VSS.n17422 VSS.n17420 1.777
R25575 VSS.n17462 VSS.n16027 1.777
R25576 VSS.n17462 VSS.n16028 1.777
R25577 VSS.n17226 VSS.n17225 1.777
R25578 VSS.n17227 VSS.n17226 1.777
R25579 VSS.n17300 VSS.n17299 1.777
R25580 VSS.n17299 VSS.n16092 1.777
R25581 VSS.n17291 VSS.n17290 1.777
R25582 VSS.n17290 VSS.n17288 1.777
R25583 VSS.n17284 VSS.n17235 1.777
R25584 VSS.n17284 VSS.n17282 1.777
R25585 VSS.n17278 VSS.n17239 1.777
R25586 VSS.n17278 VSS.n17276 1.777
R25587 VSS.n17272 VSS.n17243 1.777
R25588 VSS.n17266 VSS.n17247 1.777
R25589 VSS.n17266 VSS.n17264 1.777
R25590 VSS.n17260 VSS.n16081 1.777
R25591 VSS.n17260 VSS.n17259 1.777
R25592 VSS.n17255 VSS.n17253 1.777
R25593 VSS.n17255 VSS.n17254 1.777
R25594 VSS.n17136 VSS.n17135 1.777
R25595 VSS.n17137 VSS.n17136 1.777
R25596 VSS.n17210 VSS.n17209 1.777
R25597 VSS.n17209 VSS.n16182 1.777
R25598 VSS.n17201 VSS.n17200 1.777
R25599 VSS.n17200 VSS.n17198 1.777
R25600 VSS.n17194 VSS.n17145 1.777
R25601 VSS.n17194 VSS.n17192 1.777
R25602 VSS.n17188 VSS.n17149 1.777
R25603 VSS.n17188 VSS.n17186 1.777
R25604 VSS.n17182 VSS.n17153 1.777
R25605 VSS.n17176 VSS.n17157 1.777
R25606 VSS.n17176 VSS.n17174 1.777
R25607 VSS.n17170 VSS.n16171 1.777
R25608 VSS.n17170 VSS.n17169 1.777
R25609 VSS.n17165 VSS.n17163 1.777
R25610 VSS.n17165 VSS.n17164 1.777
R25611 VSS.n17046 VSS.n17045 1.777
R25612 VSS.n17047 VSS.n17046 1.777
R25613 VSS.n17120 VSS.n17119 1.777
R25614 VSS.n17119 VSS.n16272 1.777
R25615 VSS.n17111 VSS.n17110 1.777
R25616 VSS.n17110 VSS.n17108 1.777
R25617 VSS.n17104 VSS.n17055 1.777
R25618 VSS.n17104 VSS.n17102 1.777
R25619 VSS.n17098 VSS.n17059 1.777
R25620 VSS.n17098 VSS.n17096 1.777
R25621 VSS.n17092 VSS.n17063 1.777
R25622 VSS.n17086 VSS.n17067 1.777
R25623 VSS.n17086 VSS.n17084 1.777
R25624 VSS.n17080 VSS.n16261 1.777
R25625 VSS.n17080 VSS.n17079 1.777
R25626 VSS.n17075 VSS.n17073 1.777
R25627 VSS.n17075 VSS.n17074 1.777
R25628 VSS.n16956 VSS.n16955 1.777
R25629 VSS.n16957 VSS.n16956 1.777
R25630 VSS.n17030 VSS.n17029 1.777
R25631 VSS.n17029 VSS.n16362 1.777
R25632 VSS.n17021 VSS.n17020 1.777
R25633 VSS.n17020 VSS.n17018 1.777
R25634 VSS.n17014 VSS.n16965 1.777
R25635 VSS.n17014 VSS.n17012 1.777
R25636 VSS.n17008 VSS.n16969 1.777
R25637 VSS.n17008 VSS.n17006 1.777
R25638 VSS.n17002 VSS.n16973 1.777
R25639 VSS.n16996 VSS.n16977 1.777
R25640 VSS.n16996 VSS.n16994 1.777
R25641 VSS.n16990 VSS.n16351 1.777
R25642 VSS.n16990 VSS.n16989 1.777
R25643 VSS.n16985 VSS.n16983 1.777
R25644 VSS.n16985 VSS.n16984 1.777
R25645 VSS.n16866 VSS.n16865 1.777
R25646 VSS.n16867 VSS.n16866 1.777
R25647 VSS.n16940 VSS.n16939 1.777
R25648 VSS.n16939 VSS.n16452 1.777
R25649 VSS.n16931 VSS.n16930 1.777
R25650 VSS.n16930 VSS.n16928 1.777
R25651 VSS.n16924 VSS.n16875 1.777
R25652 VSS.n16924 VSS.n16922 1.777
R25653 VSS.n16918 VSS.n16879 1.777
R25654 VSS.n16918 VSS.n16916 1.777
R25655 VSS.n16912 VSS.n16883 1.777
R25656 VSS.n16906 VSS.n16887 1.777
R25657 VSS.n16906 VSS.n16904 1.777
R25658 VSS.n16900 VSS.n16441 1.777
R25659 VSS.n16900 VSS.n16899 1.777
R25660 VSS.n16895 VSS.n16893 1.777
R25661 VSS.n16895 VSS.n16894 1.777
R25662 VSS.n16776 VSS.n16775 1.777
R25663 VSS.n16777 VSS.n16776 1.777
R25664 VSS.n16850 VSS.n16849 1.777
R25665 VSS.n16849 VSS.n16542 1.777
R25666 VSS.n16841 VSS.n16840 1.777
R25667 VSS.n16840 VSS.n16838 1.777
R25668 VSS.n16834 VSS.n16785 1.777
R25669 VSS.n16834 VSS.n16832 1.777
R25670 VSS.n16828 VSS.n16789 1.777
R25671 VSS.n16828 VSS.n16826 1.777
R25672 VSS.n16822 VSS.n16793 1.777
R25673 VSS.n16816 VSS.n16797 1.777
R25674 VSS.n16816 VSS.n16814 1.777
R25675 VSS.n16810 VSS.n16531 1.777
R25676 VSS.n16810 VSS.n16809 1.777
R25677 VSS.n16805 VSS.n16803 1.777
R25678 VSS.n16805 VSS.n16804 1.777
R25679 VSS.n16686 VSS.n16685 1.777
R25680 VSS.n16687 VSS.n16686 1.777
R25681 VSS.n16760 VSS.n16759 1.777
R25682 VSS.n16759 VSS.n16632 1.777
R25683 VSS.n16751 VSS.n16750 1.777
R25684 VSS.n16750 VSS.n16748 1.777
R25685 VSS.n16744 VSS.n16695 1.777
R25686 VSS.n16744 VSS.n16742 1.777
R25687 VSS.n16738 VSS.n16699 1.777
R25688 VSS.n16738 VSS.n16736 1.777
R25689 VSS.n16732 VSS.n16703 1.777
R25690 VSS.n16726 VSS.n16707 1.777
R25691 VSS.n16726 VSS.n16724 1.777
R25692 VSS.n16720 VSS.n16621 1.777
R25693 VSS.n16720 VSS.n16719 1.777
R25694 VSS.n16715 VSS.n16713 1.777
R25695 VSS.n16715 VSS.n16714 1.777
R25696 VSS.n11153 VSS.n11152 1.777
R25697 VSS.n11154 VSS.n11153 1.777
R25698 VSS.n11228 VSS.n11227 1.777
R25699 VSS.n11227 VSS.n11099 1.777
R25700 VSS.n11219 VSS.n11218 1.777
R25701 VSS.n11218 VSS.n11216 1.777
R25702 VSS.n11212 VSS.n11162 1.777
R25703 VSS.n11212 VSS.n11210 1.777
R25704 VSS.n11206 VSS.n11166 1.777
R25705 VSS.n11206 VSS.n11204 1.777
R25706 VSS.n11200 VSS.n11170 1.777
R25707 VSS.n11194 VSS.n11088 1.777
R25708 VSS.n11194 VSS.n11193 1.777
R25709 VSS.n11189 VSS.n11176 1.777
R25710 VSS.n11189 VSS.n11187 1.777
R25711 VSS.n11183 VSS.n11181 1.777
R25712 VSS.n11183 VSS.n11182 1.777
R25713 VSS.n11243 VSS.n11242 1.777
R25714 VSS.n11244 VSS.n11243 1.777
R25715 VSS.n11318 VSS.n11317 1.777
R25716 VSS.n11317 VSS.n11009 1.777
R25717 VSS.n11309 VSS.n11308 1.777
R25718 VSS.n11308 VSS.n11306 1.777
R25719 VSS.n11302 VSS.n11252 1.777
R25720 VSS.n11302 VSS.n11300 1.777
R25721 VSS.n11296 VSS.n11256 1.777
R25722 VSS.n11296 VSS.n11294 1.777
R25723 VSS.n11290 VSS.n11260 1.777
R25724 VSS.n11284 VSS.n10998 1.777
R25725 VSS.n11284 VSS.n11283 1.777
R25726 VSS.n11279 VSS.n11266 1.777
R25727 VSS.n11279 VSS.n11277 1.777
R25728 VSS.n11273 VSS.n11271 1.777
R25729 VSS.n11273 VSS.n11272 1.777
R25730 VSS.n11333 VSS.n11332 1.777
R25731 VSS.n11334 VSS.n11333 1.777
R25732 VSS.n11408 VSS.n11407 1.777
R25733 VSS.n11407 VSS.n10919 1.777
R25734 VSS.n11399 VSS.n11398 1.777
R25735 VSS.n11398 VSS.n11396 1.777
R25736 VSS.n11392 VSS.n11342 1.777
R25737 VSS.n11392 VSS.n11390 1.777
R25738 VSS.n11386 VSS.n11346 1.777
R25739 VSS.n11386 VSS.n11384 1.777
R25740 VSS.n11380 VSS.n11350 1.777
R25741 VSS.n11374 VSS.n10908 1.777
R25742 VSS.n11374 VSS.n11373 1.777
R25743 VSS.n11369 VSS.n11356 1.777
R25744 VSS.n11369 VSS.n11367 1.777
R25745 VSS.n11363 VSS.n11361 1.777
R25746 VSS.n11363 VSS.n11362 1.777
R25747 VSS.n11423 VSS.n11422 1.777
R25748 VSS.n11424 VSS.n11423 1.777
R25749 VSS.n13528 VSS.n13527 1.777
R25750 VSS.n13527 VSS.n10829 1.777
R25751 VSS.n13519 VSS.n13518 1.777
R25752 VSS.n13518 VSS.n13516 1.777
R25753 VSS.n13511 VSS.n13461 1.777
R25754 VSS.n13511 VSS.n13509 1.777
R25755 VSS.n13505 VSS.n13465 1.777
R25756 VSS.n13505 VSS.n13503 1.777
R25757 VSS.n13499 VSS.n13469 1.777
R25758 VSS.n13493 VSS.n10818 1.777
R25759 VSS.n13493 VSS.n13492 1.777
R25760 VSS.n13488 VSS.n13475 1.777
R25761 VSS.n13488 VSS.n13486 1.777
R25762 VSS.n13482 VSS.n13480 1.777
R25763 VSS.n13482 VSS.n13481 1.777
R25764 VSS.n13543 VSS.n13542 1.777
R25765 VSS.n13544 VSS.n13543 1.777
R25766 VSS.n13618 VSS.n13617 1.777
R25767 VSS.n13617 VSS.n10739 1.777
R25768 VSS.n13609 VSS.n13608 1.777
R25769 VSS.n13608 VSS.n13606 1.777
R25770 VSS.n13602 VSS.n13552 1.777
R25771 VSS.n13602 VSS.n13600 1.777
R25772 VSS.n13596 VSS.n13556 1.777
R25773 VSS.n13596 VSS.n13594 1.777
R25774 VSS.n13590 VSS.n13560 1.777
R25775 VSS.n13584 VSS.n10728 1.777
R25776 VSS.n13584 VSS.n13583 1.777
R25777 VSS.n13579 VSS.n13566 1.777
R25778 VSS.n13579 VSS.n13577 1.777
R25779 VSS.n13573 VSS.n13571 1.777
R25780 VSS.n13573 VSS.n13572 1.777
R25781 VSS.n13633 VSS.n13632 1.777
R25782 VSS.n13634 VSS.n13633 1.777
R25783 VSS.n13708 VSS.n13707 1.777
R25784 VSS.n13707 VSS.n10649 1.777
R25785 VSS.n13699 VSS.n13698 1.777
R25786 VSS.n13698 VSS.n13696 1.777
R25787 VSS.n13692 VSS.n13642 1.777
R25788 VSS.n13692 VSS.n13690 1.777
R25789 VSS.n13686 VSS.n13646 1.777
R25790 VSS.n13686 VSS.n13684 1.777
R25791 VSS.n13680 VSS.n13650 1.777
R25792 VSS.n13674 VSS.n10638 1.777
R25793 VSS.n13674 VSS.n13673 1.777
R25794 VSS.n13669 VSS.n13656 1.777
R25795 VSS.n13669 VSS.n13667 1.777
R25796 VSS.n13663 VSS.n13661 1.777
R25797 VSS.n13663 VSS.n13662 1.777
R25798 VSS.n13723 VSS.n13722 1.777
R25799 VSS.n13724 VSS.n13723 1.777
R25800 VSS.n13798 VSS.n13797 1.777
R25801 VSS.n13797 VSS.n10559 1.777
R25802 VSS.n13789 VSS.n13788 1.777
R25803 VSS.n13788 VSS.n13786 1.777
R25804 VSS.n13782 VSS.n13732 1.777
R25805 VSS.n13782 VSS.n13780 1.777
R25806 VSS.n13776 VSS.n13736 1.777
R25807 VSS.n13776 VSS.n13774 1.777
R25808 VSS.n13770 VSS.n13740 1.777
R25809 VSS.n13764 VSS.n10548 1.777
R25810 VSS.n13764 VSS.n13763 1.777
R25811 VSS.n13759 VSS.n13746 1.777
R25812 VSS.n13759 VSS.n13757 1.777
R25813 VSS.n13753 VSS.n13751 1.777
R25814 VSS.n13753 VSS.n13752 1.777
R25815 VSS.n13887 VSS.n13809 1.777
R25816 VSS.n13887 VSS.n10518 1.777
R25817 VSS.n13895 VSS.n13894 1.777
R25818 VSS.n13896 VSS.n13895 1.777
R25819 VSS.n13948 VSS.n13947 1.777
R25820 VSS.n13947 VSS.n10516 1.777
R25821 VSS.n13939 VSS.n13938 1.777
R25822 VSS.n13938 VSS.n13936 1.777
R25823 VSS.n13932 VSS.n13904 1.777
R25824 VSS.n13932 VSS.n13930 1.777
R25825 VSS.n13926 VSS.n13908 1.777
R25826 VSS.n13920 VSS.n13912 1.777
R25827 VSS.n13920 VSS.n13918 1.777
R25828 VSS.n13913 VSS.n10493 1.777
R25829 VSS.n13958 VSS.n10493 1.777
R25830 VSS.n10498 VSS.n10494 1.777
R25831 VSS.n13830 VSS.n10498 1.777
R25832 VSS.n9035 VSS.n8983 1.777
R25833 VSS.n9036 VSS.n9035 1.777
R25834 VSS.n9043 VSS.n9032 1.777
R25835 VSS.n9044 VSS.n9043 1.777
R25836 VSS.n9051 VSS.n9030 1.777
R25837 VSS.n9052 VSS.n9051 1.777
R25838 VSS.n9059 VSS.n9028 1.777
R25839 VSS.n9060 VSS.n9059 1.777
R25840 VSS.n9067 VSS.n9026 1.777
R25841 VSS.n9068 VSS.n9067 1.777
R25842 VSS.n9075 VSS.n9024 1.777
R25843 VSS.n9083 VSS.n9022 1.777
R25844 VSS.n9084 VSS.n9083 1.777
R25845 VSS.n9091 VSS.n9020 1.777
R25846 VSS.n9092 VSS.n9091 1.777
R25847 VSS.n9153 VSS.n9017 1.777
R25848 VSS.n9153 VSS.n9018 1.777
R25849 VSS.n10181 VSS.n10180 1.777
R25850 VSS.n10182 VSS.n10181 1.777
R25851 VSS.n10255 VSS.n10254 1.777
R25852 VSS.n10254 VSS.n9227 1.777
R25853 VSS.n10246 VSS.n10245 1.777
R25854 VSS.n10245 VSS.n10243 1.777
R25855 VSS.n10239 VSS.n10190 1.777
R25856 VSS.n10239 VSS.n10237 1.777
R25857 VSS.n10233 VSS.n10194 1.777
R25858 VSS.n10233 VSS.n10231 1.777
R25859 VSS.n10227 VSS.n10198 1.777
R25860 VSS.n10221 VSS.n10202 1.777
R25861 VSS.n10221 VSS.n10219 1.777
R25862 VSS.n10215 VSS.n9216 1.777
R25863 VSS.n10215 VSS.n10214 1.777
R25864 VSS.n10210 VSS.n10208 1.777
R25865 VSS.n10210 VSS.n10209 1.777
R25866 VSS.n10091 VSS.n10090 1.777
R25867 VSS.n10092 VSS.n10091 1.777
R25868 VSS.n10165 VSS.n10164 1.777
R25869 VSS.n10164 VSS.n9317 1.777
R25870 VSS.n10156 VSS.n10155 1.777
R25871 VSS.n10155 VSS.n10153 1.777
R25872 VSS.n10149 VSS.n10100 1.777
R25873 VSS.n10149 VSS.n10147 1.777
R25874 VSS.n10143 VSS.n10104 1.777
R25875 VSS.n10143 VSS.n10141 1.777
R25876 VSS.n10137 VSS.n10108 1.777
R25877 VSS.n10131 VSS.n10112 1.777
R25878 VSS.n10131 VSS.n10129 1.777
R25879 VSS.n10125 VSS.n9306 1.777
R25880 VSS.n10125 VSS.n10124 1.777
R25881 VSS.n10120 VSS.n10118 1.777
R25882 VSS.n10120 VSS.n10119 1.777
R25883 VSS.n10001 VSS.n10000 1.777
R25884 VSS.n10002 VSS.n10001 1.777
R25885 VSS.n10075 VSS.n10074 1.777
R25886 VSS.n10074 VSS.n9407 1.777
R25887 VSS.n10066 VSS.n10065 1.777
R25888 VSS.n10065 VSS.n10063 1.777
R25889 VSS.n10059 VSS.n10010 1.777
R25890 VSS.n10059 VSS.n10057 1.777
R25891 VSS.n10053 VSS.n10014 1.777
R25892 VSS.n10053 VSS.n10051 1.777
R25893 VSS.n10047 VSS.n10018 1.777
R25894 VSS.n10041 VSS.n10022 1.777
R25895 VSS.n10041 VSS.n10039 1.777
R25896 VSS.n10035 VSS.n9396 1.777
R25897 VSS.n10035 VSS.n10034 1.777
R25898 VSS.n10030 VSS.n10028 1.777
R25899 VSS.n10030 VSS.n10029 1.777
R25900 VSS.n9911 VSS.n9910 1.777
R25901 VSS.n9912 VSS.n9911 1.777
R25902 VSS.n9985 VSS.n9984 1.777
R25903 VSS.n9984 VSS.n9497 1.777
R25904 VSS.n9976 VSS.n9975 1.777
R25905 VSS.n9975 VSS.n9973 1.777
R25906 VSS.n9969 VSS.n9920 1.777
R25907 VSS.n9969 VSS.n9967 1.777
R25908 VSS.n9963 VSS.n9924 1.777
R25909 VSS.n9963 VSS.n9961 1.777
R25910 VSS.n9957 VSS.n9928 1.777
R25911 VSS.n9951 VSS.n9932 1.777
R25912 VSS.n9951 VSS.n9949 1.777
R25913 VSS.n9945 VSS.n9486 1.777
R25914 VSS.n9945 VSS.n9944 1.777
R25915 VSS.n9940 VSS.n9938 1.777
R25916 VSS.n9940 VSS.n9939 1.777
R25917 VSS.n9821 VSS.n9820 1.777
R25918 VSS.n9822 VSS.n9821 1.777
R25919 VSS.n9895 VSS.n9894 1.777
R25920 VSS.n9894 VSS.n9587 1.777
R25921 VSS.n9886 VSS.n9885 1.777
R25922 VSS.n9885 VSS.n9883 1.777
R25923 VSS.n9879 VSS.n9830 1.777
R25924 VSS.n9879 VSS.n9877 1.777
R25925 VSS.n9873 VSS.n9834 1.777
R25926 VSS.n9873 VSS.n9871 1.777
R25927 VSS.n9867 VSS.n9838 1.777
R25928 VSS.n9861 VSS.n9842 1.777
R25929 VSS.n9861 VSS.n9859 1.777
R25930 VSS.n9855 VSS.n9576 1.777
R25931 VSS.n9855 VSS.n9854 1.777
R25932 VSS.n9850 VSS.n9848 1.777
R25933 VSS.n9850 VSS.n9849 1.777
R25934 VSS.n9731 VSS.n9730 1.777
R25935 VSS.n9732 VSS.n9731 1.777
R25936 VSS.n9805 VSS.n9804 1.777
R25937 VSS.n9804 VSS.n9677 1.777
R25938 VSS.n9796 VSS.n9795 1.777
R25939 VSS.n9795 VSS.n9793 1.777
R25940 VSS.n9789 VSS.n9740 1.777
R25941 VSS.n9789 VSS.n9787 1.777
R25942 VSS.n9783 VSS.n9744 1.777
R25943 VSS.n9783 VSS.n9781 1.777
R25944 VSS.n9777 VSS.n9748 1.777
R25945 VSS.n9771 VSS.n9752 1.777
R25946 VSS.n9771 VSS.n9769 1.777
R25947 VSS.n9765 VSS.n9666 1.777
R25948 VSS.n9765 VSS.n9764 1.777
R25949 VSS.n9760 VSS.n9758 1.777
R25950 VSS.n9760 VSS.n9759 1.777
R25951 VSS.n10322 VSS.n10321 1.777
R25952 VSS.n10321 VSS.n9186 1.777
R25953 VSS.n10369 VSS.n8932 1.777
R25954 VSS.n10369 VSS.n8933 1.777
R25955 VSS.n10364 VSS.n10363 1.777
R25956 VSS.n10363 VSS.n8938 1.777
R25957 VSS.n10358 VSS.n10357 1.777
R25958 VSS.n10357 VSS.n8943 1.777
R25959 VSS.n10352 VSS.n10351 1.777
R25960 VSS.n10351 VSS.n8949 1.777
R25961 VSS.n10346 VSS.n10345 1.777
R25962 VSS.n10340 VSS.n10339 1.777
R25963 VSS.n10339 VSS.n8960 1.777
R25964 VSS.n10334 VSS.n10333 1.777
R25965 VSS.n10333 VSS.n8967 1.777
R25966 VSS.n10328 VSS.n10327 1.777
R25967 VSS.n10327 VSS.n8973 1.777
R25968 VSS.n5784 VSS.n3579 1.777
R25969 VSS.n5784 VSS.n3580 1.777
R25970 VSS.n5779 VSS.n5778 1.777
R25971 VSS.n5778 VSS.n3585 1.777
R25972 VSS.n5773 VSS.n5772 1.777
R25973 VSS.n5772 VSS.n3590 1.777
R25974 VSS.n5767 VSS.n5766 1.777
R25975 VSS.n5766 VSS.n3596 1.777
R25976 VSS.n5761 VSS.n5760 1.777
R25977 VSS.n5760 VSS.n3602 1.777
R25978 VSS.n5755 VSS.n5754 1.777
R25979 VSS.n5749 VSS.n5748 1.777
R25980 VSS.n5748 VSS.n3613 1.777
R25981 VSS.n5743 VSS.n5742 1.777
R25982 VSS.n5742 VSS.n3620 1.777
R25983 VSS.n5737 VSS.n5736 1.777
R25984 VSS.n5736 VSS.n3626 1.777
R25985 VSS.n5906 VSS.n3521 1.777
R25986 VSS.n5906 VSS.n3522 1.777
R25987 VSS.n5901 VSS.n5900 1.777
R25988 VSS.n5900 VSS.n3527 1.777
R25989 VSS.n5895 VSS.n5894 1.777
R25990 VSS.n5894 VSS.n3532 1.777
R25991 VSS.n5889 VSS.n5888 1.777
R25992 VSS.n5888 VSS.n3538 1.777
R25993 VSS.n5883 VSS.n5882 1.777
R25994 VSS.n5882 VSS.n3544 1.777
R25995 VSS.n5877 VSS.n5876 1.777
R25996 VSS.n5871 VSS.n5870 1.777
R25997 VSS.n5870 VSS.n3555 1.777
R25998 VSS.n5865 VSS.n5864 1.777
R25999 VSS.n5864 VSS.n3562 1.777
R26000 VSS.n5859 VSS.n5858 1.777
R26001 VSS.n5858 VSS.n3568 1.777
R26002 VSS.n6028 VSS.n3463 1.777
R26003 VSS.n6028 VSS.n3464 1.777
R26004 VSS.n6023 VSS.n6022 1.777
R26005 VSS.n6022 VSS.n3469 1.777
R26006 VSS.n6017 VSS.n6016 1.777
R26007 VSS.n6016 VSS.n3474 1.777
R26008 VSS.n6011 VSS.n6010 1.777
R26009 VSS.n6010 VSS.n3480 1.777
R26010 VSS.n6005 VSS.n6004 1.777
R26011 VSS.n6004 VSS.n3486 1.777
R26012 VSS.n5999 VSS.n5998 1.777
R26013 VSS.n5993 VSS.n5992 1.777
R26014 VSS.n5992 VSS.n3497 1.777
R26015 VSS.n5987 VSS.n5986 1.777
R26016 VSS.n5986 VSS.n3504 1.777
R26017 VSS.n5981 VSS.n5980 1.777
R26018 VSS.n5980 VSS.n3510 1.777
R26019 VSS.n6150 VSS.n3405 1.777
R26020 VSS.n6150 VSS.n3406 1.777
R26021 VSS.n6145 VSS.n6144 1.777
R26022 VSS.n6144 VSS.n3411 1.777
R26023 VSS.n6139 VSS.n6138 1.777
R26024 VSS.n6138 VSS.n3416 1.777
R26025 VSS.n6133 VSS.n6132 1.777
R26026 VSS.n6132 VSS.n3422 1.777
R26027 VSS.n6127 VSS.n6126 1.777
R26028 VSS.n6126 VSS.n3428 1.777
R26029 VSS.n6121 VSS.n6120 1.777
R26030 VSS.n6115 VSS.n6114 1.777
R26031 VSS.n6114 VSS.n3439 1.777
R26032 VSS.n6109 VSS.n6108 1.777
R26033 VSS.n6108 VSS.n3446 1.777
R26034 VSS.n6103 VSS.n6102 1.777
R26035 VSS.n6102 VSS.n3452 1.777
R26036 VSS.n6272 VSS.n3347 1.777
R26037 VSS.n6272 VSS.n3348 1.777
R26038 VSS.n6267 VSS.n6266 1.777
R26039 VSS.n6266 VSS.n3353 1.777
R26040 VSS.n6261 VSS.n6260 1.777
R26041 VSS.n6260 VSS.n3358 1.777
R26042 VSS.n6255 VSS.n6254 1.777
R26043 VSS.n6254 VSS.n3364 1.777
R26044 VSS.n6249 VSS.n6248 1.777
R26045 VSS.n6248 VSS.n3370 1.777
R26046 VSS.n6243 VSS.n6242 1.777
R26047 VSS.n6237 VSS.n6236 1.777
R26048 VSS.n6236 VSS.n3381 1.777
R26049 VSS.n6231 VSS.n6230 1.777
R26050 VSS.n6230 VSS.n3388 1.777
R26051 VSS.n6225 VSS.n6224 1.777
R26052 VSS.n6224 VSS.n3394 1.777
R26053 VSS.n6394 VSS.n3289 1.777
R26054 VSS.n6394 VSS.n3290 1.777
R26055 VSS.n6389 VSS.n6388 1.777
R26056 VSS.n6388 VSS.n3295 1.777
R26057 VSS.n6383 VSS.n6382 1.777
R26058 VSS.n6382 VSS.n3300 1.777
R26059 VSS.n6377 VSS.n6376 1.777
R26060 VSS.n6376 VSS.n3306 1.777
R26061 VSS.n6371 VSS.n6370 1.777
R26062 VSS.n6370 VSS.n3312 1.777
R26063 VSS.n6365 VSS.n6364 1.777
R26064 VSS.n6359 VSS.n6358 1.777
R26065 VSS.n6358 VSS.n3323 1.777
R26066 VSS.n6353 VSS.n6352 1.777
R26067 VSS.n6352 VSS.n3330 1.777
R26068 VSS.n6347 VSS.n6346 1.777
R26069 VSS.n6346 VSS.n3336 1.777
R26070 VSS.n6516 VSS.n3231 1.777
R26071 VSS.n6516 VSS.n3232 1.777
R26072 VSS.n6511 VSS.n6510 1.777
R26073 VSS.n6510 VSS.n3237 1.777
R26074 VSS.n6505 VSS.n6504 1.777
R26075 VSS.n6504 VSS.n3242 1.777
R26076 VSS.n6499 VSS.n6498 1.777
R26077 VSS.n6498 VSS.n3248 1.777
R26078 VSS.n6493 VSS.n6492 1.777
R26079 VSS.n6492 VSS.n3254 1.777
R26080 VSS.n6487 VSS.n6486 1.777
R26081 VSS.n6481 VSS.n6480 1.777
R26082 VSS.n6480 VSS.n3265 1.777
R26083 VSS.n6475 VSS.n6474 1.777
R26084 VSS.n6474 VSS.n3272 1.777
R26085 VSS.n6469 VSS.n6468 1.777
R26086 VSS.n6468 VSS.n3278 1.777
R26087 VSS.n6536 VSS.n3138 1.777
R26088 VSS.n6603 VSS.n3138 1.777
R26089 VSS.n3175 VSS.n3139 1.777
R26090 VSS.n3176 VSS.n3175 1.777
R26091 VSS.n3183 VSS.n3172 1.777
R26092 VSS.n3184 VSS.n3183 1.777
R26093 VSS.n3191 VSS.n3170 1.777
R26094 VSS.n3192 VSS.n3191 1.777
R26095 VSS.n3199 VSS.n3168 1.777
R26096 VSS.n3200 VSS.n3199 1.777
R26097 VSS.n3207 VSS.n3166 1.777
R26098 VSS.n3215 VSS.n3164 1.777
R26099 VSS.n3216 VSS.n3215 1.777
R26100 VSS.n3223 VSS.n3162 1.777
R26101 VSS.n3224 VSS.n3223 1.777
R26102 VSS.n6595 VSS.n3159 1.777
R26103 VSS.n6595 VSS.n3160 1.777
R26104 VSS.n1179 VSS.n1178 1.777
R26105 VSS.n1180 VSS.n1179 1.777
R26106 VSS.n1248 VSS.n1247 1.777
R26107 VSS.n1247 VSS.n44 1.777
R26108 VSS.n1239 VSS.n1238 1.777
R26109 VSS.n1238 VSS.n1236 1.777
R26110 VSS.n1232 VSS.n1188 1.777
R26111 VSS.n1232 VSS.n1230 1.777
R26112 VSS.n1226 VSS.n1192 1.777
R26113 VSS.n1226 VSS.n1224 1.777
R26114 VSS.n1220 VSS.n1196 1.777
R26115 VSS.n1214 VSS.n1200 1.777
R26116 VSS.n1214 VSS.n1212 1.777
R26117 VSS.n1208 VSS.n33 1.777
R26118 VSS.n1208 VSS.n1207 1.777
R26119 VSS.n1256 VSS.n6 1.777
R26120 VSS.n1257 VSS.n1256 1.777
R26121 VSS.n1089 VSS.n1088 1.777
R26122 VSS.n1090 VSS.n1089 1.777
R26123 VSS.n1163 VSS.n1162 1.777
R26124 VSS.n1162 VSS.n135 1.777
R26125 VSS.n1154 VSS.n1153 1.777
R26126 VSS.n1153 VSS.n1151 1.777
R26127 VSS.n1147 VSS.n1098 1.777
R26128 VSS.n1147 VSS.n1145 1.777
R26129 VSS.n1141 VSS.n1102 1.777
R26130 VSS.n1141 VSS.n1139 1.777
R26131 VSS.n1135 VSS.n1106 1.777
R26132 VSS.n1129 VSS.n1110 1.777
R26133 VSS.n1129 VSS.n1127 1.777
R26134 VSS.n1123 VSS.n124 1.777
R26135 VSS.n1123 VSS.n1122 1.777
R26136 VSS.n1118 VSS.n1116 1.777
R26137 VSS.n1118 VSS.n1117 1.777
R26138 VSS.n999 VSS.n998 1.777
R26139 VSS.n1000 VSS.n999 1.777
R26140 VSS.n1073 VSS.n1072 1.777
R26141 VSS.n1072 VSS.n225 1.777
R26142 VSS.n1064 VSS.n1063 1.777
R26143 VSS.n1063 VSS.n1061 1.777
R26144 VSS.n1057 VSS.n1008 1.777
R26145 VSS.n1057 VSS.n1055 1.777
R26146 VSS.n1051 VSS.n1012 1.777
R26147 VSS.n1051 VSS.n1049 1.777
R26148 VSS.n1045 VSS.n1016 1.777
R26149 VSS.n1039 VSS.n1020 1.777
R26150 VSS.n1039 VSS.n1037 1.777
R26151 VSS.n1033 VSS.n214 1.777
R26152 VSS.n1033 VSS.n1032 1.777
R26153 VSS.n1028 VSS.n1026 1.777
R26154 VSS.n1028 VSS.n1027 1.777
R26155 VSS.n909 VSS.n908 1.777
R26156 VSS.n910 VSS.n909 1.777
R26157 VSS.n983 VSS.n982 1.777
R26158 VSS.n982 VSS.n315 1.777
R26159 VSS.n974 VSS.n973 1.777
R26160 VSS.n973 VSS.n971 1.777
R26161 VSS.n967 VSS.n918 1.777
R26162 VSS.n967 VSS.n965 1.777
R26163 VSS.n961 VSS.n922 1.777
R26164 VSS.n961 VSS.n959 1.777
R26165 VSS.n955 VSS.n926 1.777
R26166 VSS.n949 VSS.n930 1.777
R26167 VSS.n949 VSS.n947 1.777
R26168 VSS.n943 VSS.n304 1.777
R26169 VSS.n943 VSS.n942 1.777
R26170 VSS.n938 VSS.n936 1.777
R26171 VSS.n938 VSS.n937 1.777
R26172 VSS.n819 VSS.n818 1.777
R26173 VSS.n820 VSS.n819 1.777
R26174 VSS.n893 VSS.n892 1.777
R26175 VSS.n892 VSS.n405 1.777
R26176 VSS.n884 VSS.n883 1.777
R26177 VSS.n883 VSS.n881 1.777
R26178 VSS.n877 VSS.n828 1.777
R26179 VSS.n877 VSS.n875 1.777
R26180 VSS.n871 VSS.n832 1.777
R26181 VSS.n871 VSS.n869 1.777
R26182 VSS.n865 VSS.n836 1.777
R26183 VSS.n859 VSS.n840 1.777
R26184 VSS.n859 VSS.n857 1.777
R26185 VSS.n853 VSS.n394 1.777
R26186 VSS.n853 VSS.n852 1.777
R26187 VSS.n848 VSS.n846 1.777
R26188 VSS.n848 VSS.n847 1.777
R26189 VSS.n729 VSS.n728 1.777
R26190 VSS.n730 VSS.n729 1.777
R26191 VSS.n803 VSS.n802 1.777
R26192 VSS.n802 VSS.n495 1.777
R26193 VSS.n794 VSS.n793 1.777
R26194 VSS.n793 VSS.n791 1.777
R26195 VSS.n787 VSS.n738 1.777
R26196 VSS.n787 VSS.n785 1.777
R26197 VSS.n781 VSS.n742 1.777
R26198 VSS.n781 VSS.n779 1.777
R26199 VSS.n775 VSS.n746 1.777
R26200 VSS.n769 VSS.n750 1.777
R26201 VSS.n769 VSS.n767 1.777
R26202 VSS.n763 VSS.n484 1.777
R26203 VSS.n763 VSS.n762 1.777
R26204 VSS.n758 VSS.n756 1.777
R26205 VSS.n758 VSS.n757 1.777
R26206 VSS.n639 VSS.n638 1.777
R26207 VSS.n640 VSS.n639 1.777
R26208 VSS.n713 VSS.n712 1.777
R26209 VSS.n712 VSS.n585 1.777
R26210 VSS.n704 VSS.n703 1.777
R26211 VSS.n703 VSS.n701 1.777
R26212 VSS.n697 VSS.n648 1.777
R26213 VSS.n697 VSS.n695 1.777
R26214 VSS.n691 VSS.n652 1.777
R26215 VSS.n691 VSS.n689 1.777
R26216 VSS.n685 VSS.n656 1.777
R26217 VSS.n679 VSS.n660 1.777
R26218 VSS.n679 VSS.n677 1.777
R26219 VSS.n673 VSS.n574 1.777
R26220 VSS.n673 VSS.n672 1.777
R26221 VSS.n668 VSS.n666 1.777
R26222 VSS.n668 VSS.n667 1.777
R26223 sky130_asc_nfet_01v8_lvt_1_1/VGND sky130_asc_pnp_05v5_W3p40L3p40_7_0/VGND 1.766
R26224 VSS.n10417 VSS.n10416 1.707
R26225 VSS.n10414 VSS.n10402 1.7
R26226 VSS.n3132 VSS.n3131 1.7
R26227 VSS.n10462 VSS.n10426 1.686
R26228 VSS.n17679 VSS.n17642 1.686
R26229 VSS.n13960 VSS.n10490 1.51
R26230 VSS.n10448 VSS.n10447 1.505
R26231 VSS.n10473 VSS.n10472 1.505
R26232 VSS.n17673 VSS.n17671 1.505
R26233 VSS.n17687 VSS.n17646 1.505
R26234 VSS.n17468 VSS.n17467 1.502
R26235 VSS.n13962 VSS.n13961 1.5
R26236 VSS.n10488 sky130_asc_cap_mim_m3_1_7/VGND 1.374
R26237 VSS.n10488 VSS.n10417 1.363
R26238 VSS.n3135 VSS.n3134 1.356
R26239 VSS.n9155 VSS.n9154 1.309
R26240 VSS.n15796 VSS.n15672 1.292
R26241 VSS.n15796 VSS.n15673 1.292
R26242 VSS.n15790 VSS.n15789 1.292
R26243 VSS.n15789 VSS.n15683 1.292
R26244 VSS.n15778 VSS.n15687 1.292
R26245 VSS.n15778 VSS.n15777 1.292
R26246 VSS.n15773 VSS.n15694 1.292
R26247 VSS.n15773 VSS.n15695 1.292
R26248 VSS.n15767 VSS.n15766 1.292
R26249 VSS.n15766 VSS.n15702 1.292
R26250 VSS.n15755 VSS.n15706 1.292
R26251 VSS.n15755 VSS.n15754 1.292
R26252 sky130_asc_pnp_05v5_W3p40L3p40_8_3/xm1/Collector VSS.n15713 1.292
R26253 sky130_asc_pnp_05v5_W3p40L3p40_8_3/xm1/Collector VSS.n15714 1.292
R26254 VSS.n15745 VSS.n15744 1.292
R26255 VSS.n15744 VSS.n15721 1.292
R26256 VSS.n15733 VSS.n15725 1.292
R26257 VSS.n15733 VSS.n15732 1.292
R26258 VSS.n16021 VSS.n13997 1.292
R26259 VSS.n16021 VSS.n13998 1.292
R26260 VSS.n16015 VSS.n16014 1.292
R26261 VSS.n16014 VSS.n14005 1.292
R26262 VSS.n16003 VSS.n14009 1.292
R26263 VSS.n16003 VSS.n16002 1.292
R26264 VSS.n15888 VSS.n15561 1.292
R26265 VSS.n15888 VSS.n15562 1.292
R26266 VSS.n15882 VSS.n15881 1.292
R26267 VSS.n15881 VSS.n15571 1.292
R26268 VSS.n15870 VSS.n15575 1.292
R26269 VSS.n15870 VSS.n15869 1.292
R26270 VSS.n15865 VSS.n15582 1.292
R26271 VSS.n15865 VSS.n15583 1.292
R26272 VSS.n15859 VSS.n15858 1.292
R26273 VSS.n15858 VSS.n15590 1.292
R26274 VSS.n15847 VSS.n15594 1.292
R26275 VSS.n15847 VSS.n15846 1.292
R26276 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector VSS.n15601 1.292
R26277 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector VSS.n15602 1.292
R26278 VSS.n15837 VSS.n15836 1.292
R26279 VSS.n15836 VSS.n15609 1.292
R26280 VSS.n15825 VSS.n15613 1.292
R26281 VSS.n15825 VSS.n15824 1.292
R26282 VSS.n15820 VSS.n15620 1.292
R26283 VSS.n15820 VSS.n15621 1.292
R26284 VSS.n15814 VSS.n15813 1.292
R26285 VSS.n15813 VSS.n15628 1.292
R26286 VSS.n15802 VSS.n15632 1.292
R26287 VSS.n15802 VSS.n15801 1.292
R26288 VSS.n15458 VSS.n15457 1.292
R26289 VSS.n15457 VSS.n14130 1.292
R26290 VSS.n15469 VSS.n14126 1.292
R26291 VSS.n15469 VSS.n14128 1.292
R26292 VSS.n15476 VSS.n15475 1.292
R26293 VSS.n15476 VSS.n14120 1.292
R26294 VSS.n15487 VSS.n14115 1.292
R26295 VSS.n15488 VSS.n15487 1.292
R26296 VSS.n15493 VSS.n15492 1.292
R26297 VSS.n15492 VSS.n14109 1.292
R26298 VSS.n15504 VSS.n14105 1.292
R26299 VSS.n15504 VSS.n14107 1.292
R26300 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector VSS.n15510 1.292
R26301 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector VSS.n14099 1.292
R26302 VSS.n15521 VSS.n14094 1.292
R26303 VSS.n15522 VSS.n15521 1.292
R26304 VSS.n15527 VSS.n15526 1.292
R26305 VSS.n15526 VSS.n14088 1.292
R26306 VSS.n15538 VSS.n14084 1.292
R26307 VSS.n15538 VSS.n14086 1.292
R26308 VSS.n15545 VSS.n15544 1.292
R26309 VSS.n15545 VSS.n14078 1.292
R26310 VSS.n15556 VSS.n14074 1.292
R26311 VSS.n15557 VSS.n15556 1.292
R26312 VSS.n15229 VSS.n15085 1.292
R26313 VSS.n15229 VSS.n15086 1.292
R26314 VSS.n15223 VSS.n15222 1.292
R26315 VSS.n15222 VSS.n15096 1.292
R26316 VSS.n15211 VSS.n15100 1.292
R26317 VSS.n15211 VSS.n15210 1.292
R26318 VSS.n15206 VSS.n15107 1.292
R26319 VSS.n15206 VSS.n15108 1.292
R26320 VSS.n15200 VSS.n15199 1.292
R26321 VSS.n15199 VSS.n15115 1.292
R26322 VSS.n15188 VSS.n15119 1.292
R26323 VSS.n15188 VSS.n15187 1.292
R26324 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector VSS.n15126 1.292
R26325 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector VSS.n15127 1.292
R26326 VSS.n15178 VSS.n15177 1.292
R26327 VSS.n15177 VSS.n15134 1.292
R26328 VSS.n15166 VSS.n15138 1.292
R26329 VSS.n15166 VSS.n15165 1.292
R26330 VSS.n15161 VSS.n15145 1.292
R26331 VSS.n15161 VSS.n15146 1.292
R26332 VSS.n15155 VSS.n15154 1.292
R26333 VSS.n15154 VSS.n14139 1.292
R26334 VSS.n14140 VSS.n14137 1.292
R26335 VSS.n15452 VSS.n14137 1.292
R26336 VSS.n15321 VSS.n14974 1.292
R26337 VSS.n15321 VSS.n14975 1.292
R26338 VSS.n15315 VSS.n15314 1.292
R26339 VSS.n15314 VSS.n14984 1.292
R26340 VSS.n15303 VSS.n14988 1.292
R26341 VSS.n15303 VSS.n15302 1.292
R26342 VSS.n15298 VSS.n14995 1.292
R26343 VSS.n15298 VSS.n14996 1.292
R26344 VSS.n15292 VSS.n15291 1.292
R26345 VSS.n15291 VSS.n15003 1.292
R26346 VSS.n15280 VSS.n15007 1.292
R26347 VSS.n15280 VSS.n15279 1.292
R26348 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector VSS.n15014 1.292
R26349 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector VSS.n15015 1.292
R26350 VSS.n15270 VSS.n15269 1.292
R26351 VSS.n15269 VSS.n15022 1.292
R26352 VSS.n15258 VSS.n15026 1.292
R26353 VSS.n15258 VSS.n15257 1.292
R26354 VSS.n15253 VSS.n15033 1.292
R26355 VSS.n15253 VSS.n15034 1.292
R26356 VSS.n15247 VSS.n15246 1.292
R26357 VSS.n15246 VSS.n15041 1.292
R26358 VSS.n15235 VSS.n15045 1.292
R26359 VSS.n15235 VSS.n15234 1.292
R26360 VSS.n14878 VSS.n14877 1.292
R26361 VSS.n14878 VSS.n14297 1.292
R26362 VSS.n14889 VSS.n14292 1.292
R26363 VSS.n14890 VSS.n14889 1.292
R26364 VSS.n14895 VSS.n14894 1.292
R26365 VSS.n14894 VSS.n14286 1.292
R26366 VSS.n14906 VSS.n14282 1.292
R26367 VSS.n14906 VSS.n14284 1.292
R26368 VSS.n14913 VSS.n14912 1.292
R26369 VSS.n14913 VSS.n14276 1.292
R26370 VSS.n14924 VSS.n14271 1.292
R26371 VSS.n14925 VSS.n14924 1.292
R26372 VSS.n14929 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector 1.292
R26373 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector VSS.n14265 1.292
R26374 VSS.n14940 VSS.n14261 1.292
R26375 VSS.n14940 VSS.n14263 1.292
R26376 VSS.n14947 VSS.n14946 1.292
R26377 VSS.n14947 VSS.n14255 1.292
R26378 VSS.n14958 VSS.n14250 1.292
R26379 VSS.n14959 VSS.n14958 1.292
R26380 VSS.n14964 VSS.n14963 1.292
R26381 VSS.n14963 VSS.n14244 1.292
R26382 VSS.n15328 VSS.n14241 1.292
R26383 VSS.n15328 VSS.n14242 1.292
R26384 VSS.n14628 VSS.n14476 1.292
R26385 VSS.n14628 VSS.n14477 1.292
R26386 VSS.n14622 VSS.n14621 1.292
R26387 VSS.n14621 VSS.n14487 1.292
R26388 VSS.n14610 VSS.n14491 1.292
R26389 VSS.n14610 VSS.n14609 1.292
R26390 VSS.n14605 VSS.n14498 1.292
R26391 VSS.n14605 VSS.n14499 1.292
R26392 VSS.n14599 VSS.n14598 1.292
R26393 VSS.n14598 VSS.n14506 1.292
R26394 VSS.n14587 VSS.n14510 1.292
R26395 VSS.n14587 VSS.n14586 1.292
R26396 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector VSS.n14517 1.292
R26397 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector VSS.n14518 1.292
R26398 VSS.n14577 VSS.n14576 1.292
R26399 VSS.n14576 VSS.n14525 1.292
R26400 VSS.n14565 VSS.n14529 1.292
R26401 VSS.n14565 VSS.n14564 1.292
R26402 VSS.n14560 VSS.n14536 1.292
R26403 VSS.n14560 VSS.n14537 1.292
R26404 VSS.n14554 VSS.n14553 1.292
R26405 VSS.n14553 VSS.n14548 1.292
R26406 VSS.n14870 VSS.n14305 1.292
R26407 VSS.n14870 VSS.n14306 1.292
R26408 VSS.n14721 VSS.n14720 1.292
R26409 VSS.n14720 VSS.n14368 1.292
R26410 VSS.n14714 VSS.n14713 1.292
R26411 VSS.n14713 VSS.n14374 1.292
R26412 VSS.n14702 VSS.n14379 1.292
R26413 VSS.n14702 VSS.n14701 1.292
R26414 VSS.n14697 VSS.n14386 1.292
R26415 VSS.n14697 VSS.n14387 1.292
R26416 VSS.n14691 VSS.n14690 1.292
R26417 VSS.n14690 VSS.n14394 1.292
R26418 VSS.n14679 VSS.n14398 1.292
R26419 VSS.n14679 VSS.n14678 1.292
R26420 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Collector VSS.n14405 1.292
R26421 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Collector VSS.n14406 1.292
R26422 VSS.n14669 VSS.n14668 1.292
R26423 VSS.n14668 VSS.n14413 1.292
R26424 VSS.n14657 VSS.n14417 1.292
R26425 VSS.n14657 VSS.n14656 1.292
R26426 VSS.n14652 VSS.n14424 1.292
R26427 VSS.n14652 VSS.n14425 1.292
R26428 VSS.n14646 VSS.n14645 1.292
R26429 VSS.n14645 VSS.n14432 1.292
R26430 VSS.n14634 VSS.n14436 1.292
R26431 VSS.n14634 VSS.n14633 1.292
R26432 VSS.n12304 VSS.n11986 1.292
R26433 VSS.n12304 VSS.n11987 1.292
R26434 VSS.n12298 VSS.n12297 1.292
R26435 VSS.n12297 VSS.n11997 1.292
R26436 VSS.n12286 VSS.n12001 1.292
R26437 VSS.n12286 VSS.n12285 1.292
R26438 VSS.n12281 VSS.n12008 1.292
R26439 VSS.n12281 VSS.n12009 1.292
R26440 VSS.n12275 VSS.n12274 1.292
R26441 VSS.n12274 VSS.n12016 1.292
R26442 VSS.n12263 VSS.n12020 1.292
R26443 VSS.n12263 VSS.n12262 1.292
R26444 sky130_asc_pnp_05v5_W3p40L3p40_8_0/xm1/Collector VSS.n12027 1.292
R26445 sky130_asc_pnp_05v5_W3p40L3p40_8_0/xm1/Collector VSS.n12028 1.292
R26446 VSS.n12253 VSS.n12252 1.292
R26447 VSS.n12252 VSS.n12035 1.292
R26448 VSS.n12241 VSS.n12039 1.292
R26449 VSS.n12241 VSS.n12240 1.292
R26450 VSS.n12236 VSS.n12046 1.292
R26451 VSS.n12236 VSS.n12047 1.292
R26452 VSS.n12230 VSS.n12229 1.292
R26453 VSS.n12229 VSS.n12054 1.292
R26454 VSS.n12218 VSS.n12058 1.292
R26455 VSS.n12218 VSS.n12217 1.292
R26456 VSS.n12396 VSS.n11908 1.292
R26457 VSS.n12396 VSS.n11909 1.292
R26458 VSS.n12390 VSS.n12389 1.292
R26459 VSS.n12389 VSS.n11918 1.292
R26460 VSS.n12378 VSS.n11922 1.292
R26461 VSS.n12378 VSS.n12377 1.292
R26462 VSS.n12373 VSS.n11929 1.292
R26463 VSS.n12373 VSS.n11930 1.292
R26464 VSS.n12367 VSS.n12366 1.292
R26465 VSS.n12366 VSS.n11937 1.292
R26466 VSS.n12355 VSS.n11941 1.292
R26467 VSS.n12355 VSS.n12354 1.292
R26468 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector VSS.n11948 1.292
R26469 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector VSS.n11949 1.292
R26470 VSS.n12345 VSS.n12344 1.292
R26471 VSS.n12344 VSS.n11956 1.292
R26472 VSS.n12333 VSS.n11960 1.292
R26473 VSS.n12333 VSS.n12332 1.292
R26474 VSS.n12328 VSS.n11967 1.292
R26475 VSS.n12328 VSS.n11968 1.292
R26476 VSS.n12322 VSS.n12321 1.292
R26477 VSS.n12321 VSS.n11975 1.292
R26478 VSS.n12310 VSS.n11979 1.292
R26479 VSS.n12310 VSS.n12309 1.292
R26480 VSS.n11812 VSS.n11811 1.292
R26481 VSS.n11812 VSS.n11602 1.292
R26482 VSS.n11823 VSS.n11597 1.292
R26483 VSS.n11824 VSS.n11823 1.292
R26484 VSS.n11829 VSS.n11828 1.292
R26485 VSS.n11828 VSS.n11591 1.292
R26486 VSS.n11840 VSS.n11587 1.292
R26487 VSS.n11840 VSS.n11589 1.292
R26488 VSS.n11847 VSS.n11846 1.292
R26489 VSS.n11847 VSS.n11581 1.292
R26490 VSS.n11858 VSS.n11576 1.292
R26491 VSS.n11859 VSS.n11858 1.292
R26492 VSS.n11863 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector 1.292
R26493 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector VSS.n11570 1.292
R26494 VSS.n11874 VSS.n11566 1.292
R26495 VSS.n11874 VSS.n11568 1.292
R26496 VSS.n11881 VSS.n11880 1.292
R26497 VSS.n11881 VSS.n11560 1.292
R26498 VSS.n11892 VSS.n11555 1.292
R26499 VSS.n11893 VSS.n11892 1.292
R26500 VSS.n11898 VSS.n11897 1.292
R26501 VSS.n11897 VSS.n11549 1.292
R26502 VSS.n12403 VSS.n11546 1.292
R26503 VSS.n12403 VSS.n11547 1.292
R26504 VSS.n11677 VSS.n11669 1.292
R26505 VSS.n11678 VSS.n11677 1.292
R26506 VSS.n11683 VSS.n11682 1.292
R26507 VSS.n11682 VSS.n11663 1.292
R26508 VSS.n11694 VSS.n11659 1.292
R26509 VSS.n11694 VSS.n11661 1.292
R26510 VSS.n11701 VSS.n11700 1.292
R26511 VSS.n11701 VSS.n11653 1.292
R26512 VSS.n11712 VSS.n11648 1.292
R26513 VSS.n11713 VSS.n11712 1.292
R26514 VSS.n11718 VSS.n11717 1.292
R26515 VSS.n11717 VSS.n11642 1.292
R26516 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector VSS.n11638 1.292
R26517 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector VSS.n11640 1.292
R26518 VSS.n11735 VSS.n11734 1.292
R26519 VSS.n11735 VSS.n11632 1.292
R26520 VSS.n11746 VSS.n11627 1.292
R26521 VSS.n11747 VSS.n11746 1.292
R26522 VSS.n11752 VSS.n11751 1.292
R26523 VSS.n11751 VSS.n11621 1.292
R26524 VSS.n11763 VSS.n11616 1.292
R26525 VSS.n11763 VSS.n11619 1.292
R26526 VSS.n11770 VSS.n11612 1.292
R26527 VSS.n11770 VSS.n11610 1.292
R26528 VSS.n13302 VSS.n13301 1.292
R26529 VSS.n13301 VSS.n13251 1.292
R26530 VSS.n13290 VSS.n13253 1.292
R26531 VSS.n13290 VSS.n13289 1.292
R26532 VSS.n13285 VSS.n13261 1.292
R26533 VSS.n13285 VSS.n13262 1.292
R26534 VSS.n13279 VSS.n13278 1.292
R26535 VSS.n13278 VSS.n13273 1.292
R26536 VSS.n13455 VSS.n11431 1.292
R26537 VSS.n13455 VSS.n11432 1.292
R26538 VSS.n13449 VSS.n13448 1.292
R26539 VSS.n13448 VSS.n11439 1.292
R26540 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector VSS.n11443 1.292
R26541 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector VSS.n13437 1.292
R26542 VSS.n13433 VSS.n11450 1.292
R26543 VSS.n13433 VSS.n11451 1.292
R26544 VSS.n13427 VSS.n13426 1.292
R26545 VSS.n13426 VSS.n11458 1.292
R26546 VSS.n13415 VSS.n11462 1.292
R26547 VSS.n13415 VSS.n13414 1.292
R26548 VSS.n13410 VSS.n11469 1.292
R26549 VSS.n13410 VSS.n11470 1.292
R26550 VSS.n13404 VSS.n13403 1.292
R26551 VSS.n13403 VSS.n11477 1.292
R26552 VSS.n13156 VSS.n12578 1.292
R26553 VSS.n13157 VSS.n13156 1.292
R26554 VSS.n13162 VSS.n13161 1.292
R26555 VSS.n13161 VSS.n12572 1.292
R26556 VSS.n13173 VSS.n12568 1.292
R26557 VSS.n13173 VSS.n12570 1.292
R26558 VSS.n13180 VSS.n13179 1.292
R26559 VSS.n13180 VSS.n12562 1.292
R26560 VSS.n13191 VSS.n12557 1.292
R26561 VSS.n13192 VSS.n13191 1.292
R26562 VSS.n13197 VSS.n13196 1.292
R26563 VSS.n13196 VSS.n12551 1.292
R26564 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector VSS.n12547 1.292
R26565 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector VSS.n12549 1.292
R26566 VSS.n13214 VSS.n13213 1.292
R26567 VSS.n13214 VSS.n12541 1.292
R26568 VSS.n13225 VSS.n12536 1.292
R26569 VSS.n13226 VSS.n13225 1.292
R26570 VSS.n13231 VSS.n13230 1.292
R26571 VSS.n13230 VSS.n12528 1.292
R26572 VSS.n12529 VSS.n12526 1.292
R26573 VSS.n13243 VSS.n12526 1.292
R26574 VSS.n13309 VSS.n12521 1.292
R26575 VSS.n13309 VSS.n12519 1.292
R26576 VSS.n13053 VSS.n13052 1.292
R26577 VSS.n13052 VSS.n12894 1.292
R26578 VSS.n13041 VSS.n12896 1.292
R26579 VSS.n13041 VSS.n13040 1.292
R26580 VSS.n13036 VSS.n12904 1.292
R26581 VSS.n13036 VSS.n12905 1.292
R26582 VSS.n13030 VSS.n13029 1.292
R26583 VSS.n13029 VSS.n12912 1.292
R26584 VSS.n13018 VSS.n12916 1.292
R26585 VSS.n13018 VSS.n13017 1.292
R26586 VSS.n13013 VSS.n12923 1.292
R26587 VSS.n13013 VSS.n12924 1.292
R26588 VSS.n13007 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector 1.292
R26589 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector VSS.n12931 1.292
R26590 VSS.n12996 VSS.n12935 1.292
R26591 VSS.n12996 VSS.n12995 1.292
R26592 VSS.n12991 VSS.n12942 1.292
R26593 VSS.n12991 VSS.n12943 1.292
R26594 VSS.n12985 VSS.n12984 1.292
R26595 VSS.n12984 VSS.n12950 1.292
R26596 VSS.n12973 VSS.n12954 1.292
R26597 VSS.n12973 VSS.n12972 1.292
R26598 VSS.n12968 VSS.n12962 1.292
R26599 VSS.n12968 VSS.n12963 1.292
R26600 VSS.n12799 VSS.n12719 1.292
R26601 VSS.n12800 VSS.n12799 1.292
R26602 VSS.n12805 VSS.n12804 1.292
R26603 VSS.n12804 VSS.n12713 1.292
R26604 VSS.n12816 VSS.n12709 1.292
R26605 VSS.n12816 VSS.n12711 1.292
R26606 VSS.n12823 VSS.n12822 1.292
R26607 VSS.n12823 VSS.n12703 1.292
R26608 VSS.n12834 VSS.n12698 1.292
R26609 VSS.n12835 VSS.n12834 1.292
R26610 VSS.n12840 VSS.n12839 1.292
R26611 VSS.n12839 VSS.n12692 1.292
R26612 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Collector VSS.n12688 1.292
R26613 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Collector VSS.n12690 1.292
R26614 VSS.n12857 VSS.n12856 1.292
R26615 VSS.n12857 VSS.n12682 1.292
R26616 VSS.n12868 VSS.n12677 1.292
R26617 VSS.n12869 VSS.n12868 1.292
R26618 VSS.n12874 VSS.n12873 1.292
R26619 VSS.n12873 VSS.n12669 1.292
R26620 VSS.n12670 VSS.n12667 1.292
R26621 VSS.n12886 VSS.n12667 1.292
R26622 VSS.n13060 VSS.n12662 1.292
R26623 VSS.n13060 VSS.n12660 1.292
R26624 VSS.n7074 VSS.n7073 1.292
R26625 VSS.n7073 VSS.n7065 1.292
R26626 VSS.n7085 VSS.n7061 1.292
R26627 VSS.n7085 VSS.n7063 1.292
R26628 VSS.n7092 VSS.n7091 1.292
R26629 VSS.n7092 VSS.n7055 1.292
R26630 VSS.n7103 VSS.n7050 1.292
R26631 VSS.n7104 VSS.n7103 1.292
R26632 VSS.n7109 VSS.n7108 1.292
R26633 VSS.n7108 VSS.n7044 1.292
R26634 VSS.n7120 VSS.n7040 1.292
R26635 VSS.n7120 VSS.n7042 1.292
R26636 sky130_asc_pnp_05v5_W3p40L3p40_8_1/xm1/Collector VSS.n7126 1.292
R26637 sky130_asc_pnp_05v5_W3p40L3p40_8_1/xm1/Collector VSS.n7034 1.292
R26638 VSS.n7137 VSS.n7029 1.292
R26639 VSS.n7138 VSS.n7137 1.292
R26640 VSS.n7143 VSS.n7142 1.292
R26641 VSS.n7142 VSS.n7023 1.292
R26642 VSS.n7154 VSS.n7019 1.292
R26643 VSS.n7154 VSS.n7021 1.292
R26644 VSS.n7161 VSS.n7160 1.292
R26645 VSS.n7161 VSS.n7013 1.292
R26646 VSS.n7173 VSS.n7007 1.292
R26647 VSS.n7174 VSS.n7173 1.292
R26648 VSS.n8742 VSS.n8735 1.292
R26649 VSS.n8743 VSS.n8742 1.292
R26650 VSS.n8755 VSS.n8754 1.292
R26651 VSS.n8754 VSS.n8740 1.292
R26652 VSS.n8927 VSS.n6903 1.292
R26653 VSS.n8927 VSS.n6904 1.292
R26654 VSS.n8921 VSS.n8920 1.292
R26655 VSS.n8920 VSS.n6911 1.292
R26656 VSS.n8909 VSS.n6915 1.292
R26657 VSS.n8909 VSS.n8908 1.292
R26658 VSS.n8904 VSS.n6922 1.292
R26659 VSS.n8904 VSS.n6923 1.292
R26660 VSS.n8898 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector 1.292
R26661 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector VSS.n6930 1.292
R26662 VSS.n8887 VSS.n6934 1.292
R26663 VSS.n8887 VSS.n8886 1.292
R26664 VSS.n8882 VSS.n6941 1.292
R26665 VSS.n8882 VSS.n6942 1.292
R26666 VSS.n8876 VSS.n8875 1.292
R26667 VSS.n8875 VSS.n6949 1.292
R26668 VSS.n8864 VSS.n6953 1.292
R26669 VSS.n8864 VSS.n8863 1.292
R26670 VSS.n8859 VSS.n6960 1.292
R26671 VSS.n8859 VSS.n6961 1.292
R26672 VSS.n8639 VSS.n8638 1.292
R26673 VSS.n8639 VSS.n7316 1.292
R26674 VSS.n8650 VSS.n7311 1.292
R26675 VSS.n8651 VSS.n8650 1.292
R26676 VSS.n8656 VSS.n8655 1.292
R26677 VSS.n8655 VSS.n7305 1.292
R26678 VSS.n8667 VSS.n7301 1.292
R26679 VSS.n8667 VSS.n7303 1.292
R26680 VSS.n8674 VSS.n8673 1.292
R26681 VSS.n8674 VSS.n7295 1.292
R26682 VSS.n8685 VSS.n7290 1.292
R26683 VSS.n8686 VSS.n8685 1.292
R26684 VSS.n8690 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector 1.292
R26685 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector VSS.n7284 1.292
R26686 VSS.n8701 VSS.n7280 1.292
R26687 VSS.n8701 VSS.n7282 1.292
R26688 VSS.n8708 VSS.n8707 1.292
R26689 VSS.n8708 VSS.n7274 1.292
R26690 VSS.n8719 VSS.n7269 1.292
R26691 VSS.n8720 VSS.n8719 1.292
R26692 VSS.n8725 VSS.n8724 1.292
R26693 VSS.n8724 VSS.n7263 1.292
R26694 VSS.n8769 VSS.n7260 1.292
R26695 VSS.n8769 VSS.n7261 1.292
R26696 VSS.n8384 VSS.n8377 1.292
R26697 VSS.n8385 VSS.n8384 1.292
R26698 VSS.n8533 VSS.n8532 1.292
R26699 VSS.n8532 VSS.n8382 1.292
R26700 VSS.n8526 VSS.n8525 1.292
R26701 VSS.n8525 VSS.n8393 1.292
R26702 VSS.n8514 VSS.n8398 1.292
R26703 VSS.n8514 VSS.n8513 1.292
R26704 VSS.n8509 VSS.n8405 1.292
R26705 VSS.n8509 VSS.n8406 1.292
R26706 VSS.n8503 VSS.n8502 1.292
R26707 VSS.n8502 VSS.n8413 1.292
R26708 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector VSS.n8417 1.292
R26709 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector VSS.n8491 1.292
R26710 VSS.n8487 VSS.n8424 1.292
R26711 VSS.n8487 VSS.n8425 1.292
R26712 VSS.n8481 VSS.n8480 1.292
R26713 VSS.n8480 VSS.n8432 1.292
R26714 VSS.n8469 VSS.n8436 1.292
R26715 VSS.n8469 VSS.n8468 1.292
R26716 VSS.n8464 VSS.n8443 1.292
R26717 VSS.n8464 VSS.n8444 1.292
R26718 VSS.n8458 VSS.n8457 1.292
R26719 VSS.n8457 VSS.n8450 1.292
R26720 VSS.n8281 VSS.n8280 1.292
R26721 VSS.n8281 VSS.n7456 1.292
R26722 VSS.n8292 VSS.n7451 1.292
R26723 VSS.n8293 VSS.n8292 1.292
R26724 VSS.n8298 VSS.n8297 1.292
R26725 VSS.n8297 VSS.n7445 1.292
R26726 VSS.n8309 VSS.n7441 1.292
R26727 VSS.n8309 VSS.n7443 1.292
R26728 VSS.n8316 VSS.n8315 1.292
R26729 VSS.n8316 VSS.n7435 1.292
R26730 VSS.n8327 VSS.n7430 1.292
R26731 VSS.n8328 VSS.n8327 1.292
R26732 VSS.n8332 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector 1.292
R26733 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector VSS.n7424 1.292
R26734 VSS.n8343 VSS.n7420 1.292
R26735 VSS.n8343 VSS.n7422 1.292
R26736 VSS.n8350 VSS.n8349 1.292
R26737 VSS.n8350 VSS.n7414 1.292
R26738 VSS.n8361 VSS.n7409 1.292
R26739 VSS.n8362 VSS.n8361 1.292
R26740 VSS.n8367 VSS.n8366 1.292
R26741 VSS.n8366 VSS.n7403 1.292
R26742 VSS.n8547 VSS.n7400 1.292
R26743 VSS.n8547 VSS.n7401 1.292
R26744 VSS.n8026 VSS.n8019 1.292
R26745 VSS.n8027 VSS.n8026 1.292
R26746 VSS.n8175 VSS.n8174 1.292
R26747 VSS.n8174 VSS.n8024 1.292
R26748 VSS.n8168 VSS.n8167 1.292
R26749 VSS.n8167 VSS.n8035 1.292
R26750 VSS.n8156 VSS.n8040 1.292
R26751 VSS.n8156 VSS.n8155 1.292
R26752 VSS.n8151 VSS.n8047 1.292
R26753 VSS.n8151 VSS.n8048 1.292
R26754 VSS.n8145 VSS.n8144 1.292
R26755 VSS.n8144 VSS.n8055 1.292
R26756 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector VSS.n8059 1.292
R26757 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector VSS.n8133 1.292
R26758 VSS.n8129 VSS.n8066 1.292
R26759 VSS.n8129 VSS.n8067 1.292
R26760 VSS.n8123 VSS.n8122 1.292
R26761 VSS.n8122 VSS.n8074 1.292
R26762 VSS.n8111 VSS.n8078 1.292
R26763 VSS.n8111 VSS.n8110 1.292
R26764 VSS.n8106 VSS.n8085 1.292
R26765 VSS.n8106 VSS.n8086 1.292
R26766 VSS.n8100 VSS.n8099 1.292
R26767 VSS.n8099 VSS.n8092 1.292
R26768 VSS.n7923 VSS.n7922 1.292
R26769 VSS.n7923 VSS.n7596 1.292
R26770 VSS.n7934 VSS.n7591 1.292
R26771 VSS.n7935 VSS.n7934 1.292
R26772 VSS.n7940 VSS.n7939 1.292
R26773 VSS.n7939 VSS.n7585 1.292
R26774 VSS.n7951 VSS.n7581 1.292
R26775 VSS.n7951 VSS.n7583 1.292
R26776 VSS.n7958 VSS.n7957 1.292
R26777 VSS.n7958 VSS.n7575 1.292
R26778 VSS.n7969 VSS.n7570 1.292
R26779 VSS.n7970 VSS.n7969 1.292
R26780 VSS.n7974 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector 1.292
R26781 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector VSS.n7564 1.292
R26782 VSS.n7985 VSS.n7560 1.292
R26783 VSS.n7985 VSS.n7562 1.292
R26784 VSS.n7992 VSS.n7991 1.292
R26785 VSS.n7992 VSS.n7554 1.292
R26786 VSS.n8003 VSS.n7549 1.292
R26787 VSS.n8004 VSS.n8003 1.292
R26788 VSS.n8009 VSS.n8008 1.292
R26789 VSS.n8008 VSS.n7543 1.292
R26790 VSS.n8189 VSS.n7540 1.292
R26791 VSS.n8189 VSS.n7541 1.292
R26792 VSS.n7835 VSS.n7834 1.292
R26793 VSS.n7834 VSS.n7675 1.292
R26794 VSS.n7828 VSS.n7827 1.292
R26795 VSS.n7827 VSS.n7681 1.292
R26796 VSS.n7816 VSS.n7686 1.292
R26797 VSS.n7816 VSS.n7815 1.292
R26798 VSS.n7811 VSS.n7693 1.292
R26799 VSS.n7811 VSS.n7694 1.292
R26800 VSS.n7805 VSS.n7804 1.292
R26801 VSS.n7804 VSS.n7701 1.292
R26802 VSS.n7793 VSS.n7705 1.292
R26803 VSS.n7793 VSS.n7792 1.292
R26804 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Collector VSS.n7712 1.292
R26805 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Collector VSS.n7713 1.292
R26806 VSS.n7783 VSS.n7782 1.292
R26807 VSS.n7782 VSS.n7720 1.292
R26808 VSS.n7771 VSS.n7724 1.292
R26809 VSS.n7771 VSS.n7770 1.292
R26810 VSS.n7766 VSS.n7731 1.292
R26811 VSS.n7766 VSS.n7732 1.292
R26812 VSS.n7760 VSS.n7759 1.292
R26813 VSS.n7759 VSS.n7739 1.292
R26814 VSS.n7748 VSS.n7743 1.292
R26815 VSS.n7748 VSS.n7747 1.292
R26816 VSS.n6815 sky130_asc_pnp_05v5_W3p40L3p40_1_0/xm1/Collector 1.292
R26817 VSS.n5566 VSS.n5565 1.292
R26818 VSS.n5565 VSS.n5418 1.292
R26819 VSS.n5554 VSS.n5420 1.292
R26820 VSS.n5554 VSS.n5553 1.292
R26821 VSS.n5549 VSS.n5428 1.292
R26822 VSS.n5549 VSS.n5429 1.292
R26823 VSS.n5543 VSS.n5542 1.292
R26824 VSS.n5542 VSS.n5436 1.292
R26825 VSS.n5531 VSS.n5440 1.292
R26826 VSS.n5531 VSS.n5530 1.292
R26827 VSS.n5526 VSS.n5447 1.292
R26828 VSS.n5526 VSS.n5448 1.292
R26829 VSS.n5520 sky130_asc_pnp_05v5_W3p40L3p40_8_2/xm1/Collector 1.292
R26830 sky130_asc_pnp_05v5_W3p40L3p40_8_2/xm1/Collector VSS.n5455 1.292
R26831 VSS.n5509 VSS.n5459 1.292
R26832 VSS.n5509 VSS.n5508 1.292
R26833 VSS.n5504 VSS.n5466 1.292
R26834 VSS.n5504 VSS.n5467 1.292
R26835 VSS.n5498 VSS.n5497 1.292
R26836 VSS.n5497 VSS.n5474 1.292
R26837 VSS.n5486 VSS.n5478 1.292
R26838 VSS.n5486 VSS.n5485 1.292
R26839 VSS.n5661 VSS.n3637 1.292
R26840 VSS.n5661 VSS.n3638 1.292
R26841 VSS.n5323 VSS.n3749 1.292
R26842 VSS.n5324 VSS.n5323 1.292
R26843 VSS.n5329 VSS.n5328 1.292
R26844 VSS.n5328 VSS.n3743 1.292
R26845 VSS.n5340 VSS.n3739 1.292
R26846 VSS.n5340 VSS.n3741 1.292
R26847 VSS.n5347 VSS.n5346 1.292
R26848 VSS.n5347 VSS.n3733 1.292
R26849 VSS.n5358 VSS.n3728 1.292
R26850 VSS.n5359 VSS.n5358 1.292
R26851 VSS.n5364 VSS.n5363 1.292
R26852 VSS.n5363 VSS.n3722 1.292
R26853 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector VSS.n3718 1.292
R26854 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector VSS.n3720 1.292
R26855 VSS.n5381 VSS.n5380 1.292
R26856 VSS.n5381 VSS.n3712 1.292
R26857 VSS.n5392 VSS.n3707 1.292
R26858 VSS.n5393 VSS.n5392 1.292
R26859 VSS.n5398 VSS.n5397 1.292
R26860 VSS.n5397 VSS.n3699 1.292
R26861 VSS.n3700 VSS.n3697 1.292
R26862 VSS.n5410 VSS.n3697 1.292
R26863 VSS.n5573 VSS.n3692 1.292
R26864 VSS.n5573 VSS.n3690 1.292
R26865 VSS.n5220 VSS.n5219 1.292
R26866 VSS.n5219 VSS.n5061 1.292
R26867 VSS.n5208 VSS.n5063 1.292
R26868 VSS.n5208 VSS.n5207 1.292
R26869 VSS.n5203 VSS.n5071 1.292
R26870 VSS.n5203 VSS.n5072 1.292
R26871 VSS.n5197 VSS.n5196 1.292
R26872 VSS.n5196 VSS.n5079 1.292
R26873 VSS.n5185 VSS.n5083 1.292
R26874 VSS.n5185 VSS.n5184 1.292
R26875 VSS.n5180 VSS.n5090 1.292
R26876 VSS.n5180 VSS.n5091 1.292
R26877 VSS.n5174 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector 1.292
R26878 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector VSS.n5098 1.292
R26879 VSS.n5163 VSS.n5102 1.292
R26880 VSS.n5163 VSS.n5162 1.292
R26881 VSS.n5158 VSS.n5109 1.292
R26882 VSS.n5158 VSS.n5110 1.292
R26883 VSS.n5152 VSS.n5151 1.292
R26884 VSS.n5151 VSS.n5117 1.292
R26885 VSS.n5140 VSS.n5121 1.292
R26886 VSS.n5140 VSS.n5139 1.292
R26887 VSS.n5135 VSS.n5129 1.292
R26888 VSS.n5135 VSS.n5130 1.292
R26889 VSS.n4966 VSS.n3890 1.292
R26890 VSS.n4967 VSS.n4966 1.292
R26891 VSS.n4972 VSS.n4971 1.292
R26892 VSS.n4971 VSS.n3884 1.292
R26893 VSS.n4983 VSS.n3880 1.292
R26894 VSS.n4983 VSS.n3882 1.292
R26895 VSS.n4990 VSS.n4989 1.292
R26896 VSS.n4990 VSS.n3874 1.292
R26897 VSS.n5001 VSS.n3869 1.292
R26898 VSS.n5002 VSS.n5001 1.292
R26899 VSS.n5007 VSS.n5006 1.292
R26900 VSS.n5006 VSS.n3863 1.292
R26901 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector VSS.n3859 1.292
R26902 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector VSS.n3861 1.292
R26903 VSS.n5024 VSS.n5023 1.292
R26904 VSS.n5024 VSS.n3853 1.292
R26905 VSS.n5035 VSS.n3848 1.292
R26906 VSS.n5036 VSS.n5035 1.292
R26907 VSS.n5041 VSS.n5040 1.292
R26908 VSS.n5040 VSS.n3840 1.292
R26909 VSS.n3841 VSS.n3838 1.292
R26910 VSS.n5053 VSS.n3838 1.292
R26911 VSS.n5227 VSS.n3833 1.292
R26912 VSS.n5227 VSS.n3831 1.292
R26913 VSS.n4863 VSS.n4862 1.292
R26914 VSS.n4862 VSS.n4704 1.292
R26915 VSS.n4851 VSS.n4706 1.292
R26916 VSS.n4851 VSS.n4850 1.292
R26917 VSS.n4846 VSS.n4714 1.292
R26918 VSS.n4846 VSS.n4715 1.292
R26919 VSS.n4840 VSS.n4839 1.292
R26920 VSS.n4839 VSS.n4722 1.292
R26921 VSS.n4828 VSS.n4726 1.292
R26922 VSS.n4828 VSS.n4827 1.292
R26923 VSS.n4823 VSS.n4733 1.292
R26924 VSS.n4823 VSS.n4734 1.292
R26925 VSS.n4817 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector 1.292
R26926 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector VSS.n4741 1.292
R26927 VSS.n4806 VSS.n4745 1.292
R26928 VSS.n4806 VSS.n4805 1.292
R26929 VSS.n4801 VSS.n4752 1.292
R26930 VSS.n4801 VSS.n4753 1.292
R26931 VSS.n4795 VSS.n4794 1.292
R26932 VSS.n4794 VSS.n4760 1.292
R26933 VSS.n4783 VSS.n4764 1.292
R26934 VSS.n4783 VSS.n4782 1.292
R26935 VSS.n4778 VSS.n4772 1.292
R26936 VSS.n4778 VSS.n4773 1.292
R26937 VSS.n4609 VSS.n4031 1.292
R26938 VSS.n4610 VSS.n4609 1.292
R26939 VSS.n4615 VSS.n4614 1.292
R26940 VSS.n4614 VSS.n4025 1.292
R26941 VSS.n4626 VSS.n4021 1.292
R26942 VSS.n4626 VSS.n4023 1.292
R26943 VSS.n4633 VSS.n4632 1.292
R26944 VSS.n4633 VSS.n4015 1.292
R26945 VSS.n4644 VSS.n4010 1.292
R26946 VSS.n4645 VSS.n4644 1.292
R26947 VSS.n4650 VSS.n4649 1.292
R26948 VSS.n4649 VSS.n4004 1.292
R26949 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector VSS.n4000 1.292
R26950 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector VSS.n4002 1.292
R26951 VSS.n4667 VSS.n4666 1.292
R26952 VSS.n4667 VSS.n3994 1.292
R26953 VSS.n4678 VSS.n3989 1.292
R26954 VSS.n4679 VSS.n4678 1.292
R26955 VSS.n4684 VSS.n4683 1.292
R26956 VSS.n4683 VSS.n3981 1.292
R26957 VSS.n3982 VSS.n3979 1.292
R26958 VSS.n4696 VSS.n3979 1.292
R26959 VSS.n4870 VSS.n3974 1.292
R26960 VSS.n4870 VSS.n3972 1.292
R26961 VSS.n4506 VSS.n4505 1.292
R26962 VSS.n4505 VSS.n4347 1.292
R26963 VSS.n4494 VSS.n4349 1.292
R26964 VSS.n4494 VSS.n4493 1.292
R26965 VSS.n4489 VSS.n4357 1.292
R26966 VSS.n4489 VSS.n4358 1.292
R26967 VSS.n4483 VSS.n4482 1.292
R26968 VSS.n4482 VSS.n4365 1.292
R26969 VSS.n4471 VSS.n4369 1.292
R26970 VSS.n4471 VSS.n4470 1.292
R26971 VSS.n4466 VSS.n4376 1.292
R26972 VSS.n4466 VSS.n4377 1.292
R26973 VSS.n4460 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector 1.292
R26974 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector VSS.n4384 1.292
R26975 VSS.n4449 VSS.n4388 1.292
R26976 VSS.n4449 VSS.n4448 1.292
R26977 VSS.n4444 VSS.n4395 1.292
R26978 VSS.n4444 VSS.n4396 1.292
R26979 VSS.n4438 VSS.n4437 1.292
R26980 VSS.n4437 VSS.n4403 1.292
R26981 VSS.n4426 VSS.n4407 1.292
R26982 VSS.n4426 VSS.n4425 1.292
R26983 VSS.n4421 VSS.n4415 1.292
R26984 VSS.n4421 VSS.n4416 1.292
R26985 VSS.n4252 VSS.n4172 1.292
R26986 VSS.n4253 VSS.n4252 1.292
R26987 VSS.n4258 VSS.n4257 1.292
R26988 VSS.n4257 VSS.n4166 1.292
R26989 VSS.n4269 VSS.n4162 1.292
R26990 VSS.n4269 VSS.n4164 1.292
R26991 VSS.n4276 VSS.n4275 1.292
R26992 VSS.n4276 VSS.n4156 1.292
R26993 VSS.n4287 VSS.n4151 1.292
R26994 VSS.n4288 VSS.n4287 1.292
R26995 VSS.n4293 VSS.n4292 1.292
R26996 VSS.n4292 VSS.n4145 1.292
R26997 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Collector VSS.n4141 1.292
R26998 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Collector VSS.n4143 1.292
R26999 VSS.n4310 VSS.n4309 1.292
R27000 VSS.n4310 VSS.n4135 1.292
R27001 VSS.n4321 VSS.n4130 1.292
R27002 VSS.n4322 VSS.n4321 1.292
R27003 VSS.n4327 VSS.n4326 1.292
R27004 VSS.n4326 VSS.n4122 1.292
R27005 VSS.n4123 VSS.n4120 1.292
R27006 VSS.n4339 VSS.n4120 1.292
R27007 VSS.n4513 VSS.n4115 1.292
R27008 VSS.n4513 VSS.n4113 1.292
R27009 VSS.n2962 VSS.n2802 1.292
R27010 VSS.n2962 VSS.n2803 1.292
R27011 VSS.n2956 VSS.n2955 1.292
R27012 VSS.n2955 VSS.n2812 1.292
R27013 VSS.n2944 VSS.n2816 1.292
R27014 VSS.n2944 VSS.n2943 1.292
R27015 VSS.n2939 VSS.n2823 1.292
R27016 VSS.n2939 VSS.n2824 1.292
R27017 VSS.n2933 VSS.n2932 1.292
R27018 VSS.n2932 VSS.n2831 1.292
R27019 VSS.n2921 VSS.n2835 1.292
R27020 VSS.n2921 VSS.n2920 1.292
R27021 sky130_asc_pnp_05v5_W3p40L3p40_7_0/xm1/Collector VSS.n2842 1.292
R27022 sky130_asc_pnp_05v5_W3p40L3p40_7_0/xm1/Collector VSS.n2843 1.292
R27023 VSS.n2911 VSS.n2910 1.292
R27024 VSS.n2910 VSS.n2850 1.292
R27025 VSS.n2899 VSS.n2854 1.292
R27026 VSS.n2899 VSS.n2898 1.292
R27027 VSS.n2894 VSS.n2861 1.292
R27028 VSS.n2894 VSS.n2862 1.292
R27029 VSS.n2888 VSS.n2887 1.292
R27030 VSS.n2887 VSS.n2869 1.292
R27031 VSS.n2877 VSS.n2876 1.292
R27032 VSS.n2876 VSS.n2875 1.292
R27033 VSS.n2699 VSS.n2698 1.292
R27034 VSS.n2698 VSS.n1371 1.292
R27035 VSS.n2710 VSS.n1367 1.292
R27036 VSS.n2710 VSS.n1369 1.292
R27037 VSS.n2717 VSS.n2716 1.292
R27038 VSS.n2717 VSS.n1361 1.292
R27039 VSS.n2728 VSS.n1356 1.292
R27040 VSS.n2729 VSS.n2728 1.292
R27041 VSS.n2734 VSS.n2733 1.292
R27042 VSS.n2733 VSS.n1350 1.292
R27043 VSS.n2745 VSS.n1346 1.292
R27044 VSS.n2745 VSS.n1348 1.292
R27045 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector VSS.n2751 1.292
R27046 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Collector VSS.n1340 1.292
R27047 VSS.n2762 VSS.n1335 1.292
R27048 VSS.n2763 VSS.n2762 1.292
R27049 VSS.n2768 VSS.n2767 1.292
R27050 VSS.n2767 VSS.n1329 1.292
R27051 VSS.n2779 VSS.n1325 1.292
R27052 VSS.n2779 VSS.n1327 1.292
R27053 VSS.n2786 VSS.n2785 1.292
R27054 VSS.n2786 VSS.n1319 1.292
R27055 VSS.n2797 VSS.n1315 1.292
R27056 VSS.n2798 VSS.n2797 1.292
R27057 VSS.n2470 VSS.n2326 1.292
R27058 VSS.n2470 VSS.n2327 1.292
R27059 VSS.n2464 VSS.n2463 1.292
R27060 VSS.n2463 VSS.n2337 1.292
R27061 VSS.n2452 VSS.n2341 1.292
R27062 VSS.n2452 VSS.n2451 1.292
R27063 VSS.n2447 VSS.n2348 1.292
R27064 VSS.n2447 VSS.n2349 1.292
R27065 VSS.n2441 VSS.n2440 1.292
R27066 VSS.n2440 VSS.n2356 1.292
R27067 VSS.n2429 VSS.n2360 1.292
R27068 VSS.n2429 VSS.n2428 1.292
R27069 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector VSS.n2367 1.292
R27070 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Collector VSS.n2368 1.292
R27071 VSS.n2419 VSS.n2418 1.292
R27072 VSS.n2418 VSS.n2375 1.292
R27073 VSS.n2407 VSS.n2379 1.292
R27074 VSS.n2407 VSS.n2406 1.292
R27075 VSS.n2402 VSS.n2386 1.292
R27076 VSS.n2402 VSS.n2387 1.292
R27077 VSS.n2396 VSS.n2395 1.292
R27078 VSS.n2395 VSS.n1380 1.292
R27079 VSS.n1381 VSS.n1378 1.292
R27080 VSS.n2693 VSS.n1378 1.292
R27081 VSS.n2562 VSS.n2215 1.292
R27082 VSS.n2562 VSS.n2216 1.292
R27083 VSS.n2556 VSS.n2555 1.292
R27084 VSS.n2555 VSS.n2225 1.292
R27085 VSS.n2544 VSS.n2229 1.292
R27086 VSS.n2544 VSS.n2543 1.292
R27087 VSS.n2539 VSS.n2236 1.292
R27088 VSS.n2539 VSS.n2237 1.292
R27089 VSS.n2533 VSS.n2532 1.292
R27090 VSS.n2532 VSS.n2244 1.292
R27091 VSS.n2521 VSS.n2248 1.292
R27092 VSS.n2521 VSS.n2520 1.292
R27093 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector VSS.n2255 1.292
R27094 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Collector VSS.n2256 1.292
R27095 VSS.n2511 VSS.n2510 1.292
R27096 VSS.n2510 VSS.n2263 1.292
R27097 VSS.n2499 VSS.n2267 1.292
R27098 VSS.n2499 VSS.n2498 1.292
R27099 VSS.n2494 VSS.n2274 1.292
R27100 VSS.n2494 VSS.n2275 1.292
R27101 VSS.n2488 VSS.n2487 1.292
R27102 VSS.n2487 VSS.n2282 1.292
R27103 VSS.n2476 VSS.n2286 1.292
R27104 VSS.n2476 VSS.n2475 1.292
R27105 VSS.n2119 VSS.n2118 1.292
R27106 VSS.n2119 VSS.n1538 1.292
R27107 VSS.n2130 VSS.n1533 1.292
R27108 VSS.n2131 VSS.n2130 1.292
R27109 VSS.n2136 VSS.n2135 1.292
R27110 VSS.n2135 VSS.n1527 1.292
R27111 VSS.n2147 VSS.n1523 1.292
R27112 VSS.n2147 VSS.n1525 1.292
R27113 VSS.n2154 VSS.n2153 1.292
R27114 VSS.n2154 VSS.n1517 1.292
R27115 VSS.n2165 VSS.n1512 1.292
R27116 VSS.n2166 VSS.n2165 1.292
R27117 VSS.n2170 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector 1.292
R27118 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Collector VSS.n1506 1.292
R27119 VSS.n2181 VSS.n1502 1.292
R27120 VSS.n2181 VSS.n1504 1.292
R27121 VSS.n2188 VSS.n2187 1.292
R27122 VSS.n2188 VSS.n1496 1.292
R27123 VSS.n2199 VSS.n1491 1.292
R27124 VSS.n2200 VSS.n2199 1.292
R27125 VSS.n2205 VSS.n2204 1.292
R27126 VSS.n2204 VSS.n1485 1.292
R27127 VSS.n2569 VSS.n1482 1.292
R27128 VSS.n2569 VSS.n1483 1.292
R27129 VSS.n1869 VSS.n1717 1.292
R27130 VSS.n1869 VSS.n1718 1.292
R27131 VSS.n1863 VSS.n1862 1.292
R27132 VSS.n1862 VSS.n1728 1.292
R27133 VSS.n1851 VSS.n1732 1.292
R27134 VSS.n1851 VSS.n1850 1.292
R27135 VSS.n1846 VSS.n1739 1.292
R27136 VSS.n1846 VSS.n1740 1.292
R27137 VSS.n1840 VSS.n1839 1.292
R27138 VSS.n1839 VSS.n1747 1.292
R27139 VSS.n1828 VSS.n1751 1.292
R27140 VSS.n1828 VSS.n1827 1.292
R27141 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector VSS.n1758 1.292
R27142 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Collector VSS.n1759 1.292
R27143 VSS.n1818 VSS.n1817 1.292
R27144 VSS.n1817 VSS.n1766 1.292
R27145 VSS.n1806 VSS.n1770 1.292
R27146 VSS.n1806 VSS.n1805 1.292
R27147 VSS.n1801 VSS.n1777 1.292
R27148 VSS.n1801 VSS.n1778 1.292
R27149 VSS.n1795 VSS.n1794 1.292
R27150 VSS.n1794 VSS.n1789 1.292
R27151 VSS.n2111 VSS.n1546 1.292
R27152 VSS.n2111 VSS.n1547 1.292
R27153 VSS.n1962 VSS.n1961 1.292
R27154 VSS.n1961 VSS.n1609 1.292
R27155 VSS.n1955 VSS.n1954 1.292
R27156 VSS.n1954 VSS.n1615 1.292
R27157 VSS.n1943 VSS.n1620 1.292
R27158 VSS.n1943 VSS.n1942 1.292
R27159 VSS.n1938 VSS.n1627 1.292
R27160 VSS.n1938 VSS.n1628 1.292
R27161 VSS.n1932 VSS.n1931 1.292
R27162 VSS.n1931 VSS.n1635 1.292
R27163 VSS.n1920 VSS.n1639 1.292
R27164 VSS.n1920 VSS.n1919 1.292
R27165 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector VSS.n1646 1.292
R27166 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Collector VSS.n1647 1.292
R27167 VSS.n1910 VSS.n1909 1.292
R27168 VSS.n1909 VSS.n1654 1.292
R27169 VSS.n1898 VSS.n1658 1.292
R27170 VSS.n1898 VSS.n1897 1.292
R27171 VSS.n1893 VSS.n1665 1.292
R27172 VSS.n1893 VSS.n1666 1.292
R27173 VSS.n1887 VSS.n1886 1.292
R27174 VSS.n1886 VSS.n1673 1.292
R27175 VSS.n1875 VSS.n1677 1.292
R27176 VSS.n1875 VSS.n1874 1.292
R27177 VSS.n15670 VSS.n15669 1.28
R27178 VSS.n15892 VSS.n15891 1.28
R27179 VSS.n15454 VSS.n14136 1.28
R27180 VSS.n15083 VSS.n15082 1.28
R27181 VSS.n15334 VSS.n14236 1.28
R27182 VSS.n14865 VSS.n14864 1.28
R27183 VSS.n14474 VSS.n14473 1.28
R27184 VSS.n12104 VSS.n11984 1.28
R27185 VSS.n12409 VSS.n11541 1.28
R27186 VSS.n11804 VSS.n11775 1.28
R27187 VSS.n13398 VSS.n13397 1.28
R27188 VSS.n13315 VSS.n13314 1.28
R27189 VSS.n13149 VSS.n13148 1.28
R27190 VSS.n13066 VSS.n13065 1.28
R27191 VSS.n8853 VSS.n6968 1.28
R27192 VSS.n8764 VSS.n7254 1.28
R27193 VSS.n8631 VSS.n7324 1.28
R27194 VSS.n8542 VSS.n7394 1.28
R27195 VSS.n8273 VSS.n7464 1.28
R27196 VSS.n8184 VSS.n7534 1.28
R27197 VSS.n7915 VSS.n7604 1.28
R27198 VSS.n5579 VSS.n5578 1.28
R27199 VSS.n5316 VSS.n5315 1.28
R27200 VSS.n5233 VSS.n5232 1.28
R27201 VSS.n4959 VSS.n4958 1.28
R27202 VSS.n4876 VSS.n4875 1.28
R27203 VSS.n4602 VSS.n4601 1.28
R27204 VSS.n4519 VSS.n4518 1.28
R27205 VSS.n2966 VSS.n2965 1.28
R27206 VSS.n2695 VSS.n1377 1.28
R27207 VSS.n2324 VSS.n2323 1.28
R27208 VSS.n2575 VSS.n1477 1.28
R27209 VSS.n2106 VSS.n2105 1.28
R27210 VSS.n1715 VSS.n1714 1.28
R27211 VSS.n6900 VSS.n6881 1.245
R27212 VSS.n17328 VSS.n17312 1.244
R27213 VSS.n17391 VSS.n16051 1.244
R27214 VSS.n17394 VSS.n17393 1.244
R27215 VSS.n17396 VSS.n16048 1.244
R27216 VSS.n17457 VSS.n17456 1.244
R27217 VSS.n17450 VSS.n16049 1.244
R27218 VSS.n17449 VSS.n17447 1.244
R27219 VSS.n17444 VSS.n17400 1.244
R27220 VSS.n17404 VSS.n17403 1.244
R27221 VSS.n17438 VSS.n17437 1.244
R27222 VSS.n17408 VSS.n17406 1.244
R27223 VSS.n17434 sky130_asc_pnp_05v5_W3p40L3p40_8_3/xm1/Base 1.244
R27224 VSS.n17432 VSS.n17431 1.244
R27225 VSS.n17412 VSS.n17410 1.244
R27226 VSS.n17426 VSS.n17425 1.244
R27227 VSS.n17415 VSS.n17414 1.244
R27228 VSS.n17420 VSS.n17419 1.244
R27229 VSS.n17417 VSS.n16027 1.244
R27230 VSS.n17331 VSS.n16028 1.244
R27231 VSS.n17225 VSS.n17223 1.244
R27232 VSS.n17227 VSS.n16091 1.244
R27233 VSS.n17301 VSS.n17300 1.244
R27234 VSS.n17294 VSS.n16092 1.244
R27235 VSS.n17293 VSS.n17291 1.244
R27236 VSS.n17288 VSS.n17231 1.244
R27237 VSS.n17235 VSS.n17234 1.244
R27238 VSS.n17282 VSS.n17281 1.244
R27239 VSS.n17239 VSS.n17237 1.244
R27240 VSS.n17276 VSS.n17275 1.244
R27241 VSS.n17243 VSS.n17241 1.244
R27242 VSS.n17272 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Base 1.244
R27243 VSS.n17270 VSS.n17269 1.244
R27244 VSS.n17247 VSS.n17245 1.244
R27245 VSS.n17264 VSS.n17263 1.244
R27246 VSS.n17248 VSS.n16081 1.244
R27247 VSS.n17259 VSS.n17258 1.244
R27248 VSS.n17253 VSS.n17251 1.244
R27249 VSS.n17254 VSS.n16053 1.244
R27250 VSS.n17135 VSS.n17133 1.244
R27251 VSS.n17137 VSS.n16181 1.244
R27252 VSS.n17211 VSS.n17210 1.244
R27253 VSS.n17204 VSS.n16182 1.244
R27254 VSS.n17203 VSS.n17201 1.244
R27255 VSS.n17198 VSS.n17141 1.244
R27256 VSS.n17145 VSS.n17144 1.244
R27257 VSS.n17192 VSS.n17191 1.244
R27258 VSS.n17149 VSS.n17147 1.244
R27259 VSS.n17186 VSS.n17185 1.244
R27260 VSS.n17153 VSS.n17151 1.244
R27261 VSS.n17182 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Base 1.244
R27262 VSS.n17180 VSS.n17179 1.244
R27263 VSS.n17157 VSS.n17155 1.244
R27264 VSS.n17174 VSS.n17173 1.244
R27265 VSS.n17158 VSS.n16171 1.244
R27266 VSS.n17169 VSS.n17168 1.244
R27267 VSS.n17163 VSS.n17161 1.244
R27268 VSS.n17164 VSS.n16143 1.244
R27269 VSS.n17045 VSS.n17043 1.244
R27270 VSS.n17047 VSS.n16271 1.244
R27271 VSS.n17121 VSS.n17120 1.244
R27272 VSS.n17114 VSS.n16272 1.244
R27273 VSS.n17113 VSS.n17111 1.244
R27274 VSS.n17108 VSS.n17051 1.244
R27275 VSS.n17055 VSS.n17054 1.244
R27276 VSS.n17102 VSS.n17101 1.244
R27277 VSS.n17059 VSS.n17057 1.244
R27278 VSS.n17096 VSS.n17095 1.244
R27279 VSS.n17063 VSS.n17061 1.244
R27280 VSS.n17092 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Base 1.244
R27281 VSS.n17090 VSS.n17089 1.244
R27282 VSS.n17067 VSS.n17065 1.244
R27283 VSS.n17084 VSS.n17083 1.244
R27284 VSS.n17068 VSS.n16261 1.244
R27285 VSS.n17079 VSS.n17078 1.244
R27286 VSS.n17073 VSS.n17071 1.244
R27287 VSS.n17074 VSS.n16233 1.244
R27288 VSS.n16955 VSS.n16953 1.244
R27289 VSS.n16957 VSS.n16361 1.244
R27290 VSS.n17031 VSS.n17030 1.244
R27291 VSS.n17024 VSS.n16362 1.244
R27292 VSS.n17023 VSS.n17021 1.244
R27293 VSS.n17018 VSS.n16961 1.244
R27294 VSS.n16965 VSS.n16964 1.244
R27295 VSS.n17012 VSS.n17011 1.244
R27296 VSS.n16969 VSS.n16967 1.244
R27297 VSS.n17006 VSS.n17005 1.244
R27298 VSS.n16973 VSS.n16971 1.244
R27299 VSS.n17002 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Base 1.244
R27300 VSS.n17000 VSS.n16999 1.244
R27301 VSS.n16977 VSS.n16975 1.244
R27302 VSS.n16994 VSS.n16993 1.244
R27303 VSS.n16978 VSS.n16351 1.244
R27304 VSS.n16989 VSS.n16988 1.244
R27305 VSS.n16983 VSS.n16981 1.244
R27306 VSS.n16984 VSS.n16323 1.244
R27307 VSS.n16865 VSS.n16863 1.244
R27308 VSS.n16867 VSS.n16451 1.244
R27309 VSS.n16941 VSS.n16940 1.244
R27310 VSS.n16934 VSS.n16452 1.244
R27311 VSS.n16933 VSS.n16931 1.244
R27312 VSS.n16928 VSS.n16871 1.244
R27313 VSS.n16875 VSS.n16874 1.244
R27314 VSS.n16922 VSS.n16921 1.244
R27315 VSS.n16879 VSS.n16877 1.244
R27316 VSS.n16916 VSS.n16915 1.244
R27317 VSS.n16883 VSS.n16881 1.244
R27318 VSS.n16912 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Base 1.244
R27319 VSS.n16910 VSS.n16909 1.244
R27320 VSS.n16887 VSS.n16885 1.244
R27321 VSS.n16904 VSS.n16903 1.244
R27322 VSS.n16888 VSS.n16441 1.244
R27323 VSS.n16899 VSS.n16898 1.244
R27324 VSS.n16893 VSS.n16891 1.244
R27325 VSS.n16894 VSS.n16413 1.244
R27326 VSS.n16775 VSS.n16773 1.244
R27327 VSS.n16777 VSS.n16541 1.244
R27328 VSS.n16851 VSS.n16850 1.244
R27329 VSS.n16844 VSS.n16542 1.244
R27330 VSS.n16843 VSS.n16841 1.244
R27331 VSS.n16838 VSS.n16781 1.244
R27332 VSS.n16785 VSS.n16784 1.244
R27333 VSS.n16832 VSS.n16831 1.244
R27334 VSS.n16789 VSS.n16787 1.244
R27335 VSS.n16826 VSS.n16825 1.244
R27336 VSS.n16793 VSS.n16791 1.244
R27337 VSS.n16822 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Base 1.244
R27338 VSS.n16820 VSS.n16819 1.244
R27339 VSS.n16797 VSS.n16795 1.244
R27340 VSS.n16814 VSS.n16813 1.244
R27341 VSS.n16798 VSS.n16531 1.244
R27342 VSS.n16809 VSS.n16808 1.244
R27343 VSS.n16803 VSS.n16801 1.244
R27344 VSS.n16804 VSS.n16503 1.244
R27345 VSS.n16685 VSS.n16683 1.244
R27346 VSS.n16687 VSS.n16631 1.244
R27347 VSS.n16761 VSS.n16760 1.244
R27348 VSS.n16754 VSS.n16632 1.244
R27349 VSS.n16753 VSS.n16751 1.244
R27350 VSS.n16748 VSS.n16691 1.244
R27351 VSS.n16695 VSS.n16694 1.244
R27352 VSS.n16742 VSS.n16741 1.244
R27353 VSS.n16699 VSS.n16697 1.244
R27354 VSS.n16736 VSS.n16735 1.244
R27355 VSS.n16703 VSS.n16701 1.244
R27356 VSS.n16732 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Base 1.244
R27357 VSS.n16730 VSS.n16729 1.244
R27358 VSS.n16707 VSS.n16705 1.244
R27359 VSS.n16724 VSS.n16723 1.244
R27360 VSS.n16708 VSS.n16621 1.244
R27361 VSS.n16719 VSS.n16718 1.244
R27362 VSS.n16713 VSS.n16711 1.244
R27363 VSS.n16714 VSS.n16593 1.244
R27364 VSS.n11152 VSS.n11151 1.244
R27365 VSS.n11154 VSS.n11098 1.244
R27366 VSS.n11229 VSS.n11228 1.244
R27367 VSS.n11222 VSS.n11099 1.244
R27368 VSS.n11221 VSS.n11219 1.244
R27369 VSS.n11216 VSS.n11158 1.244
R27370 VSS.n11162 VSS.n11161 1.244
R27371 VSS.n11210 VSS.n11209 1.244
R27372 VSS.n11166 VSS.n11164 1.244
R27373 VSS.n11204 VSS.n11203 1.244
R27374 VSS.n11170 VSS.n11168 1.244
R27375 VSS.n11200 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Base 1.244
R27376 VSS.n11198 VSS.n11197 1.244
R27377 VSS.n11171 VSS.n11088 1.244
R27378 VSS.n11193 VSS.n11192 1.244
R27379 VSS.n11176 VSS.n11174 1.244
R27380 VSS.n11187 VSS.n11186 1.244
R27381 VSS.n11181 VSS.n11177 1.244
R27382 VSS.n11182 VSS.n11060 1.244
R27383 VSS.n11242 VSS.n11241 1.244
R27384 VSS.n11244 VSS.n11008 1.244
R27385 VSS.n11319 VSS.n11318 1.244
R27386 VSS.n11312 VSS.n11009 1.244
R27387 VSS.n11311 VSS.n11309 1.244
R27388 VSS.n11306 VSS.n11248 1.244
R27389 VSS.n11252 VSS.n11251 1.244
R27390 VSS.n11300 VSS.n11299 1.244
R27391 VSS.n11256 VSS.n11254 1.244
R27392 VSS.n11294 VSS.n11293 1.244
R27393 VSS.n11260 VSS.n11258 1.244
R27394 VSS.n11290 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Base 1.244
R27395 VSS.n11288 VSS.n11287 1.244
R27396 VSS.n11261 VSS.n10998 1.244
R27397 VSS.n11283 VSS.n11282 1.244
R27398 VSS.n11266 VSS.n11264 1.244
R27399 VSS.n11277 VSS.n11276 1.244
R27400 VSS.n11271 VSS.n11267 1.244
R27401 VSS.n11272 VSS.n10970 1.244
R27402 VSS.n11332 VSS.n11331 1.244
R27403 VSS.n11334 VSS.n10918 1.244
R27404 VSS.n11409 VSS.n11408 1.244
R27405 VSS.n11402 VSS.n10919 1.244
R27406 VSS.n11401 VSS.n11399 1.244
R27407 VSS.n11396 VSS.n11338 1.244
R27408 VSS.n11342 VSS.n11341 1.244
R27409 VSS.n11390 VSS.n11389 1.244
R27410 VSS.n11346 VSS.n11344 1.244
R27411 VSS.n11384 VSS.n11383 1.244
R27412 VSS.n11350 VSS.n11348 1.244
R27413 VSS.n11380 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Base 1.244
R27414 VSS.n11378 VSS.n11377 1.244
R27415 VSS.n11351 VSS.n10908 1.244
R27416 VSS.n11373 VSS.n11372 1.244
R27417 VSS.n11356 VSS.n11354 1.244
R27418 VSS.n11367 VSS.n11366 1.244
R27419 VSS.n11361 VSS.n11357 1.244
R27420 VSS.n11362 VSS.n10880 1.244
R27421 VSS.n11422 VSS.n11421 1.244
R27422 VSS.n11424 VSS.n10828 1.244
R27423 VSS.n13529 VSS.n13528 1.244
R27424 VSS.n13522 VSS.n10829 1.244
R27425 VSS.n13521 VSS.n13519 1.244
R27426 VSS.n13516 VSS.n11428 1.244
R27427 VSS.n13461 VSS.n13460 1.244
R27428 VSS.n13509 VSS.n13508 1.244
R27429 VSS.n13465 VSS.n13463 1.244
R27430 VSS.n13503 VSS.n13502 1.244
R27431 VSS.n13469 VSS.n13467 1.244
R27432 VSS.n13499 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Base 1.244
R27433 VSS.n13497 VSS.n13496 1.244
R27434 VSS.n13470 VSS.n10818 1.244
R27435 VSS.n13492 VSS.n13491 1.244
R27436 VSS.n13475 VSS.n13473 1.244
R27437 VSS.n13486 VSS.n13485 1.244
R27438 VSS.n13480 VSS.n13476 1.244
R27439 VSS.n13481 VSS.n10790 1.244
R27440 VSS.n13542 VSS.n13541 1.244
R27441 VSS.n13544 VSS.n10738 1.244
R27442 VSS.n13619 VSS.n13618 1.244
R27443 VSS.n13612 VSS.n10739 1.244
R27444 VSS.n13611 VSS.n13609 1.244
R27445 VSS.n13606 VSS.n13548 1.244
R27446 VSS.n13552 VSS.n13551 1.244
R27447 VSS.n13600 VSS.n13599 1.244
R27448 VSS.n13556 VSS.n13554 1.244
R27449 VSS.n13594 VSS.n13593 1.244
R27450 VSS.n13560 VSS.n13558 1.244
R27451 VSS.n13590 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Base 1.244
R27452 VSS.n13588 VSS.n13587 1.244
R27453 VSS.n13561 VSS.n10728 1.244
R27454 VSS.n13583 VSS.n13582 1.244
R27455 VSS.n13566 VSS.n13564 1.244
R27456 VSS.n13577 VSS.n13576 1.244
R27457 VSS.n13571 VSS.n13567 1.244
R27458 VSS.n13572 VSS.n10700 1.244
R27459 VSS.n13632 VSS.n13631 1.244
R27460 VSS.n13634 VSS.n10648 1.244
R27461 VSS.n13709 VSS.n13708 1.244
R27462 VSS.n13702 VSS.n10649 1.244
R27463 VSS.n13701 VSS.n13699 1.244
R27464 VSS.n13696 VSS.n13638 1.244
R27465 VSS.n13642 VSS.n13641 1.244
R27466 VSS.n13690 VSS.n13689 1.244
R27467 VSS.n13646 VSS.n13644 1.244
R27468 VSS.n13684 VSS.n13683 1.244
R27469 VSS.n13650 VSS.n13648 1.244
R27470 VSS.n13680 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Base 1.244
R27471 VSS.n13678 VSS.n13677 1.244
R27472 VSS.n13651 VSS.n10638 1.244
R27473 VSS.n13673 VSS.n13672 1.244
R27474 VSS.n13656 VSS.n13654 1.244
R27475 VSS.n13667 VSS.n13666 1.244
R27476 VSS.n13661 VSS.n13657 1.244
R27477 VSS.n13662 VSS.n10610 1.244
R27478 VSS.n13722 VSS.n13721 1.244
R27479 VSS.n13724 VSS.n10558 1.244
R27480 VSS.n13799 VSS.n13798 1.244
R27481 VSS.n13792 VSS.n10559 1.244
R27482 VSS.n13791 VSS.n13789 1.244
R27483 VSS.n13786 VSS.n13728 1.244
R27484 VSS.n13732 VSS.n13731 1.244
R27485 VSS.n13780 VSS.n13779 1.244
R27486 VSS.n13736 VSS.n13734 1.244
R27487 VSS.n13774 VSS.n13773 1.244
R27488 VSS.n13740 VSS.n13738 1.244
R27489 VSS.n13770 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Base 1.244
R27490 VSS.n13768 VSS.n13767 1.244
R27491 VSS.n13741 VSS.n10548 1.244
R27492 VSS.n13763 VSS.n13762 1.244
R27493 VSS.n13746 VSS.n13744 1.244
R27494 VSS.n13757 VSS.n13756 1.244
R27495 VSS.n13751 VSS.n13747 1.244
R27496 VSS.n13752 VSS.n10520 1.244
R27497 VSS.n13825 VSS.n13809 1.244
R27498 VSS.n13891 VSS.n10518 1.244
R27499 VSS.n13894 VSS.n13893 1.244
R27500 VSS.n13896 VSS.n10515 1.244
R27501 VSS.n13949 VSS.n13948 1.244
R27502 VSS.n13942 VSS.n10516 1.244
R27503 VSS.n13941 VSS.n13939 1.244
R27504 VSS.n13936 VSS.n13900 1.244
R27505 VSS.n13904 VSS.n13903 1.244
R27506 VSS.n13930 VSS.n13929 1.244
R27507 VSS.n13908 VSS.n13906 1.244
R27508 VSS.n13926 sky130_asc_pnp_05v5_W3p40L3p40_8_0/xm1/Base 1.244
R27509 VSS.n13924 VSS.n13923 1.244
R27510 VSS.n13912 VSS.n13910 1.244
R27511 VSS.n13918 VSS.n13917 1.244
R27512 VSS.n13915 VSS.n13913 1.244
R27513 VSS.n13958 VSS.n13957 1.244
R27514 VSS.n13956 VSS.n10494 1.244
R27515 VSS.n13830 VSS.n13828 1.244
R27516 VSS.n9158 VSS.n8983 1.244
R27517 VSS.n9039 VSS.n9036 1.244
R27518 VSS.n9038 VSS.n9032 1.244
R27519 VSS.n9047 VSS.n9044 1.244
R27520 VSS.n9046 VSS.n9030 1.244
R27521 VSS.n9055 VSS.n9052 1.244
R27522 VSS.n9054 VSS.n9028 1.244
R27523 VSS.n9063 VSS.n9060 1.244
R27524 VSS.n9062 VSS.n9026 1.244
R27525 VSS.n9071 VSS.n9068 1.244
R27526 VSS.n9070 VSS.n9024 1.244
R27527 sky130_asc_pnp_05v5_W3p40L3p40_8_1/xm1/Base VSS.n9075 1.244
R27528 VSS.n9079 VSS.n9076 1.244
R27529 VSS.n9078 VSS.n9022 1.244
R27530 VSS.n9087 VSS.n9084 1.244
R27531 VSS.n9086 VSS.n9020 1.244
R27532 VSS.n9095 VSS.n9092 1.244
R27533 VSS.n9094 VSS.n9017 1.244
R27534 VSS.n9149 VSS.n9018 1.244
R27535 VSS.n10180 VSS.n10178 1.244
R27536 VSS.n10182 VSS.n9226 1.244
R27537 VSS.n10256 VSS.n10255 1.244
R27538 VSS.n10249 VSS.n9227 1.244
R27539 VSS.n10248 VSS.n10246 1.244
R27540 VSS.n10243 VSS.n10186 1.244
R27541 VSS.n10190 VSS.n10189 1.244
R27542 VSS.n10237 VSS.n10236 1.244
R27543 VSS.n10194 VSS.n10192 1.244
R27544 VSS.n10231 VSS.n10230 1.244
R27545 VSS.n10198 VSS.n10196 1.244
R27546 VSS.n10227 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Base 1.244
R27547 VSS.n10225 VSS.n10224 1.244
R27548 VSS.n10202 VSS.n10200 1.244
R27549 VSS.n10219 VSS.n10218 1.244
R27550 VSS.n10203 VSS.n9216 1.244
R27551 VSS.n10214 VSS.n10213 1.244
R27552 VSS.n10208 VSS.n10206 1.244
R27553 VSS.n10209 VSS.n9188 1.244
R27554 VSS.n10090 VSS.n10088 1.244
R27555 VSS.n10092 VSS.n9316 1.244
R27556 VSS.n10166 VSS.n10165 1.244
R27557 VSS.n10159 VSS.n9317 1.244
R27558 VSS.n10158 VSS.n10156 1.244
R27559 VSS.n10153 VSS.n10096 1.244
R27560 VSS.n10100 VSS.n10099 1.244
R27561 VSS.n10147 VSS.n10146 1.244
R27562 VSS.n10104 VSS.n10102 1.244
R27563 VSS.n10141 VSS.n10140 1.244
R27564 VSS.n10108 VSS.n10106 1.244
R27565 VSS.n10137 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Base 1.244
R27566 VSS.n10135 VSS.n10134 1.244
R27567 VSS.n10112 VSS.n10110 1.244
R27568 VSS.n10129 VSS.n10128 1.244
R27569 VSS.n10113 VSS.n9306 1.244
R27570 VSS.n10124 VSS.n10123 1.244
R27571 VSS.n10118 VSS.n10116 1.244
R27572 VSS.n10119 VSS.n9278 1.244
R27573 VSS.n10000 VSS.n9998 1.244
R27574 VSS.n10002 VSS.n9406 1.244
R27575 VSS.n10076 VSS.n10075 1.244
R27576 VSS.n10069 VSS.n9407 1.244
R27577 VSS.n10068 VSS.n10066 1.244
R27578 VSS.n10063 VSS.n10006 1.244
R27579 VSS.n10010 VSS.n10009 1.244
R27580 VSS.n10057 VSS.n10056 1.244
R27581 VSS.n10014 VSS.n10012 1.244
R27582 VSS.n10051 VSS.n10050 1.244
R27583 VSS.n10018 VSS.n10016 1.244
R27584 VSS.n10047 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Base 1.244
R27585 VSS.n10045 VSS.n10044 1.244
R27586 VSS.n10022 VSS.n10020 1.244
R27587 VSS.n10039 VSS.n10038 1.244
R27588 VSS.n10023 VSS.n9396 1.244
R27589 VSS.n10034 VSS.n10033 1.244
R27590 VSS.n10028 VSS.n10026 1.244
R27591 VSS.n10029 VSS.n9368 1.244
R27592 VSS.n9910 VSS.n9908 1.244
R27593 VSS.n9912 VSS.n9496 1.244
R27594 VSS.n9986 VSS.n9985 1.244
R27595 VSS.n9979 VSS.n9497 1.244
R27596 VSS.n9978 VSS.n9976 1.244
R27597 VSS.n9973 VSS.n9916 1.244
R27598 VSS.n9920 VSS.n9919 1.244
R27599 VSS.n9967 VSS.n9966 1.244
R27600 VSS.n9924 VSS.n9922 1.244
R27601 VSS.n9961 VSS.n9960 1.244
R27602 VSS.n9928 VSS.n9926 1.244
R27603 VSS.n9957 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Base 1.244
R27604 VSS.n9955 VSS.n9954 1.244
R27605 VSS.n9932 VSS.n9930 1.244
R27606 VSS.n9949 VSS.n9948 1.244
R27607 VSS.n9933 VSS.n9486 1.244
R27608 VSS.n9944 VSS.n9943 1.244
R27609 VSS.n9938 VSS.n9936 1.244
R27610 VSS.n9939 VSS.n9458 1.244
R27611 VSS.n9820 VSS.n9818 1.244
R27612 VSS.n9822 VSS.n9586 1.244
R27613 VSS.n9896 VSS.n9895 1.244
R27614 VSS.n9889 VSS.n9587 1.244
R27615 VSS.n9888 VSS.n9886 1.244
R27616 VSS.n9883 VSS.n9826 1.244
R27617 VSS.n9830 VSS.n9829 1.244
R27618 VSS.n9877 VSS.n9876 1.244
R27619 VSS.n9834 VSS.n9832 1.244
R27620 VSS.n9871 VSS.n9870 1.244
R27621 VSS.n9838 VSS.n9836 1.244
R27622 VSS.n9867 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Base 1.244
R27623 VSS.n9865 VSS.n9864 1.244
R27624 VSS.n9842 VSS.n9840 1.244
R27625 VSS.n9859 VSS.n9858 1.244
R27626 VSS.n9843 VSS.n9576 1.244
R27627 VSS.n9854 VSS.n9853 1.244
R27628 VSS.n9848 VSS.n9846 1.244
R27629 VSS.n9849 VSS.n9548 1.244
R27630 VSS.n9730 VSS.n9728 1.244
R27631 VSS.n9732 VSS.n9676 1.244
R27632 VSS.n9806 VSS.n9805 1.244
R27633 VSS.n9799 VSS.n9677 1.244
R27634 VSS.n9798 VSS.n9796 1.244
R27635 VSS.n9793 VSS.n9736 1.244
R27636 VSS.n9740 VSS.n9739 1.244
R27637 VSS.n9787 VSS.n9786 1.244
R27638 VSS.n9744 VSS.n9742 1.244
R27639 VSS.n9781 VSS.n9780 1.244
R27640 VSS.n9748 VSS.n9746 1.244
R27641 VSS.n9777 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Base 1.244
R27642 VSS.n9775 VSS.n9774 1.244
R27643 VSS.n9752 VSS.n9750 1.244
R27644 VSS.n9769 VSS.n9768 1.244
R27645 VSS.n9753 VSS.n9666 1.244
R27646 VSS.n9764 VSS.n9763 1.244
R27647 VSS.n9758 VSS.n9756 1.244
R27648 VSS.n9759 VSS.n9638 1.244
R27649 VSS.n10322 VSS.n9181 1.244
R27650 VSS.n9186 VSS.n9185 1.244
R27651 VSS.n9184 VSS.n8932 1.244
R27652 VSS.n8937 VSS.n8933 1.244
R27653 VSS.n10365 VSS.n10364 1.244
R27654 VSS.n8942 VSS.n8938 1.244
R27655 VSS.n10359 VSS.n10358 1.244
R27656 VSS.n8948 VSS.n8943 1.244
R27657 VSS.n10353 VSS.n10352 1.244
R27658 VSS.n8954 VSS.n8949 1.244
R27659 VSS.n10347 VSS.n10346 1.244
R27660 VSS.n10345 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Base 1.244
R27661 VSS.n8961 VSS.n8959 1.244
R27662 VSS.n10341 VSS.n10340 1.244
R27663 VSS.n8966 VSS.n8960 1.244
R27664 VSS.n10335 VSS.n10334 1.244
R27665 VSS.n8972 VSS.n8967 1.244
R27666 VSS.n10329 VSS.n10328 1.244
R27667 VSS.n8978 VSS.n8973 1.244
R27668 VSS.n5668 VSS.n3579 1.244
R27669 VSS.n3584 VSS.n3580 1.244
R27670 VSS.n5780 VSS.n5779 1.244
R27671 VSS.n3589 VSS.n3585 1.244
R27672 VSS.n5774 VSS.n5773 1.244
R27673 VSS.n3595 VSS.n3590 1.244
R27674 VSS.n5768 VSS.n5767 1.244
R27675 VSS.n3601 VSS.n3596 1.244
R27676 VSS.n5762 VSS.n5761 1.244
R27677 VSS.n3607 VSS.n3602 1.244
R27678 VSS.n5756 VSS.n5755 1.244
R27679 VSS.n5754 sky130_asc_pnp_05v5_W3p40L3p40_8_2/xm1/Base 1.244
R27680 VSS.n3614 VSS.n3612 1.244
R27681 VSS.n5750 VSS.n5749 1.244
R27682 VSS.n3619 VSS.n3613 1.244
R27683 VSS.n5744 VSS.n5743 1.244
R27684 VSS.n3625 VSS.n3620 1.244
R27685 VSS.n5738 VSS.n5737 1.244
R27686 VSS.n3632 VSS.n3626 1.244
R27687 VSS.n5790 VSS.n3521 1.244
R27688 VSS.n3526 VSS.n3522 1.244
R27689 VSS.n5902 VSS.n5901 1.244
R27690 VSS.n3531 VSS.n3527 1.244
R27691 VSS.n5896 VSS.n5895 1.244
R27692 VSS.n3537 VSS.n3532 1.244
R27693 VSS.n5890 VSS.n5889 1.244
R27694 VSS.n3543 VSS.n3538 1.244
R27695 VSS.n5884 VSS.n5883 1.244
R27696 VSS.n3549 VSS.n3544 1.244
R27697 VSS.n5878 VSS.n5877 1.244
R27698 VSS.n5876 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Base 1.244
R27699 VSS.n3556 VSS.n3554 1.244
R27700 VSS.n5872 VSS.n5871 1.244
R27701 VSS.n3561 VSS.n3555 1.244
R27702 VSS.n5866 VSS.n5865 1.244
R27703 VSS.n3567 VSS.n3562 1.244
R27704 VSS.n5860 VSS.n5859 1.244
R27705 VSS.n3574 VSS.n3568 1.244
R27706 VSS.n5912 VSS.n3463 1.244
R27707 VSS.n3468 VSS.n3464 1.244
R27708 VSS.n6024 VSS.n6023 1.244
R27709 VSS.n3473 VSS.n3469 1.244
R27710 VSS.n6018 VSS.n6017 1.244
R27711 VSS.n3479 VSS.n3474 1.244
R27712 VSS.n6012 VSS.n6011 1.244
R27713 VSS.n3485 VSS.n3480 1.244
R27714 VSS.n6006 VSS.n6005 1.244
R27715 VSS.n3491 VSS.n3486 1.244
R27716 VSS.n6000 VSS.n5999 1.244
R27717 VSS.n5998 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Base 1.244
R27718 VSS.n3498 VSS.n3496 1.244
R27719 VSS.n5994 VSS.n5993 1.244
R27720 VSS.n3503 VSS.n3497 1.244
R27721 VSS.n5988 VSS.n5987 1.244
R27722 VSS.n3509 VSS.n3504 1.244
R27723 VSS.n5982 VSS.n5981 1.244
R27724 VSS.n3516 VSS.n3510 1.244
R27725 VSS.n6034 VSS.n3405 1.244
R27726 VSS.n3410 VSS.n3406 1.244
R27727 VSS.n6146 VSS.n6145 1.244
R27728 VSS.n3415 VSS.n3411 1.244
R27729 VSS.n6140 VSS.n6139 1.244
R27730 VSS.n3421 VSS.n3416 1.244
R27731 VSS.n6134 VSS.n6133 1.244
R27732 VSS.n3427 VSS.n3422 1.244
R27733 VSS.n6128 VSS.n6127 1.244
R27734 VSS.n3433 VSS.n3428 1.244
R27735 VSS.n6122 VSS.n6121 1.244
R27736 VSS.n6120 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Base 1.244
R27737 VSS.n3440 VSS.n3438 1.244
R27738 VSS.n6116 VSS.n6115 1.244
R27739 VSS.n3445 VSS.n3439 1.244
R27740 VSS.n6110 VSS.n6109 1.244
R27741 VSS.n3451 VSS.n3446 1.244
R27742 VSS.n6104 VSS.n6103 1.244
R27743 VSS.n3458 VSS.n3452 1.244
R27744 VSS.n6156 VSS.n3347 1.244
R27745 VSS.n3352 VSS.n3348 1.244
R27746 VSS.n6268 VSS.n6267 1.244
R27747 VSS.n3357 VSS.n3353 1.244
R27748 VSS.n6262 VSS.n6261 1.244
R27749 VSS.n3363 VSS.n3358 1.244
R27750 VSS.n6256 VSS.n6255 1.244
R27751 VSS.n3369 VSS.n3364 1.244
R27752 VSS.n6250 VSS.n6249 1.244
R27753 VSS.n3375 VSS.n3370 1.244
R27754 VSS.n6244 VSS.n6243 1.244
R27755 VSS.n6242 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Base 1.244
R27756 VSS.n3382 VSS.n3380 1.244
R27757 VSS.n6238 VSS.n6237 1.244
R27758 VSS.n3387 VSS.n3381 1.244
R27759 VSS.n6232 VSS.n6231 1.244
R27760 VSS.n3393 VSS.n3388 1.244
R27761 VSS.n6226 VSS.n6225 1.244
R27762 VSS.n3400 VSS.n3394 1.244
R27763 VSS.n6278 VSS.n3289 1.244
R27764 VSS.n3294 VSS.n3290 1.244
R27765 VSS.n6390 VSS.n6389 1.244
R27766 VSS.n3299 VSS.n3295 1.244
R27767 VSS.n6384 VSS.n6383 1.244
R27768 VSS.n3305 VSS.n3300 1.244
R27769 VSS.n6378 VSS.n6377 1.244
R27770 VSS.n3311 VSS.n3306 1.244
R27771 VSS.n6372 VSS.n6371 1.244
R27772 VSS.n3317 VSS.n3312 1.244
R27773 VSS.n6366 VSS.n6365 1.244
R27774 VSS.n6364 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Base 1.244
R27775 VSS.n3324 VSS.n3322 1.244
R27776 VSS.n6360 VSS.n6359 1.244
R27777 VSS.n3329 VSS.n3323 1.244
R27778 VSS.n6354 VSS.n6353 1.244
R27779 VSS.n3335 VSS.n3330 1.244
R27780 VSS.n6348 VSS.n6347 1.244
R27781 VSS.n3342 VSS.n3336 1.244
R27782 VSS.n6400 VSS.n3231 1.244
R27783 VSS.n3236 VSS.n3232 1.244
R27784 VSS.n6512 VSS.n6511 1.244
R27785 VSS.n3241 VSS.n3237 1.244
R27786 VSS.n6506 VSS.n6505 1.244
R27787 VSS.n3247 VSS.n3242 1.244
R27788 VSS.n6500 VSS.n6499 1.244
R27789 VSS.n3253 VSS.n3248 1.244
R27790 VSS.n6494 VSS.n6493 1.244
R27791 VSS.n3259 VSS.n3254 1.244
R27792 VSS.n6488 VSS.n6487 1.244
R27793 VSS.n6486 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Base 1.244
R27794 VSS.n3266 VSS.n3264 1.244
R27795 VSS.n6482 VSS.n6481 1.244
R27796 VSS.n3271 VSS.n3265 1.244
R27797 VSS.n6476 VSS.n6475 1.244
R27798 VSS.n3277 VSS.n3272 1.244
R27799 VSS.n6470 VSS.n6469 1.244
R27800 VSS.n3284 VSS.n3278 1.244
R27801 VSS.n6537 VSS.n6536 1.244
R27802 VSS.n6603 VSS.n6602 1.244
R27803 VSS.n6601 VSS.n3139 1.244
R27804 VSS.n3179 VSS.n3176 1.244
R27805 VSS.n3178 VSS.n3172 1.244
R27806 VSS.n3187 VSS.n3184 1.244
R27807 VSS.n3186 VSS.n3170 1.244
R27808 VSS.n3195 VSS.n3192 1.244
R27809 VSS.n3194 VSS.n3168 1.244
R27810 VSS.n3203 VSS.n3200 1.244
R27811 VSS.n3202 VSS.n3166 1.244
R27812 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Base VSS.n3207 1.244
R27813 VSS.n3211 VSS.n3208 1.244
R27814 VSS.n3210 VSS.n3164 1.244
R27815 VSS.n3219 VSS.n3216 1.244
R27816 VSS.n3218 VSS.n3162 1.244
R27817 VSS.n3227 VSS.n3224 1.244
R27818 VSS.n3226 VSS.n3159 1.244
R27819 VSS.n6591 VSS.n3160 1.244
R27820 VSS.n1178 VSS.n1176 1.244
R27821 VSS.n1180 VSS.n43 1.244
R27822 VSS.n1249 VSS.n1248 1.244
R27823 VSS.n1242 VSS.n44 1.244
R27824 VSS.n1241 VSS.n1239 1.244
R27825 VSS.n1236 VSS.n1184 1.244
R27826 VSS.n1188 VSS.n1187 1.244
R27827 VSS.n1230 VSS.n1229 1.244
R27828 VSS.n1192 VSS.n1190 1.244
R27829 VSS.n1224 VSS.n1223 1.244
R27830 VSS.n1196 VSS.n1194 1.244
R27831 VSS.n1220 sky130_asc_pnp_05v5_W3p40L3p40_7_0/xm1/Base 1.244
R27832 VSS.n1218 VSS.n1217 1.244
R27833 VSS.n1200 VSS.n1198 1.244
R27834 VSS.n1212 VSS.n1211 1.244
R27835 VSS.n1201 VSS.n33 1.244
R27836 VSS.n1207 VSS.n1206 1.244
R27837 VSS.n1204 VSS.n6 1.244
R27838 VSS.n1257 VSS.n4 1.244
R27839 VSS.n1262 VSS.n1261 1.244
R27840 VSS.n1088 VSS.n1086 1.244
R27841 VSS.n1090 VSS.n134 1.244
R27842 VSS.n1164 VSS.n1163 1.244
R27843 VSS.n1157 VSS.n135 1.244
R27844 VSS.n1156 VSS.n1154 1.244
R27845 VSS.n1151 VSS.n1094 1.244
R27846 VSS.n1098 VSS.n1097 1.244
R27847 VSS.n1145 VSS.n1144 1.244
R27848 VSS.n1102 VSS.n1100 1.244
R27849 VSS.n1139 VSS.n1138 1.244
R27850 VSS.n1106 VSS.n1104 1.244
R27851 VSS.n1135 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Base 1.244
R27852 VSS.n1133 VSS.n1132 1.244
R27853 VSS.n1110 VSS.n1108 1.244
R27854 VSS.n1127 VSS.n1126 1.244
R27855 VSS.n1111 VSS.n124 1.244
R27856 VSS.n1122 VSS.n1121 1.244
R27857 VSS.n1116 VSS.n1114 1.244
R27858 VSS.n1117 VSS.n96 1.244
R27859 VSS.n998 VSS.n996 1.244
R27860 VSS.n1000 VSS.n224 1.244
R27861 VSS.n1074 VSS.n1073 1.244
R27862 VSS.n1067 VSS.n225 1.244
R27863 VSS.n1066 VSS.n1064 1.244
R27864 VSS.n1061 VSS.n1004 1.244
R27865 VSS.n1008 VSS.n1007 1.244
R27866 VSS.n1055 VSS.n1054 1.244
R27867 VSS.n1012 VSS.n1010 1.244
R27868 VSS.n1049 VSS.n1048 1.244
R27869 VSS.n1016 VSS.n1014 1.244
R27870 VSS.n1045 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Base 1.244
R27871 VSS.n1043 VSS.n1042 1.244
R27872 VSS.n1020 VSS.n1018 1.244
R27873 VSS.n1037 VSS.n1036 1.244
R27874 VSS.n1021 VSS.n214 1.244
R27875 VSS.n1032 VSS.n1031 1.244
R27876 VSS.n1026 VSS.n1024 1.244
R27877 VSS.n1027 VSS.n186 1.244
R27878 VSS.n908 VSS.n906 1.244
R27879 VSS.n910 VSS.n314 1.244
R27880 VSS.n984 VSS.n983 1.244
R27881 VSS.n977 VSS.n315 1.244
R27882 VSS.n976 VSS.n974 1.244
R27883 VSS.n971 VSS.n914 1.244
R27884 VSS.n918 VSS.n917 1.244
R27885 VSS.n965 VSS.n964 1.244
R27886 VSS.n922 VSS.n920 1.244
R27887 VSS.n959 VSS.n958 1.244
R27888 VSS.n926 VSS.n924 1.244
R27889 VSS.n955 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Base 1.244
R27890 VSS.n953 VSS.n952 1.244
R27891 VSS.n930 VSS.n928 1.244
R27892 VSS.n947 VSS.n946 1.244
R27893 VSS.n931 VSS.n304 1.244
R27894 VSS.n942 VSS.n941 1.244
R27895 VSS.n936 VSS.n934 1.244
R27896 VSS.n937 VSS.n276 1.244
R27897 VSS.n818 VSS.n816 1.244
R27898 VSS.n820 VSS.n404 1.244
R27899 VSS.n894 VSS.n893 1.244
R27900 VSS.n887 VSS.n405 1.244
R27901 VSS.n886 VSS.n884 1.244
R27902 VSS.n881 VSS.n824 1.244
R27903 VSS.n828 VSS.n827 1.244
R27904 VSS.n875 VSS.n874 1.244
R27905 VSS.n832 VSS.n830 1.244
R27906 VSS.n869 VSS.n868 1.244
R27907 VSS.n836 VSS.n834 1.244
R27908 VSS.n865 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Base 1.244
R27909 VSS.n863 VSS.n862 1.244
R27910 VSS.n840 VSS.n838 1.244
R27911 VSS.n857 VSS.n856 1.244
R27912 VSS.n841 VSS.n394 1.244
R27913 VSS.n852 VSS.n851 1.244
R27914 VSS.n846 VSS.n844 1.244
R27915 VSS.n847 VSS.n366 1.244
R27916 VSS.n728 VSS.n726 1.244
R27917 VSS.n730 VSS.n494 1.244
R27918 VSS.n804 VSS.n803 1.244
R27919 VSS.n797 VSS.n495 1.244
R27920 VSS.n796 VSS.n794 1.244
R27921 VSS.n791 VSS.n734 1.244
R27922 VSS.n738 VSS.n737 1.244
R27923 VSS.n785 VSS.n784 1.244
R27924 VSS.n742 VSS.n740 1.244
R27925 VSS.n779 VSS.n778 1.244
R27926 VSS.n746 VSS.n744 1.244
R27927 VSS.n775 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Base 1.244
R27928 VSS.n773 VSS.n772 1.244
R27929 VSS.n750 VSS.n748 1.244
R27930 VSS.n767 VSS.n766 1.244
R27931 VSS.n751 VSS.n484 1.244
R27932 VSS.n762 VSS.n761 1.244
R27933 VSS.n756 VSS.n754 1.244
R27934 VSS.n757 VSS.n456 1.244
R27935 VSS.n638 VSS.n636 1.244
R27936 VSS.n640 VSS.n584 1.244
R27937 VSS.n714 VSS.n713 1.244
R27938 VSS.n707 VSS.n585 1.244
R27939 VSS.n706 VSS.n704 1.244
R27940 VSS.n701 VSS.n644 1.244
R27941 VSS.n648 VSS.n647 1.244
R27942 VSS.n695 VSS.n694 1.244
R27943 VSS.n652 VSS.n650 1.244
R27944 VSS.n689 VSS.n688 1.244
R27945 VSS.n656 VSS.n654 1.244
R27946 VSS.n685 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Base 1.244
R27947 VSS.n683 VSS.n682 1.244
R27948 VSS.n660 VSS.n658 1.244
R27949 VSS.n677 VSS.n676 1.244
R27950 VSS.n661 VSS.n574 1.244
R27951 VSS.n672 VSS.n671 1.244
R27952 VSS.n666 VSS.n664 1.244
R27953 VSS.n667 VSS.n546 1.244
R27954 VSS.n17713 VSS.n17712 1.143
R27955 VSS.n10417 VSS.n10401 1.142
R27956 VSS.n3133 VSS.n3113 1.142
R27957 VSS.n10416 VSS.n10415 1.14
R27958 VSS.n17524 sky130_asc_cap_mim_m3_1_8/VGND 1.088
R27959 VSS.n17480 sky130_asc_cap_mim_m3_1_6/VGND 1.088
R27960 VSS.n17551 VSS.n0 0.919
R27961 VSS.n15676 VSS.n15672 0.905
R27962 VSS.n15684 VSS.n15673 0.905
R27963 VSS.n15790 VSS.n15682 0.905
R27964 VSS.n15785 VSS.n15683 0.905
R27965 VSS.n15784 VSS.n15687 0.905
R27966 VSS.n15777 VSS.n15691 0.905
R27967 VSS.n15694 VSS.n15693 0.905
R27968 VSS.n15703 VSS.n15695 0.905
R27969 VSS.n15767 VSS.n15701 0.905
R27970 VSS.n15762 VSS.n15702 0.905
R27971 VSS.n15761 VSS.n15706 0.905
R27972 VSS.n15754 VSS.n15710 0.905
R27973 VSS.n15713 VSS.n15712 0.905
R27974 VSS.n15722 VSS.n15714 0.905
R27975 VSS.n15745 VSS.n15720 0.905
R27976 VSS.n15740 VSS.n15721 0.905
R27977 VSS.n15739 VSS.n15725 0.905
R27978 VSS.n15732 VSS.n15730 0.905
R27979 VSS.n15729 VSS.n13997 0.905
R27980 VSS.n14006 VSS.n13998 0.905
R27981 VSS.n16015 VSS.n14004 0.905
R27982 VSS.n16010 VSS.n14005 0.905
R27983 VSS.n16009 VSS.n14009 0.905
R27984 VSS.n16002 VSS.n14013 0.905
R27985 VSS.n15561 VSS.n14071 0.905
R27986 VSS.n15572 VSS.n15562 0.905
R27987 VSS.n15882 VSS.n15570 0.905
R27988 VSS.n15877 VSS.n15571 0.905
R27989 VSS.n15876 VSS.n15575 0.905
R27990 VSS.n15869 VSS.n15579 0.905
R27991 VSS.n15582 VSS.n15581 0.905
R27992 VSS.n15591 VSS.n15583 0.905
R27993 VSS.n15859 VSS.n15589 0.905
R27994 VSS.n15854 VSS.n15590 0.905
R27995 VSS.n15853 VSS.n15594 0.905
R27996 VSS.n15846 VSS.n15598 0.905
R27997 VSS.n15601 VSS.n15600 0.905
R27998 VSS.n15610 VSS.n15602 0.905
R27999 VSS.n15837 VSS.n15608 0.905
R28000 VSS.n15832 VSS.n15609 0.905
R28001 VSS.n15831 VSS.n15613 0.905
R28002 VSS.n15824 VSS.n15617 0.905
R28003 VSS.n15620 VSS.n15619 0.905
R28004 VSS.n15629 VSS.n15621 0.905
R28005 VSS.n15814 VSS.n15627 0.905
R28006 VSS.n15809 VSS.n15628 0.905
R28007 VSS.n15808 VSS.n15632 0.905
R28008 VSS.n15801 VSS.n15636 0.905
R28009 VSS.n15458 VSS.n14134 0.905
R28010 VSS.n15465 VSS.n14130 0.905
R28011 VSS.n15464 VSS.n14126 0.905
R28012 VSS.n14128 VSS.n14127 0.905
R28013 VSS.n15475 VSS.n14122 0.905
R28014 VSS.n15480 VSS.n14120 0.905
R28015 VSS.n15481 VSS.n14115 0.905
R28016 VSS.n15489 VSS.n15488 0.905
R28017 VSS.n15493 VSS.n14113 0.905
R28018 VSS.n15500 VSS.n14109 0.905
R28019 VSS.n15499 VSS.n14105 0.905
R28020 VSS.n14107 VSS.n14106 0.905
R28021 VSS.n15510 VSS.n14101 0.905
R28022 VSS.n15514 VSS.n14099 0.905
R28023 VSS.n15515 VSS.n14094 0.905
R28024 VSS.n15523 VSS.n15522 0.905
R28025 VSS.n15527 VSS.n14092 0.905
R28026 VSS.n15534 VSS.n14088 0.905
R28027 VSS.n15533 VSS.n14084 0.905
R28028 VSS.n14086 VSS.n14085 0.905
R28029 VSS.n15544 VSS.n14080 0.905
R28030 VSS.n15549 VSS.n14078 0.905
R28031 VSS.n15550 VSS.n14074 0.905
R28032 VSS.n15557 VSS.n14072 0.905
R28033 VSS.n15089 VSS.n15085 0.905
R28034 VSS.n15097 VSS.n15086 0.905
R28035 VSS.n15223 VSS.n15095 0.905
R28036 VSS.n15218 VSS.n15096 0.905
R28037 VSS.n15217 VSS.n15100 0.905
R28038 VSS.n15210 VSS.n15104 0.905
R28039 VSS.n15107 VSS.n15106 0.905
R28040 VSS.n15116 VSS.n15108 0.905
R28041 VSS.n15200 VSS.n15114 0.905
R28042 VSS.n15195 VSS.n15115 0.905
R28043 VSS.n15194 VSS.n15119 0.905
R28044 VSS.n15187 VSS.n15123 0.905
R28045 VSS.n15126 VSS.n15125 0.905
R28046 VSS.n15135 VSS.n15127 0.905
R28047 VSS.n15178 VSS.n15133 0.905
R28048 VSS.n15173 VSS.n15134 0.905
R28049 VSS.n15172 VSS.n15138 0.905
R28050 VSS.n15165 VSS.n15142 0.905
R28051 VSS.n15145 VSS.n15144 0.905
R28052 VSS.n15151 VSS.n15146 0.905
R28053 VSS.n15155 VSS.n15150 0.905
R28054 VSS.n15448 VSS.n14139 0.905
R28055 VSS.n15447 VSS.n14140 0.905
R28056 VSS.n15453 VSS.n15452 0.905
R28057 VSS.n14976 VSS.n14974 0.905
R28058 VSS.n14985 VSS.n14975 0.905
R28059 VSS.n15315 VSS.n14983 0.905
R28060 VSS.n15310 VSS.n14984 0.905
R28061 VSS.n15309 VSS.n14988 0.905
R28062 VSS.n15302 VSS.n14992 0.905
R28063 VSS.n14995 VSS.n14994 0.905
R28064 VSS.n15004 VSS.n14996 0.905
R28065 VSS.n15292 VSS.n15002 0.905
R28066 VSS.n15287 VSS.n15003 0.905
R28067 VSS.n15286 VSS.n15007 0.905
R28068 VSS.n15279 VSS.n15011 0.905
R28069 VSS.n15014 VSS.n15013 0.905
R28070 VSS.n15023 VSS.n15015 0.905
R28071 VSS.n15270 VSS.n15021 0.905
R28072 VSS.n15265 VSS.n15022 0.905
R28073 VSS.n15264 VSS.n15026 0.905
R28074 VSS.n15257 VSS.n15030 0.905
R28075 VSS.n15033 VSS.n15032 0.905
R28076 VSS.n15042 VSS.n15034 0.905
R28077 VSS.n15247 VSS.n15040 0.905
R28078 VSS.n15242 VSS.n15041 0.905
R28079 VSS.n15241 VSS.n15045 0.905
R28080 VSS.n15234 VSS.n15049 0.905
R28081 VSS.n14877 VSS.n14299 0.905
R28082 VSS.n14882 VSS.n14297 0.905
R28083 VSS.n14883 VSS.n14292 0.905
R28084 VSS.n14891 VSS.n14890 0.905
R28085 VSS.n14895 VSS.n14290 0.905
R28086 VSS.n14902 VSS.n14286 0.905
R28087 VSS.n14901 VSS.n14282 0.905
R28088 VSS.n14284 VSS.n14283 0.905
R28089 VSS.n14912 VSS.n14278 0.905
R28090 VSS.n14917 VSS.n14276 0.905
R28091 VSS.n14918 VSS.n14271 0.905
R28092 VSS.n14926 VSS.n14925 0.905
R28093 VSS.n14929 VSS.n14269 0.905
R28094 VSS.n14936 VSS.n14265 0.905
R28095 VSS.n14935 VSS.n14261 0.905
R28096 VSS.n14263 VSS.n14262 0.905
R28097 VSS.n14946 VSS.n14257 0.905
R28098 VSS.n14951 VSS.n14255 0.905
R28099 VSS.n14952 VSS.n14250 0.905
R28100 VSS.n14960 VSS.n14959 0.905
R28101 VSS.n14964 VSS.n14248 0.905
R28102 VSS.n14971 VSS.n14244 0.905
R28103 VSS.n14970 VSS.n14241 0.905
R28104 VSS.n15324 VSS.n14242 0.905
R28105 VSS.n14480 VSS.n14476 0.905
R28106 VSS.n14488 VSS.n14477 0.905
R28107 VSS.n14622 VSS.n14486 0.905
R28108 VSS.n14617 VSS.n14487 0.905
R28109 VSS.n14616 VSS.n14491 0.905
R28110 VSS.n14609 VSS.n14495 0.905
R28111 VSS.n14498 VSS.n14497 0.905
R28112 VSS.n14507 VSS.n14499 0.905
R28113 VSS.n14599 VSS.n14505 0.905
R28114 VSS.n14594 VSS.n14506 0.905
R28115 VSS.n14593 VSS.n14510 0.905
R28116 VSS.n14586 VSS.n14514 0.905
R28117 VSS.n14517 VSS.n14516 0.905
R28118 VSS.n14526 VSS.n14518 0.905
R28119 VSS.n14577 VSS.n14524 0.905
R28120 VSS.n14572 VSS.n14525 0.905
R28121 VSS.n14571 VSS.n14529 0.905
R28122 VSS.n14564 VSS.n14533 0.905
R28123 VSS.n14536 VSS.n14535 0.905
R28124 VSS.n14549 VSS.n14537 0.905
R28125 VSS.n14554 VSS.n14543 0.905
R28126 VSS.n14548 VSS.n14547 0.905
R28127 VSS.n14546 VSS.n14305 0.905
R28128 VSS.n14866 VSS.n14306 0.905
R28129 VSS.n14722 VSS.n14721 0.905
R28130 VSS.n14376 VSS.n14368 0.905
R28131 VSS.n14714 VSS.n14373 0.905
R28132 VSS.n14709 VSS.n14374 0.905
R28133 VSS.n14708 VSS.n14379 0.905
R28134 VSS.n14701 VSS.n14383 0.905
R28135 VSS.n14386 VSS.n14385 0.905
R28136 VSS.n14395 VSS.n14387 0.905
R28137 VSS.n14691 VSS.n14393 0.905
R28138 VSS.n14686 VSS.n14394 0.905
R28139 VSS.n14685 VSS.n14398 0.905
R28140 VSS.n14678 VSS.n14402 0.905
R28141 VSS.n14405 VSS.n14404 0.905
R28142 VSS.n14414 VSS.n14406 0.905
R28143 VSS.n14669 VSS.n14412 0.905
R28144 VSS.n14664 VSS.n14413 0.905
R28145 VSS.n14663 VSS.n14417 0.905
R28146 VSS.n14656 VSS.n14421 0.905
R28147 VSS.n14424 VSS.n14423 0.905
R28148 VSS.n14433 VSS.n14425 0.905
R28149 VSS.n14646 VSS.n14431 0.905
R28150 VSS.n14641 VSS.n14432 0.905
R28151 VSS.n14640 VSS.n14436 0.905
R28152 VSS.n14633 VSS.n14440 0.905
R28153 VSS.n11990 VSS.n11986 0.905
R28154 VSS.n11998 VSS.n11987 0.905
R28155 VSS.n12298 VSS.n11996 0.905
R28156 VSS.n12293 VSS.n11997 0.905
R28157 VSS.n12292 VSS.n12001 0.905
R28158 VSS.n12285 VSS.n12005 0.905
R28159 VSS.n12008 VSS.n12007 0.905
R28160 VSS.n12017 VSS.n12009 0.905
R28161 VSS.n12275 VSS.n12015 0.905
R28162 VSS.n12270 VSS.n12016 0.905
R28163 VSS.n12269 VSS.n12020 0.905
R28164 VSS.n12262 VSS.n12024 0.905
R28165 VSS.n12027 VSS.n12026 0.905
R28166 VSS.n12036 VSS.n12028 0.905
R28167 VSS.n12253 VSS.n12034 0.905
R28168 VSS.n12248 VSS.n12035 0.905
R28169 VSS.n12247 VSS.n12039 0.905
R28170 VSS.n12240 VSS.n12043 0.905
R28171 VSS.n12046 VSS.n12045 0.905
R28172 VSS.n12055 VSS.n12047 0.905
R28173 VSS.n12230 VSS.n12053 0.905
R28174 VSS.n12225 VSS.n12054 0.905
R28175 VSS.n12224 VSS.n12058 0.905
R28176 VSS.n12217 VSS.n12062 0.905
R28177 VSS.n11910 VSS.n11908 0.905
R28178 VSS.n11919 VSS.n11909 0.905
R28179 VSS.n12390 VSS.n11917 0.905
R28180 VSS.n12385 VSS.n11918 0.905
R28181 VSS.n12384 VSS.n11922 0.905
R28182 VSS.n12377 VSS.n11926 0.905
R28183 VSS.n11929 VSS.n11928 0.905
R28184 VSS.n11938 VSS.n11930 0.905
R28185 VSS.n12367 VSS.n11936 0.905
R28186 VSS.n12362 VSS.n11937 0.905
R28187 VSS.n12361 VSS.n11941 0.905
R28188 VSS.n12354 VSS.n11945 0.905
R28189 VSS.n11948 VSS.n11947 0.905
R28190 VSS.n11957 VSS.n11949 0.905
R28191 VSS.n12345 VSS.n11955 0.905
R28192 VSS.n12340 VSS.n11956 0.905
R28193 VSS.n12339 VSS.n11960 0.905
R28194 VSS.n12332 VSS.n11964 0.905
R28195 VSS.n11967 VSS.n11966 0.905
R28196 VSS.n11976 VSS.n11968 0.905
R28197 VSS.n12322 VSS.n11974 0.905
R28198 VSS.n12317 VSS.n11975 0.905
R28199 VSS.n12316 VSS.n11979 0.905
R28200 VSS.n12309 VSS.n11983 0.905
R28201 VSS.n11811 VSS.n11604 0.905
R28202 VSS.n11816 VSS.n11602 0.905
R28203 VSS.n11817 VSS.n11597 0.905
R28204 VSS.n11825 VSS.n11824 0.905
R28205 VSS.n11829 VSS.n11595 0.905
R28206 VSS.n11836 VSS.n11591 0.905
R28207 VSS.n11835 VSS.n11587 0.905
R28208 VSS.n11589 VSS.n11588 0.905
R28209 VSS.n11846 VSS.n11583 0.905
R28210 VSS.n11851 VSS.n11581 0.905
R28211 VSS.n11852 VSS.n11576 0.905
R28212 VSS.n11860 VSS.n11859 0.905
R28213 VSS.n11863 VSS.n11574 0.905
R28214 VSS.n11870 VSS.n11570 0.905
R28215 VSS.n11869 VSS.n11566 0.905
R28216 VSS.n11568 VSS.n11567 0.905
R28217 VSS.n11880 VSS.n11562 0.905
R28218 VSS.n11885 VSS.n11560 0.905
R28219 VSS.n11886 VSS.n11555 0.905
R28220 VSS.n11894 VSS.n11893 0.905
R28221 VSS.n11898 VSS.n11553 0.905
R28222 VSS.n11905 VSS.n11549 0.905
R28223 VSS.n11904 VSS.n11546 0.905
R28224 VSS.n12399 VSS.n11547 0.905
R28225 VSS.n11669 VSS.n11481 0.905
R28226 VSS.n11679 VSS.n11678 0.905
R28227 VSS.n11683 VSS.n11667 0.905
R28228 VSS.n11690 VSS.n11663 0.905
R28229 VSS.n11689 VSS.n11659 0.905
R28230 VSS.n11661 VSS.n11660 0.905
R28231 VSS.n11700 VSS.n11655 0.905
R28232 VSS.n11705 VSS.n11653 0.905
R28233 VSS.n11706 VSS.n11648 0.905
R28234 VSS.n11714 VSS.n11713 0.905
R28235 VSS.n11718 VSS.n11646 0.905
R28236 VSS.n11725 VSS.n11642 0.905
R28237 VSS.n11724 VSS.n11638 0.905
R28238 VSS.n11640 VSS.n11639 0.905
R28239 VSS.n11734 VSS.n11634 0.905
R28240 VSS.n11739 VSS.n11632 0.905
R28241 VSS.n11740 VSS.n11627 0.905
R28242 VSS.n11748 VSS.n11747 0.905
R28243 VSS.n11752 VSS.n11625 0.905
R28244 VSS.n11759 VSS.n11621 0.905
R28245 VSS.n11758 VSS.n11616 0.905
R28246 VSS.n11619 VSS.n11618 0.905
R28247 VSS.n11617 VSS.n11612 0.905
R28248 VSS.n11774 VSS.n11610 0.905
R28249 VSS.n13302 VSS.n12517 0.905
R28250 VSS.n13297 VSS.n13251 0.905
R28251 VSS.n13296 VSS.n13253 0.905
R28252 VSS.n13289 VSS.n13258 0.905
R28253 VSS.n13261 VSS.n13260 0.905
R28254 VSS.n13274 VSS.n13262 0.905
R28255 VSS.n13279 VSS.n13268 0.905
R28256 VSS.n13273 VSS.n13272 0.905
R28257 VSS.n13271 VSS.n11431 0.905
R28258 VSS.n11440 VSS.n11432 0.905
R28259 VSS.n13449 VSS.n11438 0.905
R28260 VSS.n13444 VSS.n11439 0.905
R28261 VSS.n13443 VSS.n11443 0.905
R28262 VSS.n13437 VSS.n11447 0.905
R28263 VSS.n11450 VSS.n11449 0.905
R28264 VSS.n11459 VSS.n11451 0.905
R28265 VSS.n13427 VSS.n11457 0.905
R28266 VSS.n13422 VSS.n11458 0.905
R28267 VSS.n13421 VSS.n11462 0.905
R28268 VSS.n13414 VSS.n11466 0.905
R28269 VSS.n11469 VSS.n11468 0.905
R28270 VSS.n11478 VSS.n11470 0.905
R28271 VSS.n13404 VSS.n11476 0.905
R28272 VSS.n13399 VSS.n11477 0.905
R28273 VSS.n13150 VSS.n12578 0.905
R28274 VSS.n13158 VSS.n13157 0.905
R28275 VSS.n13162 VSS.n12576 0.905
R28276 VSS.n13169 VSS.n12572 0.905
R28277 VSS.n13168 VSS.n12568 0.905
R28278 VSS.n12570 VSS.n12569 0.905
R28279 VSS.n13179 VSS.n12564 0.905
R28280 VSS.n13184 VSS.n12562 0.905
R28281 VSS.n13185 VSS.n12557 0.905
R28282 VSS.n13193 VSS.n13192 0.905
R28283 VSS.n13197 VSS.n12555 0.905
R28284 VSS.n13204 VSS.n12551 0.905
R28285 VSS.n13203 VSS.n12547 0.905
R28286 VSS.n12549 VSS.n12548 0.905
R28287 VSS.n13213 VSS.n12543 0.905
R28288 VSS.n13218 VSS.n12541 0.905
R28289 VSS.n13219 VSS.n12536 0.905
R28290 VSS.n13227 VSS.n13226 0.905
R28291 VSS.n13231 VSS.n12534 0.905
R28292 VSS.n13239 VSS.n12528 0.905
R28293 VSS.n13238 VSS.n12529 0.905
R28294 VSS.n13244 VSS.n13243 0.905
R28295 VSS.n13245 VSS.n12521 0.905
R28296 VSS.n13313 VSS.n12519 0.905
R28297 VSS.n13053 VSS.n12658 0.905
R28298 VSS.n13048 VSS.n12894 0.905
R28299 VSS.n13047 VSS.n12896 0.905
R28300 VSS.n13040 VSS.n12901 0.905
R28301 VSS.n12904 VSS.n12903 0.905
R28302 VSS.n12913 VSS.n12905 0.905
R28303 VSS.n13030 VSS.n12911 0.905
R28304 VSS.n13025 VSS.n12912 0.905
R28305 VSS.n13024 VSS.n12916 0.905
R28306 VSS.n13017 VSS.n12920 0.905
R28307 VSS.n12923 VSS.n12922 0.905
R28308 VSS.n12932 VSS.n12924 0.905
R28309 VSS.n13007 VSS.n12930 0.905
R28310 VSS.n13003 VSS.n12931 0.905
R28311 VSS.n13002 VSS.n12935 0.905
R28312 VSS.n12995 VSS.n12939 0.905
R28313 VSS.n12942 VSS.n12941 0.905
R28314 VSS.n12951 VSS.n12943 0.905
R28315 VSS.n12985 VSS.n12949 0.905
R28316 VSS.n12980 VSS.n12950 0.905
R28317 VSS.n12979 VSS.n12954 0.905
R28318 VSS.n12972 VSS.n12958 0.905
R28319 VSS.n12962 VSS.n12961 0.905
R28320 VSS.n12963 VSS.n12583 0.905
R28321 VSS.n12793 VSS.n12719 0.905
R28322 VSS.n12801 VSS.n12800 0.905
R28323 VSS.n12805 VSS.n12717 0.905
R28324 VSS.n12812 VSS.n12713 0.905
R28325 VSS.n12811 VSS.n12709 0.905
R28326 VSS.n12711 VSS.n12710 0.905
R28327 VSS.n12822 VSS.n12705 0.905
R28328 VSS.n12827 VSS.n12703 0.905
R28329 VSS.n12828 VSS.n12698 0.905
R28330 VSS.n12836 VSS.n12835 0.905
R28331 VSS.n12840 VSS.n12696 0.905
R28332 VSS.n12847 VSS.n12692 0.905
R28333 VSS.n12846 VSS.n12688 0.905
R28334 VSS.n12690 VSS.n12689 0.905
R28335 VSS.n12856 VSS.n12684 0.905
R28336 VSS.n12861 VSS.n12682 0.905
R28337 VSS.n12862 VSS.n12677 0.905
R28338 VSS.n12870 VSS.n12869 0.905
R28339 VSS.n12874 VSS.n12675 0.905
R28340 VSS.n12882 VSS.n12669 0.905
R28341 VSS.n12881 VSS.n12670 0.905
R28342 VSS.n12887 VSS.n12886 0.905
R28343 VSS.n12888 VSS.n12662 0.905
R28344 VSS.n13064 VSS.n12660 0.905
R28345 VSS.n7074 VSS.n7068 0.905
R28346 VSS.n7081 VSS.n7065 0.905
R28347 VSS.n7080 VSS.n7061 0.905
R28348 VSS.n7063 VSS.n7062 0.905
R28349 VSS.n7091 VSS.n7057 0.905
R28350 VSS.n7096 VSS.n7055 0.905
R28351 VSS.n7097 VSS.n7050 0.905
R28352 VSS.n7105 VSS.n7104 0.905
R28353 VSS.n7109 VSS.n7048 0.905
R28354 VSS.n7116 VSS.n7044 0.905
R28355 VSS.n7115 VSS.n7040 0.905
R28356 VSS.n7042 VSS.n7041 0.905
R28357 VSS.n7126 VSS.n7036 0.905
R28358 VSS.n7130 VSS.n7034 0.905
R28359 VSS.n7131 VSS.n7029 0.905
R28360 VSS.n7139 VSS.n7138 0.905
R28361 VSS.n7143 VSS.n7027 0.905
R28362 VSS.n7150 VSS.n7023 0.905
R28363 VSS.n7149 VSS.n7019 0.905
R28364 VSS.n7021 VSS.n7020 0.905
R28365 VSS.n7160 VSS.n7015 0.905
R28366 VSS.n7165 VSS.n7013 0.905
R28367 VSS.n7166 VSS.n7007 0.905
R28368 VSS.n7175 VSS.n7174 0.905
R28369 VSS.n8763 VSS.n8735 0.905
R28370 VSS.n8743 VSS.n8739 0.905
R28371 VSS.n8756 VSS.n8755 0.905
R28372 VSS.n8748 VSS.n8740 0.905
R28373 VSS.n8749 VSS.n6903 0.905
R28374 VSS.n6912 VSS.n6904 0.905
R28375 VSS.n8921 VSS.n6910 0.905
R28376 VSS.n8916 VSS.n6911 0.905
R28377 VSS.n8915 VSS.n6915 0.905
R28378 VSS.n8908 VSS.n6919 0.905
R28379 VSS.n6922 VSS.n6921 0.905
R28380 VSS.n6931 VSS.n6923 0.905
R28381 VSS.n8898 VSS.n6929 0.905
R28382 VSS.n8894 VSS.n6930 0.905
R28383 VSS.n8893 VSS.n6934 0.905
R28384 VSS.n8886 VSS.n6938 0.905
R28385 VSS.n6941 VSS.n6940 0.905
R28386 VSS.n6950 VSS.n6942 0.905
R28387 VSS.n8876 VSS.n6948 0.905
R28388 VSS.n8871 VSS.n6949 0.905
R28389 VSS.n8870 VSS.n6953 0.905
R28390 VSS.n8863 VSS.n6957 0.905
R28391 VSS.n6960 VSS.n6959 0.905
R28392 VSS.n7069 VSS.n6961 0.905
R28393 VSS.n8638 VSS.n7318 0.905
R28394 VSS.n8643 VSS.n7316 0.905
R28395 VSS.n8644 VSS.n7311 0.905
R28396 VSS.n8652 VSS.n8651 0.905
R28397 VSS.n8656 VSS.n7309 0.905
R28398 VSS.n8663 VSS.n7305 0.905
R28399 VSS.n8662 VSS.n7301 0.905
R28400 VSS.n7303 VSS.n7302 0.905
R28401 VSS.n8673 VSS.n7297 0.905
R28402 VSS.n8678 VSS.n7295 0.905
R28403 VSS.n8679 VSS.n7290 0.905
R28404 VSS.n8687 VSS.n8686 0.905
R28405 VSS.n8690 VSS.n7288 0.905
R28406 VSS.n8697 VSS.n7284 0.905
R28407 VSS.n8696 VSS.n7280 0.905
R28408 VSS.n7282 VSS.n7281 0.905
R28409 VSS.n8707 VSS.n7276 0.905
R28410 VSS.n8712 VSS.n7274 0.905
R28411 VSS.n8713 VSS.n7269 0.905
R28412 VSS.n8721 VSS.n8720 0.905
R28413 VSS.n8725 VSS.n7267 0.905
R28414 VSS.n8732 VSS.n7263 0.905
R28415 VSS.n8731 VSS.n7260 0.905
R28416 VSS.n8765 VSS.n7261 0.905
R28417 VSS.n8541 VSS.n8377 0.905
R28418 VSS.n8385 VSS.n8381 0.905
R28419 VSS.n8534 VSS.n8533 0.905
R28420 VSS.n8395 VSS.n8382 0.905
R28421 VSS.n8526 VSS.n8392 0.905
R28422 VSS.n8521 VSS.n8393 0.905
R28423 VSS.n8520 VSS.n8398 0.905
R28424 VSS.n8513 VSS.n8402 0.905
R28425 VSS.n8405 VSS.n8404 0.905
R28426 VSS.n8414 VSS.n8406 0.905
R28427 VSS.n8503 VSS.n8412 0.905
R28428 VSS.n8498 VSS.n8413 0.905
R28429 VSS.n8497 VSS.n8417 0.905
R28430 VSS.n8491 VSS.n8421 0.905
R28431 VSS.n8424 VSS.n8423 0.905
R28432 VSS.n8433 VSS.n8425 0.905
R28433 VSS.n8481 VSS.n8431 0.905
R28434 VSS.n8476 VSS.n8432 0.905
R28435 VSS.n8475 VSS.n8436 0.905
R28436 VSS.n8468 VSS.n8440 0.905
R28437 VSS.n8443 VSS.n8442 0.905
R28438 VSS.n8451 VSS.n8444 0.905
R28439 VSS.n8458 VSS.n8449 0.905
R28440 VSS.n8453 VSS.n8450 0.905
R28441 VSS.n8280 VSS.n7458 0.905
R28442 VSS.n8285 VSS.n7456 0.905
R28443 VSS.n8286 VSS.n7451 0.905
R28444 VSS.n8294 VSS.n8293 0.905
R28445 VSS.n8298 VSS.n7449 0.905
R28446 VSS.n8305 VSS.n7445 0.905
R28447 VSS.n8304 VSS.n7441 0.905
R28448 VSS.n7443 VSS.n7442 0.905
R28449 VSS.n8315 VSS.n7437 0.905
R28450 VSS.n8320 VSS.n7435 0.905
R28451 VSS.n8321 VSS.n7430 0.905
R28452 VSS.n8329 VSS.n8328 0.905
R28453 VSS.n8332 VSS.n7428 0.905
R28454 VSS.n8339 VSS.n7424 0.905
R28455 VSS.n8338 VSS.n7420 0.905
R28456 VSS.n7422 VSS.n7421 0.905
R28457 VSS.n8349 VSS.n7416 0.905
R28458 VSS.n8354 VSS.n7414 0.905
R28459 VSS.n8355 VSS.n7409 0.905
R28460 VSS.n8363 VSS.n8362 0.905
R28461 VSS.n8367 VSS.n7407 0.905
R28462 VSS.n8374 VSS.n7403 0.905
R28463 VSS.n8373 VSS.n7400 0.905
R28464 VSS.n8543 VSS.n7401 0.905
R28465 VSS.n8183 VSS.n8019 0.905
R28466 VSS.n8027 VSS.n8023 0.905
R28467 VSS.n8176 VSS.n8175 0.905
R28468 VSS.n8037 VSS.n8024 0.905
R28469 VSS.n8168 VSS.n8034 0.905
R28470 VSS.n8163 VSS.n8035 0.905
R28471 VSS.n8162 VSS.n8040 0.905
R28472 VSS.n8155 VSS.n8044 0.905
R28473 VSS.n8047 VSS.n8046 0.905
R28474 VSS.n8056 VSS.n8048 0.905
R28475 VSS.n8145 VSS.n8054 0.905
R28476 VSS.n8140 VSS.n8055 0.905
R28477 VSS.n8139 VSS.n8059 0.905
R28478 VSS.n8133 VSS.n8063 0.905
R28479 VSS.n8066 VSS.n8065 0.905
R28480 VSS.n8075 VSS.n8067 0.905
R28481 VSS.n8123 VSS.n8073 0.905
R28482 VSS.n8118 VSS.n8074 0.905
R28483 VSS.n8117 VSS.n8078 0.905
R28484 VSS.n8110 VSS.n8082 0.905
R28485 VSS.n8085 VSS.n8084 0.905
R28486 VSS.n8093 VSS.n8086 0.905
R28487 VSS.n8100 VSS.n8091 0.905
R28488 VSS.n8095 VSS.n8092 0.905
R28489 VSS.n7922 VSS.n7598 0.905
R28490 VSS.n7927 VSS.n7596 0.905
R28491 VSS.n7928 VSS.n7591 0.905
R28492 VSS.n7936 VSS.n7935 0.905
R28493 VSS.n7940 VSS.n7589 0.905
R28494 VSS.n7947 VSS.n7585 0.905
R28495 VSS.n7946 VSS.n7581 0.905
R28496 VSS.n7583 VSS.n7582 0.905
R28497 VSS.n7957 VSS.n7577 0.905
R28498 VSS.n7962 VSS.n7575 0.905
R28499 VSS.n7963 VSS.n7570 0.905
R28500 VSS.n7971 VSS.n7970 0.905
R28501 VSS.n7974 VSS.n7568 0.905
R28502 VSS.n7981 VSS.n7564 0.905
R28503 VSS.n7980 VSS.n7560 0.905
R28504 VSS.n7562 VSS.n7561 0.905
R28505 VSS.n7991 VSS.n7556 0.905
R28506 VSS.n7996 VSS.n7554 0.905
R28507 VSS.n7997 VSS.n7549 0.905
R28508 VSS.n8005 VSS.n8004 0.905
R28509 VSS.n8009 VSS.n7547 0.905
R28510 VSS.n8016 VSS.n7543 0.905
R28511 VSS.n8015 VSS.n7540 0.905
R28512 VSS.n8185 VSS.n7541 0.905
R28513 VSS.n7836 VSS.n7835 0.905
R28514 VSS.n7683 VSS.n7675 0.905
R28515 VSS.n7828 VSS.n7680 0.905
R28516 VSS.n7823 VSS.n7681 0.905
R28517 VSS.n7822 VSS.n7686 0.905
R28518 VSS.n7815 VSS.n7690 0.905
R28519 VSS.n7693 VSS.n7692 0.905
R28520 VSS.n7702 VSS.n7694 0.905
R28521 VSS.n7805 VSS.n7700 0.905
R28522 VSS.n7800 VSS.n7701 0.905
R28523 VSS.n7799 VSS.n7705 0.905
R28524 VSS.n7792 VSS.n7709 0.905
R28525 VSS.n7712 VSS.n7711 0.905
R28526 VSS.n7721 VSS.n7713 0.905
R28527 VSS.n7783 VSS.n7719 0.905
R28528 VSS.n7778 VSS.n7720 0.905
R28529 VSS.n7777 VSS.n7724 0.905
R28530 VSS.n7770 VSS.n7728 0.905
R28531 VSS.n7731 VSS.n7730 0.905
R28532 VSS.n7740 VSS.n7732 0.905
R28533 VSS.n7760 VSS.n7738 0.905
R28534 VSS.n7755 VSS.n7739 0.905
R28535 VSS.n7754 VSS.n7743 0.905
R28536 VSS.n7747 VSS.n7744 0.905
R28537 VSS.n6817 sky130_asc_pnp_05v5_W3p40L3p40_1_0/Collector 0.905
R28538 VSS.n5566 VSS.n3688 0.905
R28539 VSS.n5561 VSS.n5418 0.905
R28540 VSS.n5560 VSS.n5420 0.905
R28541 VSS.n5553 VSS.n5425 0.905
R28542 VSS.n5428 VSS.n5427 0.905
R28543 VSS.n5437 VSS.n5429 0.905
R28544 VSS.n5543 VSS.n5435 0.905
R28545 VSS.n5538 VSS.n5436 0.905
R28546 VSS.n5537 VSS.n5440 0.905
R28547 VSS.n5530 VSS.n5444 0.905
R28548 VSS.n5447 VSS.n5446 0.905
R28549 VSS.n5456 VSS.n5448 0.905
R28550 VSS.n5520 VSS.n5454 0.905
R28551 VSS.n5516 VSS.n5455 0.905
R28552 VSS.n5515 VSS.n5459 0.905
R28553 VSS.n5508 VSS.n5463 0.905
R28554 VSS.n5466 VSS.n5465 0.905
R28555 VSS.n5475 VSS.n5467 0.905
R28556 VSS.n5498 VSS.n5473 0.905
R28557 VSS.n5493 VSS.n5474 0.905
R28558 VSS.n5492 VSS.n5478 0.905
R28559 VSS.n5485 VSS.n5483 0.905
R28560 VSS.n5482 VSS.n3637 0.905
R28561 VSS.n3645 VSS.n3638 0.905
R28562 VSS.n5317 VSS.n3749 0.905
R28563 VSS.n5325 VSS.n5324 0.905
R28564 VSS.n5329 VSS.n3747 0.905
R28565 VSS.n5336 VSS.n3743 0.905
R28566 VSS.n5335 VSS.n3739 0.905
R28567 VSS.n3741 VSS.n3740 0.905
R28568 VSS.n5346 VSS.n3735 0.905
R28569 VSS.n5351 VSS.n3733 0.905
R28570 VSS.n5352 VSS.n3728 0.905
R28571 VSS.n5360 VSS.n5359 0.905
R28572 VSS.n5364 VSS.n3726 0.905
R28573 VSS.n5371 VSS.n3722 0.905
R28574 VSS.n5370 VSS.n3718 0.905
R28575 VSS.n3720 VSS.n3719 0.905
R28576 VSS.n5380 VSS.n3714 0.905
R28577 VSS.n5385 VSS.n3712 0.905
R28578 VSS.n5386 VSS.n3707 0.905
R28579 VSS.n5394 VSS.n5393 0.905
R28580 VSS.n5398 VSS.n3705 0.905
R28581 VSS.n5406 VSS.n3699 0.905
R28582 VSS.n5405 VSS.n3700 0.905
R28583 VSS.n5411 VSS.n5410 0.905
R28584 VSS.n5412 VSS.n3692 0.905
R28585 VSS.n5577 VSS.n3690 0.905
R28586 VSS.n5220 VSS.n3829 0.905
R28587 VSS.n5215 VSS.n5061 0.905
R28588 VSS.n5214 VSS.n5063 0.905
R28589 VSS.n5207 VSS.n5068 0.905
R28590 VSS.n5071 VSS.n5070 0.905
R28591 VSS.n5080 VSS.n5072 0.905
R28592 VSS.n5197 VSS.n5078 0.905
R28593 VSS.n5192 VSS.n5079 0.905
R28594 VSS.n5191 VSS.n5083 0.905
R28595 VSS.n5184 VSS.n5087 0.905
R28596 VSS.n5090 VSS.n5089 0.905
R28597 VSS.n5099 VSS.n5091 0.905
R28598 VSS.n5174 VSS.n5097 0.905
R28599 VSS.n5170 VSS.n5098 0.905
R28600 VSS.n5169 VSS.n5102 0.905
R28601 VSS.n5162 VSS.n5106 0.905
R28602 VSS.n5109 VSS.n5108 0.905
R28603 VSS.n5118 VSS.n5110 0.905
R28604 VSS.n5152 VSS.n5116 0.905
R28605 VSS.n5147 VSS.n5117 0.905
R28606 VSS.n5146 VSS.n5121 0.905
R28607 VSS.n5139 VSS.n5125 0.905
R28608 VSS.n5129 VSS.n5128 0.905
R28609 VSS.n5130 VSS.n3754 0.905
R28610 VSS.n4960 VSS.n3890 0.905
R28611 VSS.n4968 VSS.n4967 0.905
R28612 VSS.n4972 VSS.n3888 0.905
R28613 VSS.n4979 VSS.n3884 0.905
R28614 VSS.n4978 VSS.n3880 0.905
R28615 VSS.n3882 VSS.n3881 0.905
R28616 VSS.n4989 VSS.n3876 0.905
R28617 VSS.n4994 VSS.n3874 0.905
R28618 VSS.n4995 VSS.n3869 0.905
R28619 VSS.n5003 VSS.n5002 0.905
R28620 VSS.n5007 VSS.n3867 0.905
R28621 VSS.n5014 VSS.n3863 0.905
R28622 VSS.n5013 VSS.n3859 0.905
R28623 VSS.n3861 VSS.n3860 0.905
R28624 VSS.n5023 VSS.n3855 0.905
R28625 VSS.n5028 VSS.n3853 0.905
R28626 VSS.n5029 VSS.n3848 0.905
R28627 VSS.n5037 VSS.n5036 0.905
R28628 VSS.n5041 VSS.n3846 0.905
R28629 VSS.n5049 VSS.n3840 0.905
R28630 VSS.n5048 VSS.n3841 0.905
R28631 VSS.n5054 VSS.n5053 0.905
R28632 VSS.n5055 VSS.n3833 0.905
R28633 VSS.n5231 VSS.n3831 0.905
R28634 VSS.n4863 VSS.n3970 0.905
R28635 VSS.n4858 VSS.n4704 0.905
R28636 VSS.n4857 VSS.n4706 0.905
R28637 VSS.n4850 VSS.n4711 0.905
R28638 VSS.n4714 VSS.n4713 0.905
R28639 VSS.n4723 VSS.n4715 0.905
R28640 VSS.n4840 VSS.n4721 0.905
R28641 VSS.n4835 VSS.n4722 0.905
R28642 VSS.n4834 VSS.n4726 0.905
R28643 VSS.n4827 VSS.n4730 0.905
R28644 VSS.n4733 VSS.n4732 0.905
R28645 VSS.n4742 VSS.n4734 0.905
R28646 VSS.n4817 VSS.n4740 0.905
R28647 VSS.n4813 VSS.n4741 0.905
R28648 VSS.n4812 VSS.n4745 0.905
R28649 VSS.n4805 VSS.n4749 0.905
R28650 VSS.n4752 VSS.n4751 0.905
R28651 VSS.n4761 VSS.n4753 0.905
R28652 VSS.n4795 VSS.n4759 0.905
R28653 VSS.n4790 VSS.n4760 0.905
R28654 VSS.n4789 VSS.n4764 0.905
R28655 VSS.n4782 VSS.n4768 0.905
R28656 VSS.n4772 VSS.n4771 0.905
R28657 VSS.n4773 VSS.n3895 0.905
R28658 VSS.n4603 VSS.n4031 0.905
R28659 VSS.n4611 VSS.n4610 0.905
R28660 VSS.n4615 VSS.n4029 0.905
R28661 VSS.n4622 VSS.n4025 0.905
R28662 VSS.n4621 VSS.n4021 0.905
R28663 VSS.n4023 VSS.n4022 0.905
R28664 VSS.n4632 VSS.n4017 0.905
R28665 VSS.n4637 VSS.n4015 0.905
R28666 VSS.n4638 VSS.n4010 0.905
R28667 VSS.n4646 VSS.n4645 0.905
R28668 VSS.n4650 VSS.n4008 0.905
R28669 VSS.n4657 VSS.n4004 0.905
R28670 VSS.n4656 VSS.n4000 0.905
R28671 VSS.n4002 VSS.n4001 0.905
R28672 VSS.n4666 VSS.n3996 0.905
R28673 VSS.n4671 VSS.n3994 0.905
R28674 VSS.n4672 VSS.n3989 0.905
R28675 VSS.n4680 VSS.n4679 0.905
R28676 VSS.n4684 VSS.n3987 0.905
R28677 VSS.n4692 VSS.n3981 0.905
R28678 VSS.n4691 VSS.n3982 0.905
R28679 VSS.n4697 VSS.n4696 0.905
R28680 VSS.n4698 VSS.n3974 0.905
R28681 VSS.n4874 VSS.n3972 0.905
R28682 VSS.n4506 VSS.n4111 0.905
R28683 VSS.n4501 VSS.n4347 0.905
R28684 VSS.n4500 VSS.n4349 0.905
R28685 VSS.n4493 VSS.n4354 0.905
R28686 VSS.n4357 VSS.n4356 0.905
R28687 VSS.n4366 VSS.n4358 0.905
R28688 VSS.n4483 VSS.n4364 0.905
R28689 VSS.n4478 VSS.n4365 0.905
R28690 VSS.n4477 VSS.n4369 0.905
R28691 VSS.n4470 VSS.n4373 0.905
R28692 VSS.n4376 VSS.n4375 0.905
R28693 VSS.n4385 VSS.n4377 0.905
R28694 VSS.n4460 VSS.n4383 0.905
R28695 VSS.n4456 VSS.n4384 0.905
R28696 VSS.n4455 VSS.n4388 0.905
R28697 VSS.n4448 VSS.n4392 0.905
R28698 VSS.n4395 VSS.n4394 0.905
R28699 VSS.n4404 VSS.n4396 0.905
R28700 VSS.n4438 VSS.n4402 0.905
R28701 VSS.n4433 VSS.n4403 0.905
R28702 VSS.n4432 VSS.n4407 0.905
R28703 VSS.n4425 VSS.n4411 0.905
R28704 VSS.n4415 VSS.n4414 0.905
R28705 VSS.n4416 VSS.n4036 0.905
R28706 VSS.n4246 VSS.n4172 0.905
R28707 VSS.n4254 VSS.n4253 0.905
R28708 VSS.n4258 VSS.n4170 0.905
R28709 VSS.n4265 VSS.n4166 0.905
R28710 VSS.n4264 VSS.n4162 0.905
R28711 VSS.n4164 VSS.n4163 0.905
R28712 VSS.n4275 VSS.n4158 0.905
R28713 VSS.n4280 VSS.n4156 0.905
R28714 VSS.n4281 VSS.n4151 0.905
R28715 VSS.n4289 VSS.n4288 0.905
R28716 VSS.n4293 VSS.n4149 0.905
R28717 VSS.n4300 VSS.n4145 0.905
R28718 VSS.n4299 VSS.n4141 0.905
R28719 VSS.n4143 VSS.n4142 0.905
R28720 VSS.n4309 VSS.n4137 0.905
R28721 VSS.n4314 VSS.n4135 0.905
R28722 VSS.n4315 VSS.n4130 0.905
R28723 VSS.n4323 VSS.n4322 0.905
R28724 VSS.n4327 VSS.n4128 0.905
R28725 VSS.n4335 VSS.n4122 0.905
R28726 VSS.n4334 VSS.n4123 0.905
R28727 VSS.n4340 VSS.n4339 0.905
R28728 VSS.n4341 VSS.n4115 0.905
R28729 VSS.n4517 VSS.n4113 0.905
R28730 VSS.n2802 VSS.n1312 0.905
R28731 VSS.n2813 VSS.n2803 0.905
R28732 VSS.n2956 VSS.n2811 0.905
R28733 VSS.n2951 VSS.n2812 0.905
R28734 VSS.n2950 VSS.n2816 0.905
R28735 VSS.n2943 VSS.n2820 0.905
R28736 VSS.n2823 VSS.n2822 0.905
R28737 VSS.n2832 VSS.n2824 0.905
R28738 VSS.n2933 VSS.n2830 0.905
R28739 VSS.n2928 VSS.n2831 0.905
R28740 VSS.n2927 VSS.n2835 0.905
R28741 VSS.n2920 VSS.n2839 0.905
R28742 VSS.n2842 VSS.n2841 0.905
R28743 VSS.n2851 VSS.n2843 0.905
R28744 VSS.n2911 VSS.n2849 0.905
R28745 VSS.n2906 VSS.n2850 0.905
R28746 VSS.n2905 VSS.n2854 0.905
R28747 VSS.n2898 VSS.n2858 0.905
R28748 VSS.n2861 VSS.n2860 0.905
R28749 VSS.n2870 VSS.n2862 0.905
R28750 VSS.n2888 VSS.n2868 0.905
R28751 VSS.n2883 VSS.n2869 0.905
R28752 VSS.n2882 VSS.n2877 0.905
R28753 VSS.n2875 VSS.n1269 0.905
R28754 VSS.n2699 VSS.n1375 0.905
R28755 VSS.n2706 VSS.n1371 0.905
R28756 VSS.n2705 VSS.n1367 0.905
R28757 VSS.n1369 VSS.n1368 0.905
R28758 VSS.n2716 VSS.n1363 0.905
R28759 VSS.n2721 VSS.n1361 0.905
R28760 VSS.n2722 VSS.n1356 0.905
R28761 VSS.n2730 VSS.n2729 0.905
R28762 VSS.n2734 VSS.n1354 0.905
R28763 VSS.n2741 VSS.n1350 0.905
R28764 VSS.n2740 VSS.n1346 0.905
R28765 VSS.n1348 VSS.n1347 0.905
R28766 VSS.n2751 VSS.n1342 0.905
R28767 VSS.n2755 VSS.n1340 0.905
R28768 VSS.n2756 VSS.n1335 0.905
R28769 VSS.n2764 VSS.n2763 0.905
R28770 VSS.n2768 VSS.n1333 0.905
R28771 VSS.n2775 VSS.n1329 0.905
R28772 VSS.n2774 VSS.n1325 0.905
R28773 VSS.n1327 VSS.n1326 0.905
R28774 VSS.n2785 VSS.n1321 0.905
R28775 VSS.n2790 VSS.n1319 0.905
R28776 VSS.n2791 VSS.n1315 0.905
R28777 VSS.n2798 VSS.n1313 0.905
R28778 VSS.n2330 VSS.n2326 0.905
R28779 VSS.n2338 VSS.n2327 0.905
R28780 VSS.n2464 VSS.n2336 0.905
R28781 VSS.n2459 VSS.n2337 0.905
R28782 VSS.n2458 VSS.n2341 0.905
R28783 VSS.n2451 VSS.n2345 0.905
R28784 VSS.n2348 VSS.n2347 0.905
R28785 VSS.n2357 VSS.n2349 0.905
R28786 VSS.n2441 VSS.n2355 0.905
R28787 VSS.n2436 VSS.n2356 0.905
R28788 VSS.n2435 VSS.n2360 0.905
R28789 VSS.n2428 VSS.n2364 0.905
R28790 VSS.n2367 VSS.n2366 0.905
R28791 VSS.n2376 VSS.n2368 0.905
R28792 VSS.n2419 VSS.n2374 0.905
R28793 VSS.n2414 VSS.n2375 0.905
R28794 VSS.n2413 VSS.n2379 0.905
R28795 VSS.n2406 VSS.n2383 0.905
R28796 VSS.n2386 VSS.n2385 0.905
R28797 VSS.n2392 VSS.n2387 0.905
R28798 VSS.n2396 VSS.n2391 0.905
R28799 VSS.n2689 VSS.n1380 0.905
R28800 VSS.n2688 VSS.n1381 0.905
R28801 VSS.n2694 VSS.n2693 0.905
R28802 VSS.n2217 VSS.n2215 0.905
R28803 VSS.n2226 VSS.n2216 0.905
R28804 VSS.n2556 VSS.n2224 0.905
R28805 VSS.n2551 VSS.n2225 0.905
R28806 VSS.n2550 VSS.n2229 0.905
R28807 VSS.n2543 VSS.n2233 0.905
R28808 VSS.n2236 VSS.n2235 0.905
R28809 VSS.n2245 VSS.n2237 0.905
R28810 VSS.n2533 VSS.n2243 0.905
R28811 VSS.n2528 VSS.n2244 0.905
R28812 VSS.n2527 VSS.n2248 0.905
R28813 VSS.n2520 VSS.n2252 0.905
R28814 VSS.n2255 VSS.n2254 0.905
R28815 VSS.n2264 VSS.n2256 0.905
R28816 VSS.n2511 VSS.n2262 0.905
R28817 VSS.n2506 VSS.n2263 0.905
R28818 VSS.n2505 VSS.n2267 0.905
R28819 VSS.n2498 VSS.n2271 0.905
R28820 VSS.n2274 VSS.n2273 0.905
R28821 VSS.n2283 VSS.n2275 0.905
R28822 VSS.n2488 VSS.n2281 0.905
R28823 VSS.n2483 VSS.n2282 0.905
R28824 VSS.n2482 VSS.n2286 0.905
R28825 VSS.n2475 VSS.n2290 0.905
R28826 VSS.n2118 VSS.n1540 0.905
R28827 VSS.n2123 VSS.n1538 0.905
R28828 VSS.n2124 VSS.n1533 0.905
R28829 VSS.n2132 VSS.n2131 0.905
R28830 VSS.n2136 VSS.n1531 0.905
R28831 VSS.n2143 VSS.n1527 0.905
R28832 VSS.n2142 VSS.n1523 0.905
R28833 VSS.n1525 VSS.n1524 0.905
R28834 VSS.n2153 VSS.n1519 0.905
R28835 VSS.n2158 VSS.n1517 0.905
R28836 VSS.n2159 VSS.n1512 0.905
R28837 VSS.n2167 VSS.n2166 0.905
R28838 VSS.n2170 VSS.n1510 0.905
R28839 VSS.n2177 VSS.n1506 0.905
R28840 VSS.n2176 VSS.n1502 0.905
R28841 VSS.n1504 VSS.n1503 0.905
R28842 VSS.n2187 VSS.n1498 0.905
R28843 VSS.n2192 VSS.n1496 0.905
R28844 VSS.n2193 VSS.n1491 0.905
R28845 VSS.n2201 VSS.n2200 0.905
R28846 VSS.n2205 VSS.n1489 0.905
R28847 VSS.n2212 VSS.n1485 0.905
R28848 VSS.n2211 VSS.n1482 0.905
R28849 VSS.n2565 VSS.n1483 0.905
R28850 VSS.n1721 VSS.n1717 0.905
R28851 VSS.n1729 VSS.n1718 0.905
R28852 VSS.n1863 VSS.n1727 0.905
R28853 VSS.n1858 VSS.n1728 0.905
R28854 VSS.n1857 VSS.n1732 0.905
R28855 VSS.n1850 VSS.n1736 0.905
R28856 VSS.n1739 VSS.n1738 0.905
R28857 VSS.n1748 VSS.n1740 0.905
R28858 VSS.n1840 VSS.n1746 0.905
R28859 VSS.n1835 VSS.n1747 0.905
R28860 VSS.n1834 VSS.n1751 0.905
R28861 VSS.n1827 VSS.n1755 0.905
R28862 VSS.n1758 VSS.n1757 0.905
R28863 VSS.n1767 VSS.n1759 0.905
R28864 VSS.n1818 VSS.n1765 0.905
R28865 VSS.n1813 VSS.n1766 0.905
R28866 VSS.n1812 VSS.n1770 0.905
R28867 VSS.n1805 VSS.n1774 0.905
R28868 VSS.n1777 VSS.n1776 0.905
R28869 VSS.n1790 VSS.n1778 0.905
R28870 VSS.n1795 VSS.n1784 0.905
R28871 VSS.n1789 VSS.n1788 0.905
R28872 VSS.n1787 VSS.n1546 0.905
R28873 VSS.n2107 VSS.n1547 0.905
R28874 VSS.n1963 VSS.n1962 0.905
R28875 VSS.n1617 VSS.n1609 0.905
R28876 VSS.n1955 VSS.n1614 0.905
R28877 VSS.n1950 VSS.n1615 0.905
R28878 VSS.n1949 VSS.n1620 0.905
R28879 VSS.n1942 VSS.n1624 0.905
R28880 VSS.n1627 VSS.n1626 0.905
R28881 VSS.n1636 VSS.n1628 0.905
R28882 VSS.n1932 VSS.n1634 0.905
R28883 VSS.n1927 VSS.n1635 0.905
R28884 VSS.n1926 VSS.n1639 0.905
R28885 VSS.n1919 VSS.n1643 0.905
R28886 VSS.n1646 VSS.n1645 0.905
R28887 VSS.n1655 VSS.n1647 0.905
R28888 VSS.n1910 VSS.n1653 0.905
R28889 VSS.n1905 VSS.n1654 0.905
R28890 VSS.n1904 VSS.n1658 0.905
R28891 VSS.n1897 VSS.n1662 0.905
R28892 VSS.n1665 VSS.n1664 0.905
R28893 VSS.n1674 VSS.n1666 0.905
R28894 VSS.n1887 VSS.n1672 0.905
R28895 VSS.n1882 VSS.n1673 0.905
R28896 VSS.n1881 VSS.n1677 0.905
R28897 VSS.n1874 VSS.n1681 0.905
R28898 VSS.n3127 VSS.n3124 0.861
R28899 VSS.n3129 VSS.n3128 0.861
R28900 VSS.n3134 VSS.n3133 0.855
R28901 VSS.n16771 VSS.n16770 0.785
R28902 VSS.n16861 VSS.n16860 0.785
R28903 VSS.n16951 VSS.n16950 0.785
R28904 VSS.n17041 VSS.n17040 0.785
R28905 VSS.n17131 VSS.n17130 0.785
R28906 VSS.n17221 VSS.n17220 0.785
R28907 VSS.n17311 VSS.n17310 0.785
R28908 VSS.n11238 VSS.n11237 0.785
R28909 VSS.n11328 VSS.n11327 0.785
R28910 VSS.n11418 VSS.n11417 0.785
R28911 VSS.n13538 VSS.n13537 0.785
R28912 VSS.n13628 VSS.n13627 0.785
R28913 VSS.n13718 VSS.n13717 0.785
R28914 VSS.n13808 VSS.n13807 0.785
R28915 VSS.n9816 VSS.n9815 0.785
R28916 VSS.n9906 VSS.n9905 0.785
R28917 VSS.n9996 VSS.n9995 0.785
R28918 VSS.n10086 VSS.n10085 0.785
R28919 VSS.n10176 VSS.n10175 0.785
R28920 VSS.n10318 VSS.n10265 0.785
R28921 VSS.n9161 VSS.n9160 0.785
R28922 VSS.n6519 VSS.n6518 0.785
R28923 VSS.n6397 VSS.n6396 0.785
R28924 VSS.n6275 VSS.n6274 0.785
R28925 VSS.n6153 VSS.n6152 0.785
R28926 VSS.n6031 VSS.n6030 0.785
R28927 VSS.n5909 VSS.n5908 0.785
R28928 VSS.n5787 VSS.n5786 0.785
R28929 VSS.n724 VSS.n723 0.785
R28930 VSS.n814 VSS.n813 0.785
R28931 VSS.n904 VSS.n903 0.785
R28932 VSS.n994 VSS.n993 0.785
R28933 VSS.n1084 VSS.n1083 0.785
R28934 VSS.n1174 VSS.n1173 0.785
R28935 VSS.n3048 VSS.n3047 0.784
R28936 VSS.n10443 VSS.n10428 0.752
R28937 VSS.n10468 VSS.n10467 0.752
R28938 VSS.n17678 VSS.n17677 0.752
R28939 VSS.n17684 VSS.n17648 0.752
R28940 VSS.n17304 VSS.n16055 0.735
R28941 VSS.n17214 VSS.n16145 0.735
R28942 VSS.n17124 VSS.n16235 0.735
R28943 VSS.n17034 VSS.n16325 0.735
R28944 VSS.n16944 VSS.n16415 0.735
R28945 VSS.n16854 VSS.n16505 0.735
R28946 VSS.n16764 VSS.n16595 0.735
R28947 VSS.n10259 VSS.n9190 0.735
R28948 VSS.n10169 VSS.n9280 0.735
R28949 VSS.n10079 VSS.n9370 0.735
R28950 VSS.n9989 VSS.n9460 0.735
R28951 VSS.n9899 VSS.n9550 0.735
R28952 VSS.n9809 VSS.n9640 0.735
R28953 VSS.n10326 VSS.n8977 0.735
R28954 VSS.n5735 VSS.n3630 0.735
R28955 VSS.n5857 VSS.n3572 0.735
R28956 VSS.n5979 VSS.n3514 0.735
R28957 VSS.n6101 VSS.n3456 0.735
R28958 VSS.n6223 VSS.n3398 0.735
R28959 VSS.n6345 VSS.n3340 0.735
R28960 VSS.n6467 VSS.n3282 0.735
R28961 VSS.n6597 VSS.n6596 0.735
R28962 VSS.n1255 VSS.n7 0.735
R28963 VSS.n1167 VSS.n98 0.735
R28964 VSS.n1077 VSS.n188 0.735
R28965 VSS.n987 VSS.n278 0.735
R28966 VSS.n897 VSS.n368 0.735
R28967 VSS.n807 VSS.n458 0.735
R28968 VSS.n717 VSS.n548 0.735
R28969 VSS.n3048 VSS.n1265 0.535
R28970 sky130_asc_pnp_05v5_W3p40L3p40_8_3/xm1/Base VSS.n17432 0.533
R28971 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Base VSS.n17270 0.533
R28972 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Base VSS.n17180 0.533
R28973 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Base VSS.n17090 0.533
R28974 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Base VSS.n17000 0.533
R28975 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Base VSS.n16910 0.533
R28976 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Base VSS.n16820 0.533
R28977 sky130_asc_pnp_05v5_W3p40L3p40_8_3/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Base VSS.n16730 0.533
R28978 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Base VSS.n11198 0.533
R28979 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Base VSS.n11288 0.533
R28980 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Base VSS.n11378 0.533
R28981 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Base VSS.n13497 0.533
R28982 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Base VSS.n13588 0.533
R28983 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Base VSS.n13678 0.533
R28984 sky130_asc_pnp_05v5_W3p40L3p40_8_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Base VSS.n13768 0.533
R28985 sky130_asc_pnp_05v5_W3p40L3p40_8_0/xm1/Base VSS.n13924 0.533
R28986 VSS.n9076 sky130_asc_pnp_05v5_W3p40L3p40_8_1/xm1/Base 0.533
R28987 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Base VSS.n10225 0.533
R28988 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Base VSS.n10135 0.533
R28989 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Base VSS.n10045 0.533
R28990 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Base VSS.n9955 0.533
R28991 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Base VSS.n9865 0.533
R28992 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Base VSS.n9775 0.533
R28993 VSS.n8961 sky130_asc_pnp_05v5_W3p40L3p40_8_1/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Base 0.533
R28994 VSS.n3614 sky130_asc_pnp_05v5_W3p40L3p40_8_2/xm1/Base 0.533
R28995 VSS.n3556 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Base 0.533
R28996 VSS.n3498 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Base 0.533
R28997 VSS.n3440 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Base 0.533
R28998 VSS.n3382 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Base 0.533
R28999 VSS.n3324 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Base 0.533
R29000 VSS.n3266 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Base 0.533
R29001 VSS.n3208 sky130_asc_pnp_05v5_W3p40L3p40_8_2/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_6/Base 0.533
R29002 sky130_asc_pnp_05v5_W3p40L3p40_7_0/xm1/Base VSS.n1218 0.533
R29003 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0/Base VSS.n1133 0.533
R29004 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1/Base VSS.n1043 0.533
R29005 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2/Base VSS.n953 0.533
R29006 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3/Base VSS.n863 0.533
R29007 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4/Base VSS.n773 0.533
R29008 sky130_asc_pnp_05v5_W3p40L3p40_7_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_5/Base VSS.n683 0.533
R29009 VSS.n17712 VSS.n17711 0.485
R29010 VSS.n17712 VSS.n17637 0.485
R29011 VSS.n17712 VSS.n17633 0.485
R29012 VSS.n17712 VSS.n17618 0.481
R29013 VSS.n17712 VSS.n17623 0.481
R29014 VSS.n17712 VSS.n17625 0.481
R29015 VSS.n17609 VSS.n17607 0.438
R29016 VSS.n17704 sky130_asc_nfet_01v8_lvt_1_0/VGND 0.426
R29017 sky130_asc_cap_mim_m3_1_4/VGND VSS.n17704 0.422
R29018 VSS.n10456 VSS.n10431 0.414
R29019 VSS.n10482 VSS.n10420 0.414
R29020 VSS.n17662 VSS.n17655 0.414
R29021 VSS.n17695 VSS.n17643 0.413
R29022 VSS.n17525 sky130_asc_res_xhigh_po_2p85_2_0/VGND 0.403
R29023 VSS.n10452 VSS.n10430 0.382
R29024 VSS.n10477 VSS.n10422 0.382
R29025 VSS.n17667 VSS.n17653 0.382
R29026 VSS.n17693 VSS.n17692 0.382
R29027 VSS.n6896 VSS.n6882 0.372
R29028 VSS.n16024 VSS.n16023 0.357
R29029 VSS.n13513 VSS.n13457 0.357
R29030 VSS.n10371 VSS.n8929 0.357
R29031 VSS.n5664 VSS.n5663 0.357
R29032 VSS.n1263 VSS.n1262 0.355
R29033 VSS.n10447 VSS.n10429 0.35
R29034 VSS.n10472 VSS.n10424 0.35
R29035 VSS.n17673 VSS.n17672 0.35
R29036 VSS.n17687 VSS.n17686 0.349
R29037 VSS.n6607 sky130_asc_res_xhigh_po_2p85_1_0/VGND 0.333
R29038 VSS.n6607 sky130_asc_res_xhigh_po_2p85_1_0/Rout 0.331
R29039 VSS.n17525 sky130_asc_res_xhigh_po_2p85_2_0/Rout 0.331
R29040 VSS.n17550 sky130_asc_res_xhigh_po_2p85_2_1/Rout 0.33
R29041 VSS.n10463 VSS.n10428 0.317
R29042 VSS.n17650 VSS.n17648 0.317
R29043 VSS.n14631 VSS.n14630 0.296
R29044 VSS.n14867 VSS.n14298 0.296
R29045 VSS.n15325 VSS.n15323 0.296
R29046 VSS.n15232 VSS.n15231 0.296
R29047 VSS.n15455 VSS.n14135 0.296
R29048 VSS.n15890 VSS.n15559 0.296
R29049 VSS.n15799 VSS.n15798 0.296
R29050 VSS.n13063 VSS.n12659 0.296
R29051 VSS.n12959 VSS.n12584 0.296
R29052 VSS.n13312 VSS.n12518 0.296
R29053 VSS.n13400 VSS.n11480 0.296
R29054 VSS.n11773 VSS.n11603 0.296
R29055 VSS.n12400 VSS.n12398 0.296
R29056 VSS.n12307 VSS.n12306 0.296
R29057 VSS.n7745 VSS.n7597 0.296
R29058 VSS.n8186 VSS.n8018 0.296
R29059 VSS.n8096 VSS.n7457 0.296
R29060 VSS.n8544 VSS.n8376 0.296
R29061 VSS.n8454 VSS.n7317 0.296
R29062 VSS.n8766 VSS.n8734 0.296
R29063 VSS.n7071 VSS.n7070 0.296
R29064 VSS.n4516 VSS.n4112 0.296
R29065 VSS.n4412 VSS.n4037 0.296
R29066 VSS.n4873 VSS.n3971 0.296
R29067 VSS.n4769 VSS.n3896 0.296
R29068 VSS.n5230 VSS.n3830 0.296
R29069 VSS.n5126 VSS.n3755 0.296
R29070 VSS.n5576 VSS.n3689 0.296
R29071 VSS.n1872 VSS.n1871 0.296
R29072 VSS.n2108 VSS.n1539 0.296
R29073 VSS.n2566 VSS.n2564 0.296
R29074 VSS.n2473 VSS.n2472 0.296
R29075 VSS.n2696 VSS.n1376 0.296
R29076 VSS.n2964 VSS.n2800 0.296
R29077 VSS.n14630 VSS.n14629 0.29
R29078 VSS.n14879 VSS.n14298 0.29
R29079 VSS.n15323 VSS.n15322 0.29
R29080 VSS.n15231 VSS.n15230 0.29
R29081 VSS.n15456 VSS.n15455 0.29
R29082 VSS.n15890 VSS.n15889 0.29
R29083 VSS.n15798 VSS.n15797 0.29
R29084 VSS.n13051 VSS.n12659 0.29
R29085 VSS.n12584 VSS.n12579 0.29
R29086 VSS.n13300 VSS.n12518 0.29
R29087 VSS.n11670 VSS.n11480 0.29
R29088 VSS.n11813 VSS.n11603 0.29
R29089 VSS.n12398 VSS.n12397 0.29
R29090 VSS.n12306 VSS.n12305 0.29
R29091 VSS.n7924 VSS.n7597 0.29
R29092 VSS.n8025 VSS.n8018 0.29
R29093 VSS.n8282 VSS.n7457 0.29
R29094 VSS.n8383 VSS.n8376 0.29
R29095 VSS.n8640 VSS.n7317 0.29
R29096 VSS.n8741 VSS.n8734 0.29
R29097 VSS.n7072 VSS.n7071 0.29
R29098 VSS.n4504 VSS.n4112 0.29
R29099 VSS.n4037 VSS.n4032 0.29
R29100 VSS.n4861 VSS.n3971 0.29
R29101 VSS.n3896 VSS.n3891 0.29
R29102 VSS.n5218 VSS.n3830 0.29
R29103 VSS.n3755 VSS.n3750 0.29
R29104 VSS.n5564 VSS.n3689 0.29
R29105 VSS.n1871 VSS.n1870 0.29
R29106 VSS.n2120 VSS.n1539 0.29
R29107 VSS.n2564 VSS.n2563 0.29
R29108 VSS.n2472 VSS.n2471 0.29
R29109 VSS.n2697 VSS.n2696 0.29
R29110 VSS.n2964 VSS.n2963 0.29
R29111 VSS.n15998 VSS.n14014 0.258
R29112 VSS.n12213 VSS.n12063 0.258
R29113 VSS.n7178 VSS.n7005 0.258
R29114 VSS.n3648 VSS.n3644 0.258
R29115 VSS.n3045 VSS.n3044 0.258
R29116 VSS.n17513 VSS.t154 0.219
R29117 VSS.n17469 VSS.t156 0.219
R29118 VSS.n10403 VSS.t160 0.219
R29119 VSS.n6884 VSS.t106 0.219
R29120 VSS.n3115 VSS.t178 0.219
R29121 VSS.n13965 VSS.n10400 0.219
R29122 VSS.n17485 VSS.n17484 0.219
R29123 VSS.n17481 sky130_asc_pnp_05v5_W3p40L3p40_8_3/VGND 0.208
R29124 VSS.n10489 sky130_asc_pnp_05v5_W3p40L3p40_8_0/VGND 0.208
R29125 VSS.n6882 sky130_asc_cap_mim_m3_1_5/VGND 0.208
R29126 sky130_asc_pnp_05v5_W3p40L3p40_7_0/VGND VSS.n17600 0.207
R29127 VSS.n13962 VSS.n10489 0.198
R29128 VSS.n17522 VSS.n17521 0.196
R29129 VSS.n17514 VSS.n17513 0.196
R29130 VSS.n17515 VSS.n17514 0.196
R29131 VSS.n17516 VSS.n17515 0.196
R29132 VSS.n17517 VSS.n17516 0.196
R29133 VSS.n17518 VSS.n17517 0.196
R29134 VSS.n17519 VSS.n17518 0.196
R29135 VSS.n17478 VSS.n17477 0.196
R29136 VSS.n17470 VSS.n17469 0.196
R29137 VSS.n17471 VSS.n17470 0.196
R29138 VSS.n17472 VSS.n17471 0.196
R29139 VSS.n17473 VSS.n17472 0.196
R29140 VSS.n17474 VSS.n17473 0.196
R29141 VSS.n17475 VSS.n17474 0.196
R29142 VSS.n10412 VSS.n10411 0.196
R29143 VSS.n10404 VSS.n10403 0.196
R29144 VSS.n10405 VSS.n10404 0.196
R29145 VSS.n10406 VSS.n10405 0.196
R29146 VSS.n10407 VSS.n10406 0.196
R29147 VSS.n10408 VSS.n10407 0.196
R29148 VSS.n10409 VSS.n10408 0.196
R29149 VSS.n6885 VSS.n6884 0.196
R29150 VSS.n6886 VSS.n6885 0.196
R29151 VSS.n6887 VSS.n6886 0.196
R29152 VSS.n6888 VSS.n6887 0.196
R29153 VSS.n6889 VSS.n6888 0.196
R29154 VSS.n6890 VSS.n6889 0.196
R29155 VSS.n6891 VSS.n6890 0.196
R29156 VSS.n3116 VSS.n3115 0.196
R29157 VSS.n3117 VSS.n3116 0.196
R29158 VSS.n3118 VSS.n3117 0.196
R29159 VSS.n3119 VSS.n3118 0.196
R29160 VSS.n3120 VSS.n3119 0.196
R29161 VSS.n3121 VSS.n3120 0.196
R29162 VSS.n3122 VSS.n3121 0.196
R29163 VSS.n3123 VSS.n3122 0.196
R29164 VSS.n10465 VSS.n10427 0.19
R29165 VSS.n10466 VSS.n10465 0.19
R29166 VSS.n17681 VSS.n17649 0.19
R29167 VSS.n17682 VSS.n17681 0.19
R29168 VSS.n17482 VSS.n17481 0.184
R29169 VSS.n17523 VSS.n17519 0.173
R29170 VSS.n17479 VSS.n17475 0.173
R29171 VSS.n1266 sky130_asc_pnp_05v5_W3p40L3p40_7_0/Collector 0.167
R29172 VSS.n10486 VSS.n10485 0.163
R29173 VSS.n16000 VSS.n15999 0.148
R29174 VSS.n16770 VSS.n16592 0.148
R29175 VSS.n16860 VSS.n16502 0.148
R29176 VSS.n16950 VSS.n16412 0.148
R29177 VSS.n17040 VSS.n16322 0.148
R29178 VSS.n17130 VSS.n16232 0.148
R29179 VSS.n17220 VSS.n16142 0.148
R29180 VSS.n17310 VSS.n16052 0.148
R29181 VSS.n17333 VSS.n17332 0.148
R29182 VSS.n12215 VSS.n12214 0.148
R29183 VSS.n11237 VSS.n11059 0.148
R29184 VSS.n11327 VSS.n10969 0.148
R29185 VSS.n11417 VSS.n10879 0.148
R29186 VSS.n13537 VSS.n10789 0.148
R29187 VSS.n13627 VSS.n10699 0.148
R29188 VSS.n13717 VSS.n10609 0.148
R29189 VSS.n13807 VSS.n10519 0.148
R29190 VSS.n13833 VSS.n13832 0.148
R29191 VSS.n7177 VSS.n7176 0.148
R29192 VSS.n9815 VSS.n9637 0.148
R29193 VSS.n9905 VSS.n9547 0.148
R29194 VSS.n9995 VSS.n9457 0.148
R29195 VSS.n10085 VSS.n9367 0.148
R29196 VSS.n10175 VSS.n9277 0.148
R29197 VSS.n10265 VSS.n9187 0.148
R29198 VSS.n9161 VSS.n8980 0.148
R29199 VSS.n9150 VSS.n9097 0.148
R29200 VSS.n3647 VSS.n3646 0.148
R29201 VSS.n6592 VSS.n6519 0.148
R29202 VSS.n6397 VSS.n3286 0.148
R29203 VSS.n6275 VSS.n3344 0.148
R29204 VSS.n6153 VSS.n3402 0.148
R29205 VSS.n6031 VSS.n3460 0.148
R29206 VSS.n5909 VSS.n3518 0.148
R29207 VSS.n5787 VSS.n3576 0.148
R29208 VSS.n5665 VSS.n3634 0.148
R29209 VSS.n723 VSS.n545 0.148
R29210 VSS.n813 VSS.n455 0.148
R29211 VSS.n903 VSS.n365 0.148
R29212 VSS.n993 VSS.n275 0.148
R29213 VSS.n1083 VSS.n185 0.148
R29214 VSS.n1173 VSS.n95 0.148
R29215 VSS.n10457 VSS.n10455 0.144
R29216 VSS.n10451 VSS.n10450 0.144
R29217 VSS.n10446 VSS.n10445 0.144
R29218 VSS.n10471 VSS.n10470 0.144
R29219 VSS.n10476 VSS.n10475 0.144
R29220 VSS.n10481 VSS.n10480 0.144
R29221 VSS.n17664 VSS.n17663 0.144
R29222 VSS.n17669 VSS.n17668 0.144
R29223 VSS.n17675 VSS.n17674 0.144
R29224 VSS.n17688 VSS.n17647 0.144
R29225 VSS.n17690 VSS.n17645 0.144
R29226 VSS.n17698 VSS.n17697 0.144
R29227 VSS.n16771 VSS.n16543 0.142
R29228 VSS.n16861 VSS.n16453 0.142
R29229 VSS.n16951 VSS.n16363 0.142
R29230 VSS.n17041 VSS.n16273 0.142
R29231 VSS.n17131 VSS.n16183 0.142
R29232 VSS.n17221 VSS.n16093 0.142
R29233 VSS.n17388 VSS.n17311 0.142
R29234 VSS.n11238 VSS.n11010 0.142
R29235 VSS.n11328 VSS.n10920 0.142
R29236 VSS.n11418 VSS.n10830 0.142
R29237 VSS.n13538 VSS.n10740 0.142
R29238 VSS.n13628 VSS.n10650 0.142
R29239 VSS.n13718 VSS.n10560 0.142
R29240 VSS.n13888 VSS.n13808 0.142
R29241 VSS.n9816 VSS.n9588 0.142
R29242 VSS.n9906 VSS.n9498 0.142
R29243 VSS.n9996 VSS.n9408 0.142
R29244 VSS.n10086 VSS.n9318 0.142
R29245 VSS.n10176 VSS.n9228 0.142
R29246 VSS.n10320 VSS.n10318 0.142
R29247 VSS.n9160 VSS.n8981 0.142
R29248 VSS.n6518 VSS.n6517 0.142
R29249 VSS.n6396 VSS.n6395 0.142
R29250 VSS.n6274 VSS.n6273 0.142
R29251 VSS.n6152 VSS.n6151 0.142
R29252 VSS.n6030 VSS.n6029 0.142
R29253 VSS.n5908 VSS.n5907 0.142
R29254 VSS.n5786 VSS.n5785 0.142
R29255 VSS.n724 VSS.n496 0.142
R29256 VSS.n814 VSS.n406 0.142
R29257 VSS.n904 VSS.n316 0.142
R29258 VSS.n994 VSS.n226 0.142
R29259 VSS.n1084 VSS.n136 0.142
R29260 VSS.n1174 VSS.n45 0.142
R29261 VSS.n6894 VSS.n6891 0.136
R29262 VSS.n1260 VSS.n1259 0.135
R29263 VSS.n14712 VSS.n14377 0.13
R29264 VSS.n14710 VSS.n14378 0.13
R29265 VSS.n14699 VSS.n14698 0.13
R29266 VSS.n14689 VSS.n14396 0.13
R29267 VSS.n14687 VSS.n14397 0.13
R29268 VSS.n14676 VSS.n14675 0.13
R29269 VSS.n14667 VSS.n14415 0.13
R29270 VSS.n14665 VSS.n14416 0.13
R29271 VSS.n14654 VSS.n14653 0.13
R29272 VSS.n14644 VSS.n14434 0.13
R29273 VSS.n14642 VSS.n14435 0.13
R29274 VSS.n14620 VSS.n14489 0.13
R29275 VSS.n14618 VSS.n14490 0.13
R29276 VSS.n14607 VSS.n14606 0.13
R29277 VSS.n14597 VSS.n14508 0.13
R29278 VSS.n14595 VSS.n14509 0.13
R29279 VSS.n14584 VSS.n14583 0.13
R29280 VSS.n14575 VSS.n14527 0.13
R29281 VSS.n14573 VSS.n14528 0.13
R29282 VSS.n14562 VSS.n14561 0.13
R29283 VSS.n14552 VSS.n14550 0.13
R29284 VSS.n14869 VSS.n14307 0.13
R29285 VSS.n14881 VSS.n14293 0.13
R29286 VSS.n14893 VSS.n14892 0.13
R29287 VSS.n14905 VSS.n14903 0.13
R29288 VSS.n14914 VSS.n14277 0.13
R29289 VSS.n14916 VSS.n14272 0.13
R29290 VSS.n14928 VSS.n14927 0.13
R29291 VSS.n14939 VSS.n14937 0.13
R29292 VSS.n14948 VSS.n14256 0.13
R29293 VSS.n14950 VSS.n14251 0.13
R29294 VSS.n14962 VSS.n14961 0.13
R29295 VSS.n15327 VSS.n14972 0.13
R29296 VSS.n15313 VSS.n14986 0.13
R29297 VSS.n15311 VSS.n14987 0.13
R29298 VSS.n15300 VSS.n15299 0.13
R29299 VSS.n15290 VSS.n15005 0.13
R29300 VSS.n15288 VSS.n15006 0.13
R29301 VSS.n15277 VSS.n15276 0.13
R29302 VSS.n15268 VSS.n15024 0.13
R29303 VSS.n15266 VSS.n15025 0.13
R29304 VSS.n15255 VSS.n15254 0.13
R29305 VSS.n15245 VSS.n15043 0.13
R29306 VSS.n15243 VSS.n15044 0.13
R29307 VSS.n15221 VSS.n15098 0.13
R29308 VSS.n15219 VSS.n15099 0.13
R29309 VSS.n15208 VSS.n15207 0.13
R29310 VSS.n15198 VSS.n15117 0.13
R29311 VSS.n15196 VSS.n15118 0.13
R29312 VSS.n15185 VSS.n15184 0.13
R29313 VSS.n15176 VSS.n15136 0.13
R29314 VSS.n15174 VSS.n15137 0.13
R29315 VSS.n15163 VSS.n15162 0.13
R29316 VSS.n15153 VSS.n15152 0.13
R29317 VSS.n15450 VSS.n15449 0.13
R29318 VSS.n15468 VSS.n15466 0.13
R29319 VSS.n15477 VSS.n14121 0.13
R29320 VSS.n15479 VSS.n14116 0.13
R29321 VSS.n15491 VSS.n15490 0.13
R29322 VSS.n15503 VSS.n15501 0.13
R29323 VSS.n15511 VSS.n14100 0.13
R29324 VSS.n15513 VSS.n14095 0.13
R29325 VSS.n15525 VSS.n15524 0.13
R29326 VSS.n15537 VSS.n15535 0.13
R29327 VSS.n15546 VSS.n14079 0.13
R29328 VSS.n15548 VSS.n14073 0.13
R29329 VSS.n15880 VSS.n15573 0.13
R29330 VSS.n15878 VSS.n15574 0.13
R29331 VSS.n15867 VSS.n15866 0.13
R29332 VSS.n15857 VSS.n15592 0.13
R29333 VSS.n15855 VSS.n15593 0.13
R29334 VSS.n15844 VSS.n15843 0.13
R29335 VSS.n15835 VSS.n15611 0.13
R29336 VSS.n15833 VSS.n15612 0.13
R29337 VSS.n15822 VSS.n15821 0.13
R29338 VSS.n15812 VSS.n15630 0.13
R29339 VSS.n15810 VSS.n15631 0.13
R29340 VSS.n15788 VSS.n15685 0.13
R29341 VSS.n15786 VSS.n15686 0.13
R29342 VSS.n15775 VSS.n15774 0.13
R29343 VSS.n15765 VSS.n15704 0.13
R29344 VSS.n15763 VSS.n15705 0.13
R29345 VSS.n15752 VSS.n15751 0.13
R29346 VSS.n15743 VSS.n15723 0.13
R29347 VSS.n15741 VSS.n15724 0.13
R29348 VSS.n16013 VSS.n14007 0.13
R29349 VSS.n16011 VSS.n14008 0.13
R29350 VSS.n16757 VSS.n16689 0.13
R29351 VSS.n16755 VSS.n16690 0.13
R29352 VSS.n16746 VSS.n16745 0.13
R29353 VSS.n16740 VSS.n16739 0.13
R29354 VSS.n16734 VSS.n16733 0.13
R29355 VSS.n16728 VSS.n16727 0.13
R29356 VSS.n16722 VSS.n16721 0.13
R29357 VSS.n16717 VSS.n16716 0.13
R29358 VSS.n16847 VSS.n16779 0.13
R29359 VSS.n16845 VSS.n16780 0.13
R29360 VSS.n16836 VSS.n16835 0.13
R29361 VSS.n16830 VSS.n16829 0.13
R29362 VSS.n16824 VSS.n16823 0.13
R29363 VSS.n16818 VSS.n16817 0.13
R29364 VSS.n16812 VSS.n16811 0.13
R29365 VSS.n16807 VSS.n16806 0.13
R29366 VSS.n16937 VSS.n16869 0.13
R29367 VSS.n16935 VSS.n16870 0.13
R29368 VSS.n16926 VSS.n16925 0.13
R29369 VSS.n16920 VSS.n16919 0.13
R29370 VSS.n16914 VSS.n16913 0.13
R29371 VSS.n16908 VSS.n16907 0.13
R29372 VSS.n16902 VSS.n16901 0.13
R29373 VSS.n16897 VSS.n16896 0.13
R29374 VSS.n17027 VSS.n16959 0.13
R29375 VSS.n17025 VSS.n16960 0.13
R29376 VSS.n17016 VSS.n17015 0.13
R29377 VSS.n17010 VSS.n17009 0.13
R29378 VSS.n17004 VSS.n17003 0.13
R29379 VSS.n16998 VSS.n16997 0.13
R29380 VSS.n16992 VSS.n16991 0.13
R29381 VSS.n16987 VSS.n16986 0.13
R29382 VSS.n17117 VSS.n17049 0.13
R29383 VSS.n17115 VSS.n17050 0.13
R29384 VSS.n17106 VSS.n17105 0.13
R29385 VSS.n17100 VSS.n17099 0.13
R29386 VSS.n17094 VSS.n17093 0.13
R29387 VSS.n17088 VSS.n17087 0.13
R29388 VSS.n17082 VSS.n17081 0.13
R29389 VSS.n17077 VSS.n17076 0.13
R29390 VSS.n17207 VSS.n17139 0.13
R29391 VSS.n17205 VSS.n17140 0.13
R29392 VSS.n17196 VSS.n17195 0.13
R29393 VSS.n17190 VSS.n17189 0.13
R29394 VSS.n17184 VSS.n17183 0.13
R29395 VSS.n17178 VSS.n17177 0.13
R29396 VSS.n17172 VSS.n17171 0.13
R29397 VSS.n17167 VSS.n17166 0.13
R29398 VSS.n17297 VSS.n17229 0.13
R29399 VSS.n17295 VSS.n17230 0.13
R29400 VSS.n17286 VSS.n17285 0.13
R29401 VSS.n17280 VSS.n17279 0.13
R29402 VSS.n17274 VSS.n17273 0.13
R29403 VSS.n17268 VSS.n17267 0.13
R29404 VSS.n17262 VSS.n17261 0.13
R29405 VSS.n17257 VSS.n17256 0.13
R29406 VSS.n17390 VSS.n16050 0.13
R29407 VSS.n17453 VSS.n17398 0.13
R29408 VSS.n17451 VSS.n17399 0.13
R29409 VSS.n17442 VSS.n17441 0.13
R29410 VSS.n17436 VSS.n17435 0.13
R29411 VSS.n17430 VSS.n17429 0.13
R29412 VSS.n17424 VSS.n17423 0.13
R29413 VSS.n12803 VSS.n12802 0.13
R29414 VSS.n12815 VSS.n12813 0.13
R29415 VSS.n12824 VSS.n12704 0.13
R29416 VSS.n12826 VSS.n12699 0.13
R29417 VSS.n12838 VSS.n12837 0.13
R29418 VSS.n12850 VSS.n12848 0.13
R29419 VSS.n12858 VSS.n12683 0.13
R29420 VSS.n12860 VSS.n12678 0.13
R29421 VSS.n12872 VSS.n12871 0.13
R29422 VSS.n12884 VSS.n12883 0.13
R29423 VSS.n13061 VSS.n12661 0.13
R29424 VSS.n13049 VSS.n12895 0.13
R29425 VSS.n13038 VSS.n13037 0.13
R29426 VSS.n13028 VSS.n12914 0.13
R29427 VSS.n13026 VSS.n12915 0.13
R29428 VSS.n13015 VSS.n13014 0.13
R29429 VSS.n13006 VSS.n12933 0.13
R29430 VSS.n13004 VSS.n12934 0.13
R29431 VSS.n12993 VSS.n12992 0.13
R29432 VSS.n12983 VSS.n12952 0.13
R29433 VSS.n12981 VSS.n12953 0.13
R29434 VSS.n12970 VSS.n12969 0.13
R29435 VSS.n13160 VSS.n13159 0.13
R29436 VSS.n13172 VSS.n13170 0.13
R29437 VSS.n13181 VSS.n12563 0.13
R29438 VSS.n13183 VSS.n12558 0.13
R29439 VSS.n13195 VSS.n13194 0.13
R29440 VSS.n13207 VSS.n13205 0.13
R29441 VSS.n13215 VSS.n12542 0.13
R29442 VSS.n13217 VSS.n12537 0.13
R29443 VSS.n13229 VSS.n13228 0.13
R29444 VSS.n13241 VSS.n13240 0.13
R29445 VSS.n13310 VSS.n12520 0.13
R29446 VSS.n13298 VSS.n13252 0.13
R29447 VSS.n13287 VSS.n13286 0.13
R29448 VSS.n13277 VSS.n13275 0.13
R29449 VSS.n13447 VSS.n11441 0.13
R29450 VSS.n13445 VSS.n11442 0.13
R29451 VSS.n13435 VSS.n13434 0.13
R29452 VSS.n13425 VSS.n11460 0.13
R29453 VSS.n13423 VSS.n11461 0.13
R29454 VSS.n13412 VSS.n13411 0.13
R29455 VSS.n13402 VSS.n11479 0.13
R29456 VSS.n11681 VSS.n11680 0.13
R29457 VSS.n11693 VSS.n11691 0.13
R29458 VSS.n11702 VSS.n11654 0.13
R29459 VSS.n11704 VSS.n11649 0.13
R29460 VSS.n11716 VSS.n11715 0.13
R29461 VSS.n11728 VSS.n11726 0.13
R29462 VSS.n11736 VSS.n11633 0.13
R29463 VSS.n11738 VSS.n11628 0.13
R29464 VSS.n11750 VSS.n11749 0.13
R29465 VSS.n11762 VSS.n11760 0.13
R29466 VSS.n11771 VSS.n11611 0.13
R29467 VSS.n11815 VSS.n11598 0.13
R29468 VSS.n11827 VSS.n11826 0.13
R29469 VSS.n11839 VSS.n11837 0.13
R29470 VSS.n11848 VSS.n11582 0.13
R29471 VSS.n11850 VSS.n11577 0.13
R29472 VSS.n11862 VSS.n11861 0.13
R29473 VSS.n11873 VSS.n11871 0.13
R29474 VSS.n11882 VSS.n11561 0.13
R29475 VSS.n11884 VSS.n11556 0.13
R29476 VSS.n11896 VSS.n11895 0.13
R29477 VSS.n12402 VSS.n11906 0.13
R29478 VSS.n12388 VSS.n11920 0.13
R29479 VSS.n12386 VSS.n11921 0.13
R29480 VSS.n12375 VSS.n12374 0.13
R29481 VSS.n12365 VSS.n11939 0.13
R29482 VSS.n12363 VSS.n11940 0.13
R29483 VSS.n12352 VSS.n12351 0.13
R29484 VSS.n12343 VSS.n11958 0.13
R29485 VSS.n12341 VSS.n11959 0.13
R29486 VSS.n12330 VSS.n12329 0.13
R29487 VSS.n12320 VSS.n11977 0.13
R29488 VSS.n12318 VSS.n11978 0.13
R29489 VSS.n12296 VSS.n11999 0.13
R29490 VSS.n12294 VSS.n12000 0.13
R29491 VSS.n12283 VSS.n12282 0.13
R29492 VSS.n12273 VSS.n12018 0.13
R29493 VSS.n12271 VSS.n12019 0.13
R29494 VSS.n12260 VSS.n12259 0.13
R29495 VSS.n12251 VSS.n12037 0.13
R29496 VSS.n12249 VSS.n12038 0.13
R29497 VSS.n12238 VSS.n12237 0.13
R29498 VSS.n12228 VSS.n12056 0.13
R29499 VSS.n12226 VSS.n12057 0.13
R29500 VSS.n11225 VSS.n11156 0.13
R29501 VSS.n11223 VSS.n11157 0.13
R29502 VSS.n11214 VSS.n11213 0.13
R29503 VSS.n11208 VSS.n11207 0.13
R29504 VSS.n11202 VSS.n11201 0.13
R29505 VSS.n11196 VSS.n11195 0.13
R29506 VSS.n11191 VSS.n11190 0.13
R29507 VSS.n11185 VSS.n11184 0.13
R29508 VSS.n11315 VSS.n11246 0.13
R29509 VSS.n11313 VSS.n11247 0.13
R29510 VSS.n11304 VSS.n11303 0.13
R29511 VSS.n11298 VSS.n11297 0.13
R29512 VSS.n11292 VSS.n11291 0.13
R29513 VSS.n11286 VSS.n11285 0.13
R29514 VSS.n11281 VSS.n11280 0.13
R29515 VSS.n11275 VSS.n11274 0.13
R29516 VSS.n11405 VSS.n11336 0.13
R29517 VSS.n11403 VSS.n11337 0.13
R29518 VSS.n11394 VSS.n11393 0.13
R29519 VSS.n11388 VSS.n11387 0.13
R29520 VSS.n11382 VSS.n11381 0.13
R29521 VSS.n11376 VSS.n11375 0.13
R29522 VSS.n11371 VSS.n11370 0.13
R29523 VSS.n11365 VSS.n11364 0.13
R29524 VSS.n13525 VSS.n11426 0.13
R29525 VSS.n13523 VSS.n11427 0.13
R29526 VSS.n13507 VSS.n13506 0.13
R29527 VSS.n13501 VSS.n13500 0.13
R29528 VSS.n13495 VSS.n13494 0.13
R29529 VSS.n13490 VSS.n13489 0.13
R29530 VSS.n13484 VSS.n13483 0.13
R29531 VSS.n13615 VSS.n13546 0.13
R29532 VSS.n13613 VSS.n13547 0.13
R29533 VSS.n13604 VSS.n13603 0.13
R29534 VSS.n13598 VSS.n13597 0.13
R29535 VSS.n13592 VSS.n13591 0.13
R29536 VSS.n13586 VSS.n13585 0.13
R29537 VSS.n13581 VSS.n13580 0.13
R29538 VSS.n13575 VSS.n13574 0.13
R29539 VSS.n13705 VSS.n13636 0.13
R29540 VSS.n13703 VSS.n13637 0.13
R29541 VSS.n13694 VSS.n13693 0.13
R29542 VSS.n13688 VSS.n13687 0.13
R29543 VSS.n13682 VSS.n13681 0.13
R29544 VSS.n13676 VSS.n13675 0.13
R29545 VSS.n13671 VSS.n13670 0.13
R29546 VSS.n13665 VSS.n13664 0.13
R29547 VSS.n13795 VSS.n13726 0.13
R29548 VSS.n13793 VSS.n13727 0.13
R29549 VSS.n13784 VSS.n13783 0.13
R29550 VSS.n13778 VSS.n13777 0.13
R29551 VSS.n13772 VSS.n13771 0.13
R29552 VSS.n13766 VSS.n13765 0.13
R29553 VSS.n13761 VSS.n13760 0.13
R29554 VSS.n13755 VSS.n13754 0.13
R29555 VSS.n13890 VSS.n10517 0.13
R29556 VSS.n13945 VSS.n13898 0.13
R29557 VSS.n13943 VSS.n13899 0.13
R29558 VSS.n13934 VSS.n13933 0.13
R29559 VSS.n13928 VSS.n13927 0.13
R29560 VSS.n13922 VSS.n13921 0.13
R29561 VSS.n13916 VSS.n10491 0.13
R29562 VSS.n7826 VSS.n7684 0.13
R29563 VSS.n7824 VSS.n7685 0.13
R29564 VSS.n7813 VSS.n7812 0.13
R29565 VSS.n7803 VSS.n7703 0.13
R29566 VSS.n7801 VSS.n7704 0.13
R29567 VSS.n7790 VSS.n7789 0.13
R29568 VSS.n7781 VSS.n7722 0.13
R29569 VSS.n7779 VSS.n7723 0.13
R29570 VSS.n7768 VSS.n7767 0.13
R29571 VSS.n7758 VSS.n7741 0.13
R29572 VSS.n7756 VSS.n7742 0.13
R29573 VSS.n7926 VSS.n7592 0.13
R29574 VSS.n7938 VSS.n7937 0.13
R29575 VSS.n7950 VSS.n7948 0.13
R29576 VSS.n7959 VSS.n7576 0.13
R29577 VSS.n7961 VSS.n7571 0.13
R29578 VSS.n7973 VSS.n7972 0.13
R29579 VSS.n7984 VSS.n7982 0.13
R29580 VSS.n7993 VSS.n7555 0.13
R29581 VSS.n7995 VSS.n7550 0.13
R29582 VSS.n8007 VSS.n8006 0.13
R29583 VSS.n8188 VSS.n8017 0.13
R29584 VSS.n8030 VSS.n8029 0.13
R29585 VSS.n8166 VSS.n8038 0.13
R29586 VSS.n8164 VSS.n8039 0.13
R29587 VSS.n8153 VSS.n8152 0.13
R29588 VSS.n8143 VSS.n8057 0.13
R29589 VSS.n8141 VSS.n8058 0.13
R29590 VSS.n8131 VSS.n8130 0.13
R29591 VSS.n8121 VSS.n8076 0.13
R29592 VSS.n8119 VSS.n8077 0.13
R29593 VSS.n8108 VSS.n8107 0.13
R29594 VSS.n8098 VSS.n8094 0.13
R29595 VSS.n8284 VSS.n7452 0.13
R29596 VSS.n8296 VSS.n8295 0.13
R29597 VSS.n8308 VSS.n8306 0.13
R29598 VSS.n8317 VSS.n7436 0.13
R29599 VSS.n8319 VSS.n7431 0.13
R29600 VSS.n8331 VSS.n8330 0.13
R29601 VSS.n8342 VSS.n8340 0.13
R29602 VSS.n8351 VSS.n7415 0.13
R29603 VSS.n8353 VSS.n7410 0.13
R29604 VSS.n8365 VSS.n8364 0.13
R29605 VSS.n8546 VSS.n8375 0.13
R29606 VSS.n8388 VSS.n8387 0.13
R29607 VSS.n8524 VSS.n8396 0.13
R29608 VSS.n8522 VSS.n8397 0.13
R29609 VSS.n8511 VSS.n8510 0.13
R29610 VSS.n8501 VSS.n8415 0.13
R29611 VSS.n8499 VSS.n8416 0.13
R29612 VSS.n8489 VSS.n8488 0.13
R29613 VSS.n8479 VSS.n8434 0.13
R29614 VSS.n8477 VSS.n8435 0.13
R29615 VSS.n8466 VSS.n8465 0.13
R29616 VSS.n8456 VSS.n8452 0.13
R29617 VSS.n8642 VSS.n7312 0.13
R29618 VSS.n8654 VSS.n8653 0.13
R29619 VSS.n8666 VSS.n8664 0.13
R29620 VSS.n8675 VSS.n7296 0.13
R29621 VSS.n8677 VSS.n7291 0.13
R29622 VSS.n8689 VSS.n8688 0.13
R29623 VSS.n8700 VSS.n8698 0.13
R29624 VSS.n8709 VSS.n7275 0.13
R29625 VSS.n8711 VSS.n7270 0.13
R29626 VSS.n8723 VSS.n8722 0.13
R29627 VSS.n8768 VSS.n8733 0.13
R29628 VSS.n8747 VSS.n8745 0.13
R29629 VSS.n8919 VSS.n6913 0.13
R29630 VSS.n8917 VSS.n6914 0.13
R29631 VSS.n8906 VSS.n8905 0.13
R29632 VSS.n8897 VSS.n6932 0.13
R29633 VSS.n8895 VSS.n6933 0.13
R29634 VSS.n8884 VSS.n8883 0.13
R29635 VSS.n8874 VSS.n6951 0.13
R29636 VSS.n8872 VSS.n6952 0.13
R29637 VSS.n8861 VSS.n8860 0.13
R29638 VSS.n7084 VSS.n7082 0.13
R29639 VSS.n7093 VSS.n7056 0.13
R29640 VSS.n7095 VSS.n7051 0.13
R29641 VSS.n7107 VSS.n7106 0.13
R29642 VSS.n7119 VSS.n7117 0.13
R29643 VSS.n7127 VSS.n7035 0.13
R29644 VSS.n7129 VSS.n7030 0.13
R29645 VSS.n7141 VSS.n7140 0.13
R29646 VSS.n7153 VSS.n7151 0.13
R29647 VSS.n7162 VSS.n7014 0.13
R29648 VSS.n7164 VSS.n7008 0.13
R29649 VSS.n9802 VSS.n9734 0.13
R29650 VSS.n9800 VSS.n9735 0.13
R29651 VSS.n9791 VSS.n9790 0.13
R29652 VSS.n9785 VSS.n9784 0.13
R29653 VSS.n9779 VSS.n9778 0.13
R29654 VSS.n9773 VSS.n9772 0.13
R29655 VSS.n9767 VSS.n9766 0.13
R29656 VSS.n9762 VSS.n9761 0.13
R29657 VSS.n9892 VSS.n9824 0.13
R29658 VSS.n9890 VSS.n9825 0.13
R29659 VSS.n9881 VSS.n9880 0.13
R29660 VSS.n9875 VSS.n9874 0.13
R29661 VSS.n9869 VSS.n9868 0.13
R29662 VSS.n9863 VSS.n9862 0.13
R29663 VSS.n9857 VSS.n9856 0.13
R29664 VSS.n9852 VSS.n9851 0.13
R29665 VSS.n9982 VSS.n9914 0.13
R29666 VSS.n9980 VSS.n9915 0.13
R29667 VSS.n9971 VSS.n9970 0.13
R29668 VSS.n9965 VSS.n9964 0.13
R29669 VSS.n9959 VSS.n9958 0.13
R29670 VSS.n9953 VSS.n9952 0.13
R29671 VSS.n9947 VSS.n9946 0.13
R29672 VSS.n9942 VSS.n9941 0.13
R29673 VSS.n10072 VSS.n10004 0.13
R29674 VSS.n10070 VSS.n10005 0.13
R29675 VSS.n10061 VSS.n10060 0.13
R29676 VSS.n10055 VSS.n10054 0.13
R29677 VSS.n10049 VSS.n10048 0.13
R29678 VSS.n10043 VSS.n10042 0.13
R29679 VSS.n10037 VSS.n10036 0.13
R29680 VSS.n10032 VSS.n10031 0.13
R29681 VSS.n10162 VSS.n10094 0.13
R29682 VSS.n10160 VSS.n10095 0.13
R29683 VSS.n10151 VSS.n10150 0.13
R29684 VSS.n10145 VSS.n10144 0.13
R29685 VSS.n10139 VSS.n10138 0.13
R29686 VSS.n10133 VSS.n10132 0.13
R29687 VSS.n10127 VSS.n10126 0.13
R29688 VSS.n10122 VSS.n10121 0.13
R29689 VSS.n10252 VSS.n10184 0.13
R29690 VSS.n10250 VSS.n10185 0.13
R29691 VSS.n10241 VSS.n10240 0.13
R29692 VSS.n10235 VSS.n10234 0.13
R29693 VSS.n10229 VSS.n10228 0.13
R29694 VSS.n10223 VSS.n10222 0.13
R29695 VSS.n10217 VSS.n10216 0.13
R29696 VSS.n10212 VSS.n10211 0.13
R29697 VSS.n8940 VSS.n8939 0.13
R29698 VSS.n8946 VSS.n8945 0.13
R29699 VSS.n8952 VSS.n8951 0.13
R29700 VSS.n8957 VSS.n8956 0.13
R29701 VSS.n8964 VSS.n8963 0.13
R29702 VSS.n8970 VSS.n8969 0.13
R29703 VSS.n8976 VSS.n8975 0.13
R29704 VSS.n9041 VSS.n9040 0.13
R29705 VSS.n9049 VSS.n9048 0.13
R29706 VSS.n9057 VSS.n9056 0.13
R29707 VSS.n9065 VSS.n9064 0.13
R29708 VSS.n9073 VSS.n9072 0.13
R29709 VSS.n9081 VSS.n9080 0.13
R29710 VSS.n9089 VSS.n9088 0.13
R29711 VSS.n9152 VSS.n9096 0.13
R29712 VSS.n4256 VSS.n4255 0.13
R29713 VSS.n4268 VSS.n4266 0.13
R29714 VSS.n4277 VSS.n4157 0.13
R29715 VSS.n4279 VSS.n4152 0.13
R29716 VSS.n4291 VSS.n4290 0.13
R29717 VSS.n4303 VSS.n4301 0.13
R29718 VSS.n4311 VSS.n4136 0.13
R29719 VSS.n4313 VSS.n4131 0.13
R29720 VSS.n4325 VSS.n4324 0.13
R29721 VSS.n4337 VSS.n4336 0.13
R29722 VSS.n4514 VSS.n4114 0.13
R29723 VSS.n4502 VSS.n4348 0.13
R29724 VSS.n4491 VSS.n4490 0.13
R29725 VSS.n4481 VSS.n4367 0.13
R29726 VSS.n4479 VSS.n4368 0.13
R29727 VSS.n4468 VSS.n4467 0.13
R29728 VSS.n4459 VSS.n4386 0.13
R29729 VSS.n4457 VSS.n4387 0.13
R29730 VSS.n4446 VSS.n4445 0.13
R29731 VSS.n4436 VSS.n4405 0.13
R29732 VSS.n4434 VSS.n4406 0.13
R29733 VSS.n4423 VSS.n4422 0.13
R29734 VSS.n4613 VSS.n4612 0.13
R29735 VSS.n4625 VSS.n4623 0.13
R29736 VSS.n4634 VSS.n4016 0.13
R29737 VSS.n4636 VSS.n4011 0.13
R29738 VSS.n4648 VSS.n4647 0.13
R29739 VSS.n4660 VSS.n4658 0.13
R29740 VSS.n4668 VSS.n3995 0.13
R29741 VSS.n4670 VSS.n3990 0.13
R29742 VSS.n4682 VSS.n4681 0.13
R29743 VSS.n4694 VSS.n4693 0.13
R29744 VSS.n4871 VSS.n3973 0.13
R29745 VSS.n4859 VSS.n4705 0.13
R29746 VSS.n4848 VSS.n4847 0.13
R29747 VSS.n4838 VSS.n4724 0.13
R29748 VSS.n4836 VSS.n4725 0.13
R29749 VSS.n4825 VSS.n4824 0.13
R29750 VSS.n4816 VSS.n4743 0.13
R29751 VSS.n4814 VSS.n4744 0.13
R29752 VSS.n4803 VSS.n4802 0.13
R29753 VSS.n4793 VSS.n4762 0.13
R29754 VSS.n4791 VSS.n4763 0.13
R29755 VSS.n4780 VSS.n4779 0.13
R29756 VSS.n4970 VSS.n4969 0.13
R29757 VSS.n4982 VSS.n4980 0.13
R29758 VSS.n4991 VSS.n3875 0.13
R29759 VSS.n4993 VSS.n3870 0.13
R29760 VSS.n5005 VSS.n5004 0.13
R29761 VSS.n5017 VSS.n5015 0.13
R29762 VSS.n5025 VSS.n3854 0.13
R29763 VSS.n5027 VSS.n3849 0.13
R29764 VSS.n5039 VSS.n5038 0.13
R29765 VSS.n5051 VSS.n5050 0.13
R29766 VSS.n5228 VSS.n3832 0.13
R29767 VSS.n5216 VSS.n5062 0.13
R29768 VSS.n5205 VSS.n5204 0.13
R29769 VSS.n5195 VSS.n5081 0.13
R29770 VSS.n5193 VSS.n5082 0.13
R29771 VSS.n5182 VSS.n5181 0.13
R29772 VSS.n5173 VSS.n5100 0.13
R29773 VSS.n5171 VSS.n5101 0.13
R29774 VSS.n5160 VSS.n5159 0.13
R29775 VSS.n5150 VSS.n5119 0.13
R29776 VSS.n5148 VSS.n5120 0.13
R29777 VSS.n5137 VSS.n5136 0.13
R29778 VSS.n5327 VSS.n5326 0.13
R29779 VSS.n5339 VSS.n5337 0.13
R29780 VSS.n5348 VSS.n3734 0.13
R29781 VSS.n5350 VSS.n3729 0.13
R29782 VSS.n5362 VSS.n5361 0.13
R29783 VSS.n5374 VSS.n5372 0.13
R29784 VSS.n5382 VSS.n3713 0.13
R29785 VSS.n5384 VSS.n3708 0.13
R29786 VSS.n5396 VSS.n5395 0.13
R29787 VSS.n5408 VSS.n5407 0.13
R29788 VSS.n5574 VSS.n3691 0.13
R29789 VSS.n5562 VSS.n5419 0.13
R29790 VSS.n5551 VSS.n5550 0.13
R29791 VSS.n5541 VSS.n5438 0.13
R29792 VSS.n5539 VSS.n5439 0.13
R29793 VSS.n5528 VSS.n5527 0.13
R29794 VSS.n5519 VSS.n5457 0.13
R29795 VSS.n5517 VSS.n5458 0.13
R29796 VSS.n5506 VSS.n5505 0.13
R29797 VSS.n5496 VSS.n5476 0.13
R29798 VSS.n5494 VSS.n5477 0.13
R29799 VSS.n3174 VSS.n3137 0.13
R29800 VSS.n3181 VSS.n3180 0.13
R29801 VSS.n3189 VSS.n3188 0.13
R29802 VSS.n3197 VSS.n3196 0.13
R29803 VSS.n3205 VSS.n3204 0.13
R29804 VSS.n3213 VSS.n3212 0.13
R29805 VSS.n3221 VSS.n3220 0.13
R29806 VSS.n6594 VSS.n3228 0.13
R29807 VSS.n3239 VSS.n3238 0.13
R29808 VSS.n3245 VSS.n3244 0.13
R29809 VSS.n3251 VSS.n3250 0.13
R29810 VSS.n3257 VSS.n3256 0.13
R29811 VSS.n3262 VSS.n3261 0.13
R29812 VSS.n3269 VSS.n3268 0.13
R29813 VSS.n3275 VSS.n3274 0.13
R29814 VSS.n3281 VSS.n3280 0.13
R29815 VSS.n3297 VSS.n3296 0.13
R29816 VSS.n3303 VSS.n3302 0.13
R29817 VSS.n3309 VSS.n3308 0.13
R29818 VSS.n3315 VSS.n3314 0.13
R29819 VSS.n3320 VSS.n3319 0.13
R29820 VSS.n3327 VSS.n3326 0.13
R29821 VSS.n3333 VSS.n3332 0.13
R29822 VSS.n3339 VSS.n3338 0.13
R29823 VSS.n3355 VSS.n3354 0.13
R29824 VSS.n3361 VSS.n3360 0.13
R29825 VSS.n3367 VSS.n3366 0.13
R29826 VSS.n3373 VSS.n3372 0.13
R29827 VSS.n3378 VSS.n3377 0.13
R29828 VSS.n3385 VSS.n3384 0.13
R29829 VSS.n3391 VSS.n3390 0.13
R29830 VSS.n3397 VSS.n3396 0.13
R29831 VSS.n3413 VSS.n3412 0.13
R29832 VSS.n3419 VSS.n3418 0.13
R29833 VSS.n3425 VSS.n3424 0.13
R29834 VSS.n3431 VSS.n3430 0.13
R29835 VSS.n3436 VSS.n3435 0.13
R29836 VSS.n3443 VSS.n3442 0.13
R29837 VSS.n3449 VSS.n3448 0.13
R29838 VSS.n3455 VSS.n3454 0.13
R29839 VSS.n3471 VSS.n3470 0.13
R29840 VSS.n3477 VSS.n3476 0.13
R29841 VSS.n3483 VSS.n3482 0.13
R29842 VSS.n3489 VSS.n3488 0.13
R29843 VSS.n3494 VSS.n3493 0.13
R29844 VSS.n3501 VSS.n3500 0.13
R29845 VSS.n3507 VSS.n3506 0.13
R29846 VSS.n3513 VSS.n3512 0.13
R29847 VSS.n3529 VSS.n3528 0.13
R29848 VSS.n3535 VSS.n3534 0.13
R29849 VSS.n3541 VSS.n3540 0.13
R29850 VSS.n3547 VSS.n3546 0.13
R29851 VSS.n3552 VSS.n3551 0.13
R29852 VSS.n3559 VSS.n3558 0.13
R29853 VSS.n3565 VSS.n3564 0.13
R29854 VSS.n3571 VSS.n3570 0.13
R29855 VSS.n3587 VSS.n3586 0.13
R29856 VSS.n3593 VSS.n3592 0.13
R29857 VSS.n3599 VSS.n3598 0.13
R29858 VSS.n3605 VSS.n3604 0.13
R29859 VSS.n3610 VSS.n3609 0.13
R29860 VSS.n3617 VSS.n3616 0.13
R29861 VSS.n3623 VSS.n3622 0.13
R29862 VSS.n3629 VSS.n3628 0.13
R29863 VSS.n1953 VSS.n1618 0.13
R29864 VSS.n1951 VSS.n1619 0.13
R29865 VSS.n1940 VSS.n1939 0.13
R29866 VSS.n1930 VSS.n1637 0.13
R29867 VSS.n1928 VSS.n1638 0.13
R29868 VSS.n1917 VSS.n1916 0.13
R29869 VSS.n1908 VSS.n1656 0.13
R29870 VSS.n1906 VSS.n1657 0.13
R29871 VSS.n1895 VSS.n1894 0.13
R29872 VSS.n1885 VSS.n1675 0.13
R29873 VSS.n1883 VSS.n1676 0.13
R29874 VSS.n1861 VSS.n1730 0.13
R29875 VSS.n1859 VSS.n1731 0.13
R29876 VSS.n1848 VSS.n1847 0.13
R29877 VSS.n1838 VSS.n1749 0.13
R29878 VSS.n1836 VSS.n1750 0.13
R29879 VSS.n1825 VSS.n1824 0.13
R29880 VSS.n1816 VSS.n1768 0.13
R29881 VSS.n1814 VSS.n1769 0.13
R29882 VSS.n1803 VSS.n1802 0.13
R29883 VSS.n1793 VSS.n1791 0.13
R29884 VSS.n2110 VSS.n1548 0.13
R29885 VSS.n2122 VSS.n1534 0.13
R29886 VSS.n2134 VSS.n2133 0.13
R29887 VSS.n2146 VSS.n2144 0.13
R29888 VSS.n2155 VSS.n1518 0.13
R29889 VSS.n2157 VSS.n1513 0.13
R29890 VSS.n2169 VSS.n2168 0.13
R29891 VSS.n2180 VSS.n2178 0.13
R29892 VSS.n2189 VSS.n1497 0.13
R29893 VSS.n2191 VSS.n1492 0.13
R29894 VSS.n2203 VSS.n2202 0.13
R29895 VSS.n2568 VSS.n2213 0.13
R29896 VSS.n2554 VSS.n2227 0.13
R29897 VSS.n2552 VSS.n2228 0.13
R29898 VSS.n2541 VSS.n2540 0.13
R29899 VSS.n2531 VSS.n2246 0.13
R29900 VSS.n2529 VSS.n2247 0.13
R29901 VSS.n2518 VSS.n2517 0.13
R29902 VSS.n2509 VSS.n2265 0.13
R29903 VSS.n2507 VSS.n2266 0.13
R29904 VSS.n2496 VSS.n2495 0.13
R29905 VSS.n2486 VSS.n2284 0.13
R29906 VSS.n2484 VSS.n2285 0.13
R29907 VSS.n2462 VSS.n2339 0.13
R29908 VSS.n2460 VSS.n2340 0.13
R29909 VSS.n2449 VSS.n2448 0.13
R29910 VSS.n2439 VSS.n2358 0.13
R29911 VSS.n2437 VSS.n2359 0.13
R29912 VSS.n2426 VSS.n2425 0.13
R29913 VSS.n2417 VSS.n2377 0.13
R29914 VSS.n2415 VSS.n2378 0.13
R29915 VSS.n2404 VSS.n2403 0.13
R29916 VSS.n2394 VSS.n2393 0.13
R29917 VSS.n2691 VSS.n2690 0.13
R29918 VSS.n2709 VSS.n2707 0.13
R29919 VSS.n2718 VSS.n1362 0.13
R29920 VSS.n2720 VSS.n1357 0.13
R29921 VSS.n2732 VSS.n2731 0.13
R29922 VSS.n2744 VSS.n2742 0.13
R29923 VSS.n2752 VSS.n1341 0.13
R29924 VSS.n2754 VSS.n1336 0.13
R29925 VSS.n2766 VSS.n2765 0.13
R29926 VSS.n2778 VSS.n2776 0.13
R29927 VSS.n2787 VSS.n1320 0.13
R29928 VSS.n2789 VSS.n1314 0.13
R29929 VSS.n2954 VSS.n2814 0.13
R29930 VSS.n2952 VSS.n2815 0.13
R29931 VSS.n2941 VSS.n2940 0.13
R29932 VSS.n2931 VSS.n2833 0.13
R29933 VSS.n2929 VSS.n2834 0.13
R29934 VSS.n2918 VSS.n2917 0.13
R29935 VSS.n2909 VSS.n2852 0.13
R29936 VSS.n2907 VSS.n2853 0.13
R29937 VSS.n2896 VSS.n2895 0.13
R29938 VSS.n2886 VSS.n2871 0.13
R29939 VSS.n2884 VSS.n2872 0.13
R29940 VSS.n710 VSS.n642 0.13
R29941 VSS.n708 VSS.n643 0.13
R29942 VSS.n699 VSS.n698 0.13
R29943 VSS.n693 VSS.n692 0.13
R29944 VSS.n687 VSS.n686 0.13
R29945 VSS.n681 VSS.n680 0.13
R29946 VSS.n675 VSS.n674 0.13
R29947 VSS.n670 VSS.n669 0.13
R29948 VSS.n800 VSS.n732 0.13
R29949 VSS.n798 VSS.n733 0.13
R29950 VSS.n789 VSS.n788 0.13
R29951 VSS.n783 VSS.n782 0.13
R29952 VSS.n777 VSS.n776 0.13
R29953 VSS.n771 VSS.n770 0.13
R29954 VSS.n765 VSS.n764 0.13
R29955 VSS.n760 VSS.n759 0.13
R29956 VSS.n890 VSS.n822 0.13
R29957 VSS.n888 VSS.n823 0.13
R29958 VSS.n879 VSS.n878 0.13
R29959 VSS.n873 VSS.n872 0.13
R29960 VSS.n867 VSS.n866 0.13
R29961 VSS.n861 VSS.n860 0.13
R29962 VSS.n855 VSS.n854 0.13
R29963 VSS.n850 VSS.n849 0.13
R29964 VSS.n980 VSS.n912 0.13
R29965 VSS.n978 VSS.n913 0.13
R29966 VSS.n969 VSS.n968 0.13
R29967 VSS.n963 VSS.n962 0.13
R29968 VSS.n957 VSS.n956 0.13
R29969 VSS.n951 VSS.n950 0.13
R29970 VSS.n945 VSS.n944 0.13
R29971 VSS.n940 VSS.n939 0.13
R29972 VSS.n1070 VSS.n1002 0.13
R29973 VSS.n1068 VSS.n1003 0.13
R29974 VSS.n1059 VSS.n1058 0.13
R29975 VSS.n1053 VSS.n1052 0.13
R29976 VSS.n1047 VSS.n1046 0.13
R29977 VSS.n1041 VSS.n1040 0.13
R29978 VSS.n1035 VSS.n1034 0.13
R29979 VSS.n1030 VSS.n1029 0.13
R29980 VSS.n1160 VSS.n1092 0.13
R29981 VSS.n1158 VSS.n1093 0.13
R29982 VSS.n1149 VSS.n1148 0.13
R29983 VSS.n1143 VSS.n1142 0.13
R29984 VSS.n1137 VSS.n1136 0.13
R29985 VSS.n1131 VSS.n1130 0.13
R29986 VSS.n1125 VSS.n1124 0.13
R29987 VSS.n1120 VSS.n1119 0.13
R29988 VSS.n1245 VSS.n1182 0.13
R29989 VSS.n1243 VSS.n1183 0.13
R29990 VSS.n1234 VSS.n1233 0.13
R29991 VSS.n1228 VSS.n1227 0.13
R29992 VSS.n1222 VSS.n1221 0.13
R29993 VSS.n1216 VSS.n1215 0.13
R29994 VSS.n1210 VSS.n1209 0.13
R29995 VSS.n1205 VSS.n5 0.13
R29996 VSS.n10413 VSS.n10409 0.119
R29997 VSS.n13829 VSS.n10490 0.116
R29998 VSS.n17722 VSS.n0 0.116
R29999 VSS.n17553 VSS.n17549 0.115
R30000 VSS.n17556 VSS.n17509 0.115
R30001 VSS.n17559 VSS.n13989 0.115
R30002 VSS.n17562 VSS.n10396 0.115
R30003 VSS.n17565 VSS.n6631 0.115
R30004 VSS.n17568 VSS.n3108 0.115
R30005 VSS.n17571 VSS.n3081 0.115
R30006 VSS.n17576 VSS.n17575 0.115
R30007 VSS.n6900 sky130_asc_pnp_05v5_W3p40L3p40_1_0/VGND 0.11
R30008 VSS.n17573 VSS.n17572 0.106
R30009 VSS.n17570 VSS.n17569 0.106
R30010 VSS.n17567 VSS.n17566 0.106
R30011 VSS.n17564 VSS.n17563 0.106
R30012 VSS.n17561 VSS.n17560 0.106
R30013 VSS.n17558 VSS.n17557 0.106
R30014 VSS.n17555 VSS.n17554 0.106
R30015 VSS.n17552 VSS.n17551 0.106
R30016 VSS.n17714 VSS.n17713 0.106
R30017 VSS.n17715 VSS.n17714 0.106
R30018 VSS.n17716 VSS.n17715 0.106
R30019 VSS.n17717 VSS.n17716 0.106
R30020 VSS.n17718 VSS.n17717 0.106
R30021 VSS.n17719 VSS.n17718 0.106
R30022 VSS.n17720 VSS.n17719 0.106
R30023 VSS.n17721 VSS.n17720 0.106
R30024 VSS.n17722 VSS.n17721 0.106
R30025 VSS.n10414 VSS.n10413 0.106
R30026 VSS.t207 VSS.t184 0.101
R30027 VSS.t225 VSS.t167 0.101
R30028 VSS.t154 VSS.t206 0.101
R30029 VSS.t146 VSS.t153 0.101
R30030 VSS.t123 VSS.t175 0.101
R30031 VSS.t110 VSS.t122 0.101
R30032 VSS.t191 VSS.t135 0.101
R30033 VSS.t108 VSS.t163 0.101
R30034 VSS.t102 VSS.t112 0.101
R30035 VSS.t95 VSS.t213 0.101
R30036 VSS.t133 VSS.t179 0.101
R30037 VSS.t116 VSS.t157 0.101
R30038 VSS.t156 VSS.t200 0.101
R30039 VSS.t105 VSS.t150 0.101
R30040 VSS.t125 VSS.t170 0.101
R30041 VSS.t220 VSS.t115 0.101
R30042 VSS.t228 VSS.t129 0.101
R30043 VSS.t114 VSS.t155 0.101
R30044 VSS.t215 VSS.t104 0.101
R30045 VSS.t171 VSS.t210 0.101
R30046 VSS.t136 VSS.t183 0.101
R30047 VSS.t120 VSS.t161 0.101
R30048 VSS.t160 VSS.t203 0.101
R30049 VSS.t109 VSS.t152 0.101
R30050 VSS.t128 VSS.t173 0.101
R30051 VSS.t221 VSS.t118 0.101
R30052 VSS.t231 VSS.t131 0.101
R30053 VSS.t117 VSS.t159 0.101
R30054 VSS.t217 VSS.t107 0.101
R30055 VSS.t174 VSS.t212 0.101
R30056 VSS.n13513 VSS.n13512 0.101
R30057 VSS.t229 VSS.t196 0.101
R30058 VSS.t106 VSS.t218 0.101
R30059 VSS.t121 VSS.t226 0.101
R30060 VSS.t232 VSS.t198 0.101
R30061 VSS.t189 VSS.t149 0.101
R30062 VSS.t201 VSS.t168 0.101
R30063 VSS.t151 VSS.t113 0.101
R30064 VSS.t103 VSS.t214 0.101
R30065 VSS.t137 VSS.t98 0.101
R30066 VSS.t139 VSS.t99 0.101
R30067 VSS.t178 VSS.t216 0.101
R30068 VSS.t190 VSS.t223 0.101
R30069 VSS.t140 VSS.t185 0.101
R30070 VSS.t148 VSS.t192 0.101
R30071 VSS.t164 VSS.t205 0.101
R30072 VSS.t132 VSS.t177 0.101
R30073 VSS.t134 VSS.t181 0.101
R30074 VSS.t224 VSS.t126 0.101
R30075 VSS.t97 VSS.t142 0.101
R30076 VSS.t195 VSS.t94 0.101
R30077 VSS.n8929 VSS.n6901 0.1
R30078 VSS.n16023 VSS.n16022 0.098
R30079 VSS.n17464 VSS.n17463 0.096
R30080 VSS.n5663 VSS.n5662 0.091
R30081 VSS.n17703 VSS.n17641 0.089
R30082 VSS.n3135 sky130_asc_cap_mim_m3_1_9/VGND 0.081
R30083 VSS.n10413 VSS.n10412 0.077
R30084 VSS.n13457 VSS.n13456 0.073
R30085 VSS.n10371 VSS.n8930 0.071
R30086 VSS.n3131 VSS.n3130 0.071
R30087 VSS.n15999 sky130_asc_pnp_05v5_W3p40L3p40_8_3/Collector 0.066
R30088 VSS.n17333 sky130_asc_pnp_05v5_W3p40L3p40_8_3/Base 0.066
R30089 VSS.n12214 sky130_asc_pnp_05v5_W3p40L3p40_8_0/Collector 0.066
R30090 VSS.n13833 sky130_asc_pnp_05v5_W3p40L3p40_8_0/Base 0.066
R30091 VSS.n7177 sky130_asc_pnp_05v5_W3p40L3p40_8_1/Collector 0.066
R30092 VSS.n9097 sky130_asc_pnp_05v5_W3p40L3p40_8_1/Base 0.066
R30093 VSS.n3647 sky130_asc_pnp_05v5_W3p40L3p40_8_2/Collector 0.066
R30094 VSS.n3047 VSS.n3046 0.061
R30095 VSS.n6894 VSS.n6893 0.059
R30096 VSS.n10371 VSS.n10370 0.058
R30097 VSS.n13457 VSS.n11429 0.057
R30098 VSS.n17466 VSS.n17465 0.056
R30099 VSS.n3046 sky130_asc_pnp_05v5_W3p40L3p40_7_0/Collector 0.052
R30100 VSS.n6897 VSS.n6895 0.05
R30101 VSS.n3051 VSS.n1 0.047
R30102 VSS.n17520 sky130_asc_cap_mim_m3_1_8/Cout 0.047
R30103 VSS.n17476 sky130_asc_cap_mim_m3_1_6/Cout 0.047
R30104 VSS.n10410 sky130_asc_cap_mim_m3_1_7/Cout 0.047
R30105 VSS.n6892 sky130_asc_cap_mim_m3_1_5/Cout 0.047
R30106 VSS.n2873 VSS.n1266 0.046
R30107 VSS.n5664 sky130_asc_pnp_05v5_W3p40L3p40_8_2/Base 0.042
R30108 VSS.n10445 VSS.n10442 0.04
R30109 VSS.n10470 VSS.n10425 0.04
R30110 VSS.n17676 VSS.n17675 0.04
R30111 VSS.n17683 VSS.n17647 0.04
R30112 VSS.n5663 VSS.n3635 0.039
R30113 VSS.n17550 sky130_asc_res_xhigh_po_2p85_2_1/VGND 0.039
R30114 VSS.n10450 VSS.n10441 0.035
R30115 VSS.n10475 VSS.n10423 0.035
R30116 VSS.n17669 VSS.n17652 0.035
R30117 VSS.n17690 VSS.n17689 0.035
R30118 VSS.n16023 VSS.n13995 0.032
R30119 VSS.n17464 VSS.n16024 0.03
R30120 VSS.n8929 VSS.n8928 0.03
R30121 VSS.n0 VSS 0.03
R30122 VSS.n10455 VSS.n10440 0.029
R30123 VSS.n10480 VSS.n10421 0.029
R30124 VSS.n17664 VSS.n17654 0.029
R30125 VSS.n17697 VSS.n17644 0.029
R30126 VSS.n13514 VSS.n13513 0.028
R30127 VSS.n17708 VSS.n17707 0.026
R30128 VSS.n17579 VSS.n17578 0.025
R30129 VSS.n3079 VSS.n3078 0.025
R30130 VSS.n3106 VSS.n3105 0.025
R30131 VSS.n6629 VSS.n6628 0.025
R30132 VSS.n10394 VSS.n10393 0.025
R30133 VSS.n13987 VSS.n13986 0.025
R30134 VSS.n17507 VSS.n17506 0.025
R30135 VSS.n17547 VSS.n17546 0.025
R30136 VSS.n17545 VSS.n17544 0.025
R30137 VSS.n17505 VSS.n17504 0.025
R30138 VSS.n13985 VSS.n13984 0.025
R30139 VSS.n10392 VSS.n10391 0.025
R30140 VSS.n6627 VSS.n6626 0.025
R30141 VSS.n3104 VSS.n3103 0.025
R30142 VSS.n3077 VSS.n3076 0.025
R30143 VSS.n17581 VSS.n17580 0.025
R30144 VSS.n17710 VSS.n17709 0.025
R30145 VSS.n17613 VSS.n17612 0.025
R30146 VSS.n17615 VSS.n17614 0.025
R30147 VSS.n17628 VSS.n17627 0.025
R30148 VSS.n6898 VSS.n6883 0.025
R30149 VSS.n10459 VSS.n10458 0.024
R30150 VSS.n10485 VSS.n10419 0.024
R30151 VSS.n17659 VSS.n17656 0.024
R30152 VSS.n17699 VSS.n17641 0.024
R30153 VSS.n17521 VSS.t207 0.023
R30154 VSS.n17522 VSS.t225 0.023
R30155 VSS.n17523 VSS.n17522 0.023
R30156 VSS.n17513 VSS.t146 0.023
R30157 VSS.n17514 VSS.t123 0.023
R30158 VSS.n17515 VSS.t110 0.023
R30159 VSS.n17516 VSS.t191 0.023
R30160 VSS.n17517 VSS.t108 0.023
R30161 VSS.n17518 VSS.t102 0.023
R30162 VSS.n17519 VSS.t95 0.023
R30163 VSS.n17477 VSS.t133 0.023
R30164 VSS.n17478 VSS.t116 0.023
R30165 VSS.n17479 VSS.n17478 0.023
R30166 VSS.n17469 VSS.t105 0.023
R30167 VSS.n17470 VSS.t125 0.023
R30168 VSS.n17471 VSS.t220 0.023
R30169 VSS.n17472 VSS.t228 0.023
R30170 VSS.n17473 VSS.t114 0.023
R30171 VSS.n17474 VSS.t215 0.023
R30172 VSS.n17475 VSS.t171 0.023
R30173 VSS.n10411 VSS.t136 0.023
R30174 VSS.n10412 VSS.t120 0.023
R30175 VSS.n10403 VSS.t109 0.023
R30176 VSS.n10404 VSS.t128 0.023
R30177 VSS.n10405 VSS.t221 0.023
R30178 VSS.n10406 VSS.t231 0.023
R30179 VSS.n10407 VSS.t117 0.023
R30180 VSS.n10408 VSS.t217 0.023
R30181 VSS.n10409 VSS.t174 0.023
R30182 VSS.n6893 VSS.t229 0.023
R30183 VSS.n6884 VSS.t121 0.023
R30184 VSS.n6885 VSS.t232 0.023
R30185 VSS.n6886 VSS.t189 0.023
R30186 VSS.n6887 VSS.t201 0.023
R30187 VSS.n6888 VSS.t151 0.023
R30188 VSS.n6889 VSS.t103 0.023
R30189 VSS.n6890 VSS.t137 0.023
R30190 VSS.n6891 VSS.t139 0.023
R30191 VSS.n3115 VSS.t190 0.023
R30192 VSS.n3116 VSS.t140 0.023
R30193 VSS.n3117 VSS.t148 0.023
R30194 VSS.n3118 VSS.t164 0.023
R30195 VSS.n3119 VSS.t132 0.023
R30196 VSS.n3120 VSS.t134 0.023
R30197 VSS.n3121 VSS.t224 0.023
R30198 VSS.n3122 VSS.t97 0.023
R30199 VSS.n3123 VSS.t195 0.023
R30200 VSS.n5665 VSS.n5664 0.023
R30201 VSS.n17597 VSS.n17596 0.023
R30202 VSS.n3061 VSS.n3060 0.023
R30203 VSS.n3088 VSS.n3087 0.023
R30204 VSS.n6611 VSS.n6610 0.023
R30205 VSS.n10376 VSS.n10375 0.023
R30206 VSS.n13969 VSS.n13968 0.023
R30207 VSS.n17489 VSS.n17488 0.023
R30208 VSS.n17529 VSS.n17528 0.023
R30209 VSS.n17531 VSS.n17512 0.021
R30210 VSS.n17491 VSS.n13992 0.021
R30211 VSS.n13971 VSS.n10399 0.021
R30212 VSS.n10378 VSS.n6634 0.021
R30213 VSS.n6613 VSS.n3111 0.021
R30214 VSS.n3090 VSS.n3084 0.021
R30215 VSS.n3063 VSS.n3057 0.021
R30216 VSS.n17594 VSS.n3052 0.021
R30217 VSS.n17620 VSS.n17619 0.021
R30218 VSS.n17615 VSS.n17610 0.021
R30219 VSS.n17710 VSS.n17640 0.021
R30220 VSS.n17607 VSS.n17606 0.021
R30221 VSS.n17602 VSS.n17601 0.021
R30222 VSS.n17482 VSS.n17468 0.021
R30223 VSS.n10458 VSS.n10457 0.021
R30224 VSS.n10481 VSS.n10419 0.021
R30225 VSS.n3050 VSS.n1265 0.021
R30226 VSS.n17663 VSS.n17656 0.021
R30227 VSS.n17699 VSS.n17698 0.021
R30228 VSS.n17521 VSS.n17520 0.02
R30229 VSS.n17477 VSS.n17476 0.02
R30230 VSS.n10411 VSS.n10410 0.02
R30231 VSS.n6893 VSS.n6892 0.02
R30232 VSS.n17531 VSS.n17530 0.02
R30233 VSS.n17491 VSS.n17490 0.02
R30234 VSS.n13971 VSS.n13970 0.02
R30235 VSS.n10378 VSS.n10377 0.02
R30236 VSS.n6613 VSS.n6612 0.02
R30237 VSS.n3090 VSS.n3089 0.02
R30238 VSS.n3063 VSS.n3062 0.02
R30239 VSS.n17595 VSS.n17594 0.02
R30240 VSS.n3124 VSS.n3123 0.02
R30241 VSS.n17577 VSS.n17576 0.019
R30242 VSS.n3081 VSS.n3080 0.019
R30243 VSS.n3108 VSS.n3107 0.019
R30244 VSS.n6631 VSS.n6630 0.019
R30245 VSS.n10396 VSS.n10395 0.019
R30246 VSS.n13989 VSS.n13988 0.019
R30247 VSS.n17509 VSS.n17508 0.019
R30248 VSS.n17549 VSS.n17548 0.019
R30249 VSS.n17618 VSS.n17617 0.019
R30250 VSS.n17623 VSS.n17622 0.019
R30251 VSS.n17607 VSS.n17605 0.019
R30252 VSS.n3132 VSS.n3112 0.019
R30253 VSS.n3047 VSS.n1266 0.019
R30254 sky130_asc_res_xhigh_po_2p85_1_0/Rout VSS.n6606 0.018
R30255 VSS.n14375 VSS.n14369 0.017
R30256 VSS.n14712 VSS.n14711 0.017
R30257 VSS.n14700 VSS.n14378 0.017
R30258 VSS.n14698 VSS.n14384 0.017
R30259 VSS.n14689 VSS.n14688 0.017
R30260 VSS.n14677 VSS.n14397 0.017
R30261 VSS.n14675 VSS.n14403 0.017
R30262 VSS.n14667 VSS.n14666 0.017
R30263 VSS.n14655 VSS.n14416 0.017
R30264 VSS.n14653 VSS.n14422 0.017
R30265 VSS.n14644 VSS.n14643 0.017
R30266 VSS.n14632 VSS.n14435 0.017
R30267 VSS.n14629 VSS.n14475 0.017
R30268 VSS.n14620 VSS.n14619 0.017
R30269 VSS.n14608 VSS.n14490 0.017
R30270 VSS.n14606 VSS.n14496 0.017
R30271 VSS.n14597 VSS.n14596 0.017
R30272 VSS.n14585 VSS.n14509 0.017
R30273 VSS.n14583 VSS.n14515 0.017
R30274 VSS.n14575 VSS.n14574 0.017
R30275 VSS.n14563 VSS.n14528 0.017
R30276 VSS.n14561 VSS.n14534 0.017
R30277 VSS.n14552 VSS.n14551 0.017
R30278 VSS.n14869 VSS.n14868 0.017
R30279 VSS.n14880 VSS.n14879 0.017
R30280 VSS.n14293 VSS.n14291 0.017
R30281 VSS.n14893 VSS.n14285 0.017
R30282 VSS.n14905 VSS.n14904 0.017
R30283 VSS.n14915 VSS.n14914 0.017
R30284 VSS.n14272 VSS.n14270 0.017
R30285 VSS.n14928 VSS.n14264 0.017
R30286 VSS.n14939 VSS.n14938 0.017
R30287 VSS.n14949 VSS.n14948 0.017
R30288 VSS.n14251 VSS.n14249 0.017
R30289 VSS.n14962 VSS.n14243 0.017
R30290 VSS.n15327 VSS.n15326 0.017
R30291 VSS.n15322 VSS.n14973 0.017
R30292 VSS.n15313 VSS.n15312 0.017
R30293 VSS.n15301 VSS.n14987 0.017
R30294 VSS.n15299 VSS.n14993 0.017
R30295 VSS.n15290 VSS.n15289 0.017
R30296 VSS.n15278 VSS.n15006 0.017
R30297 VSS.n15276 VSS.n15012 0.017
R30298 VSS.n15268 VSS.n15267 0.017
R30299 VSS.n15256 VSS.n15025 0.017
R30300 VSS.n15254 VSS.n15031 0.017
R30301 VSS.n15245 VSS.n15244 0.017
R30302 VSS.n15233 VSS.n15044 0.017
R30303 VSS.n15230 VSS.n15084 0.017
R30304 VSS.n15221 VSS.n15220 0.017
R30305 VSS.n15209 VSS.n15099 0.017
R30306 VSS.n15207 VSS.n15105 0.017
R30307 VSS.n15198 VSS.n15197 0.017
R30308 VSS.n15186 VSS.n15118 0.017
R30309 VSS.n15184 VSS.n15124 0.017
R30310 VSS.n15176 VSS.n15175 0.017
R30311 VSS.n15164 VSS.n15137 0.017
R30312 VSS.n15162 VSS.n15143 0.017
R30313 VSS.n15153 VSS.n14138 0.017
R30314 VSS.n15451 VSS.n15450 0.017
R30315 VSS.n15456 VSS.n14129 0.017
R30316 VSS.n15468 VSS.n15467 0.017
R30317 VSS.n15478 VSS.n15477 0.017
R30318 VSS.n14116 VSS.n14114 0.017
R30319 VSS.n15491 VSS.n14108 0.017
R30320 VSS.n15503 VSS.n15502 0.017
R30321 VSS.n15512 VSS.n15511 0.017
R30322 VSS.n14095 VSS.n14093 0.017
R30323 VSS.n15525 VSS.n14087 0.017
R30324 VSS.n15537 VSS.n15536 0.017
R30325 VSS.n15547 VSS.n15546 0.017
R30326 VSS.n15558 VSS.n14073 0.017
R30327 VSS.n15889 VSS.n15560 0.017
R30328 VSS.n15880 VSS.n15879 0.017
R30329 VSS.n15868 VSS.n15574 0.017
R30330 VSS.n15866 VSS.n15580 0.017
R30331 VSS.n15857 VSS.n15856 0.017
R30332 VSS.n15845 VSS.n15593 0.017
R30333 VSS.n15843 VSS.n15599 0.017
R30334 VSS.n15835 VSS.n15834 0.017
R30335 VSS.n15823 VSS.n15612 0.017
R30336 VSS.n15821 VSS.n15618 0.017
R30337 VSS.n15812 VSS.n15811 0.017
R30338 VSS.n15800 VSS.n15631 0.017
R30339 VSS.n15797 VSS.n15671 0.017
R30340 VSS.n15788 VSS.n15787 0.017
R30341 VSS.n15776 VSS.n15686 0.017
R30342 VSS.n15774 VSS.n15692 0.017
R30343 VSS.n15765 VSS.n15764 0.017
R30344 VSS.n15753 VSS.n15705 0.017
R30345 VSS.n15751 VSS.n15711 0.017
R30346 VSS.n15743 VSS.n15742 0.017
R30347 VSS.n15731 VSS.n15724 0.017
R30348 VSS.n16022 VSS.n13996 0.017
R30349 VSS.n16013 VSS.n16012 0.017
R30350 VSS.n16001 VSS.n14008 0.017
R30351 VSS.n16688 VSS.n16633 0.017
R30352 VSS.n16757 VSS.n16756 0.017
R30353 VSS.n16747 VSS.n16690 0.017
R30354 VSS.n16745 VSS.n16692 0.017
R30355 VSS.n16739 VSS.n16698 0.017
R30356 VSS.n16733 VSS.n16702 0.017
R30357 VSS.n16727 VSS.n16706 0.017
R30358 VSS.n16721 VSS.n16709 0.017
R30359 VSS.n16716 VSS.n16712 0.017
R30360 VSS.n16778 VSS.n16543 0.017
R30361 VSS.n16847 VSS.n16846 0.017
R30362 VSS.n16837 VSS.n16780 0.017
R30363 VSS.n16835 VSS.n16782 0.017
R30364 VSS.n16829 VSS.n16788 0.017
R30365 VSS.n16823 VSS.n16792 0.017
R30366 VSS.n16817 VSS.n16796 0.017
R30367 VSS.n16811 VSS.n16799 0.017
R30368 VSS.n16806 VSS.n16802 0.017
R30369 VSS.n16868 VSS.n16453 0.017
R30370 VSS.n16937 VSS.n16936 0.017
R30371 VSS.n16927 VSS.n16870 0.017
R30372 VSS.n16925 VSS.n16872 0.017
R30373 VSS.n16919 VSS.n16878 0.017
R30374 VSS.n16913 VSS.n16882 0.017
R30375 VSS.n16907 VSS.n16886 0.017
R30376 VSS.n16901 VSS.n16889 0.017
R30377 VSS.n16896 VSS.n16892 0.017
R30378 VSS.n16958 VSS.n16363 0.017
R30379 VSS.n17027 VSS.n17026 0.017
R30380 VSS.n17017 VSS.n16960 0.017
R30381 VSS.n17015 VSS.n16962 0.017
R30382 VSS.n17009 VSS.n16968 0.017
R30383 VSS.n17003 VSS.n16972 0.017
R30384 VSS.n16997 VSS.n16976 0.017
R30385 VSS.n16991 VSS.n16979 0.017
R30386 VSS.n16986 VSS.n16982 0.017
R30387 VSS.n17048 VSS.n16273 0.017
R30388 VSS.n17117 VSS.n17116 0.017
R30389 VSS.n17107 VSS.n17050 0.017
R30390 VSS.n17105 VSS.n17052 0.017
R30391 VSS.n17099 VSS.n17058 0.017
R30392 VSS.n17093 VSS.n17062 0.017
R30393 VSS.n17087 VSS.n17066 0.017
R30394 VSS.n17081 VSS.n17069 0.017
R30395 VSS.n17076 VSS.n17072 0.017
R30396 VSS.n17138 VSS.n16183 0.017
R30397 VSS.n17207 VSS.n17206 0.017
R30398 VSS.n17197 VSS.n17140 0.017
R30399 VSS.n17195 VSS.n17142 0.017
R30400 VSS.n17189 VSS.n17148 0.017
R30401 VSS.n17183 VSS.n17152 0.017
R30402 VSS.n17177 VSS.n17156 0.017
R30403 VSS.n17171 VSS.n17159 0.017
R30404 VSS.n17166 VSS.n17162 0.017
R30405 VSS.n17228 VSS.n16093 0.017
R30406 VSS.n17297 VSS.n17296 0.017
R30407 VSS.n17287 VSS.n17230 0.017
R30408 VSS.n17285 VSS.n17232 0.017
R30409 VSS.n17279 VSS.n17238 0.017
R30410 VSS.n17273 VSS.n17242 0.017
R30411 VSS.n17267 VSS.n17246 0.017
R30412 VSS.n17261 VSS.n17249 0.017
R30413 VSS.n17256 VSS.n17252 0.017
R30414 VSS.n17389 VSS.n17388 0.017
R30415 VSS.n17397 VSS.n16050 0.017
R30416 VSS.n17453 VSS.n17452 0.017
R30417 VSS.n17443 VSS.n17399 0.017
R30418 VSS.n17441 VSS.n17401 0.017
R30419 VSS.n17435 VSS.n17407 0.017
R30420 VSS.n17429 VSS.n17411 0.017
R30421 VSS.n17423 VSS.n16025 0.017
R30422 VSS.n17463 VSS.n16026 0.017
R30423 VSS.n12720 VSS.n12718 0.017
R30424 VSS.n12803 VSS.n12712 0.017
R30425 VSS.n12815 VSS.n12814 0.017
R30426 VSS.n12825 VSS.n12824 0.017
R30427 VSS.n12699 VSS.n12697 0.017
R30428 VSS.n12838 VSS.n12691 0.017
R30429 VSS.n12850 VSS.n12849 0.017
R30430 VSS.n12859 VSS.n12858 0.017
R30431 VSS.n12678 VSS.n12676 0.017
R30432 VSS.n12872 VSS.n12668 0.017
R30433 VSS.n12885 VSS.n12884 0.017
R30434 VSS.n13062 VSS.n13061 0.017
R30435 VSS.n13051 VSS.n13050 0.017
R30436 VSS.n13039 VSS.n12895 0.017
R30437 VSS.n13037 VSS.n12902 0.017
R30438 VSS.n13028 VSS.n13027 0.017
R30439 VSS.n13016 VSS.n12915 0.017
R30440 VSS.n13014 VSS.n12921 0.017
R30441 VSS.n13006 VSS.n13005 0.017
R30442 VSS.n12994 VSS.n12934 0.017
R30443 VSS.n12992 VSS.n12940 0.017
R30444 VSS.n12983 VSS.n12982 0.017
R30445 VSS.n12971 VSS.n12953 0.017
R30446 VSS.n12969 VSS.n12960 0.017
R30447 VSS.n12579 VSS.n12577 0.017
R30448 VSS.n13160 VSS.n12571 0.017
R30449 VSS.n13172 VSS.n13171 0.017
R30450 VSS.n13182 VSS.n13181 0.017
R30451 VSS.n12558 VSS.n12556 0.017
R30452 VSS.n13195 VSS.n12550 0.017
R30453 VSS.n13207 VSS.n13206 0.017
R30454 VSS.n13216 VSS.n13215 0.017
R30455 VSS.n12537 VSS.n12535 0.017
R30456 VSS.n13229 VSS.n12527 0.017
R30457 VSS.n13242 VSS.n13241 0.017
R30458 VSS.n13311 VSS.n13310 0.017
R30459 VSS.n13300 VSS.n13299 0.017
R30460 VSS.n13288 VSS.n13252 0.017
R30461 VSS.n13286 VSS.n13259 0.017
R30462 VSS.n13277 VSS.n13276 0.017
R30463 VSS.n13456 VSS.n11430 0.017
R30464 VSS.n13447 VSS.n13446 0.017
R30465 VSS.n13436 VSS.n11442 0.017
R30466 VSS.n13434 VSS.n11448 0.017
R30467 VSS.n13425 VSS.n13424 0.017
R30468 VSS.n13413 VSS.n11461 0.017
R30469 VSS.n13411 VSS.n11467 0.017
R30470 VSS.n13402 VSS.n13401 0.017
R30471 VSS.n11670 VSS.n11668 0.017
R30472 VSS.n11681 VSS.n11662 0.017
R30473 VSS.n11693 VSS.n11692 0.017
R30474 VSS.n11703 VSS.n11702 0.017
R30475 VSS.n11649 VSS.n11647 0.017
R30476 VSS.n11716 VSS.n11641 0.017
R30477 VSS.n11728 VSS.n11727 0.017
R30478 VSS.n11737 VSS.n11736 0.017
R30479 VSS.n11628 VSS.n11626 0.017
R30480 VSS.n11750 VSS.n11620 0.017
R30481 VSS.n11762 VSS.n11761 0.017
R30482 VSS.n11772 VSS.n11771 0.017
R30483 VSS.n11814 VSS.n11813 0.017
R30484 VSS.n11598 VSS.n11596 0.017
R30485 VSS.n11827 VSS.n11590 0.017
R30486 VSS.n11839 VSS.n11838 0.017
R30487 VSS.n11849 VSS.n11848 0.017
R30488 VSS.n11577 VSS.n11575 0.017
R30489 VSS.n11862 VSS.n11569 0.017
R30490 VSS.n11873 VSS.n11872 0.017
R30491 VSS.n11883 VSS.n11882 0.017
R30492 VSS.n11556 VSS.n11554 0.017
R30493 VSS.n11896 VSS.n11548 0.017
R30494 VSS.n12402 VSS.n12401 0.017
R30495 VSS.n12397 VSS.n11907 0.017
R30496 VSS.n12388 VSS.n12387 0.017
R30497 VSS.n12376 VSS.n11921 0.017
R30498 VSS.n12374 VSS.n11927 0.017
R30499 VSS.n12365 VSS.n12364 0.017
R30500 VSS.n12353 VSS.n11940 0.017
R30501 VSS.n12351 VSS.n11946 0.017
R30502 VSS.n12343 VSS.n12342 0.017
R30503 VSS.n12331 VSS.n11959 0.017
R30504 VSS.n12329 VSS.n11965 0.017
R30505 VSS.n12320 VSS.n12319 0.017
R30506 VSS.n12308 VSS.n11978 0.017
R30507 VSS.n12305 VSS.n11985 0.017
R30508 VSS.n12296 VSS.n12295 0.017
R30509 VSS.n12284 VSS.n12000 0.017
R30510 VSS.n12282 VSS.n12006 0.017
R30511 VSS.n12273 VSS.n12272 0.017
R30512 VSS.n12261 VSS.n12019 0.017
R30513 VSS.n12259 VSS.n12025 0.017
R30514 VSS.n12251 VSS.n12250 0.017
R30515 VSS.n12239 VSS.n12038 0.017
R30516 VSS.n12237 VSS.n12044 0.017
R30517 VSS.n12228 VSS.n12227 0.017
R30518 VSS.n12216 VSS.n12057 0.017
R30519 VSS.n11155 VSS.n11100 0.017
R30520 VSS.n11225 VSS.n11224 0.017
R30521 VSS.n11215 VSS.n11157 0.017
R30522 VSS.n11213 VSS.n11159 0.017
R30523 VSS.n11207 VSS.n11165 0.017
R30524 VSS.n11201 VSS.n11169 0.017
R30525 VSS.n11195 VSS.n11172 0.017
R30526 VSS.n11190 VSS.n11175 0.017
R30527 VSS.n11184 VSS.n11178 0.017
R30528 VSS.n11245 VSS.n11010 0.017
R30529 VSS.n11315 VSS.n11314 0.017
R30530 VSS.n11305 VSS.n11247 0.017
R30531 VSS.n11303 VSS.n11249 0.017
R30532 VSS.n11297 VSS.n11255 0.017
R30533 VSS.n11291 VSS.n11259 0.017
R30534 VSS.n11285 VSS.n11262 0.017
R30535 VSS.n11280 VSS.n11265 0.017
R30536 VSS.n11274 VSS.n11268 0.017
R30537 VSS.n11335 VSS.n10920 0.017
R30538 VSS.n11405 VSS.n11404 0.017
R30539 VSS.n11395 VSS.n11337 0.017
R30540 VSS.n11393 VSS.n11339 0.017
R30541 VSS.n11387 VSS.n11345 0.017
R30542 VSS.n11381 VSS.n11349 0.017
R30543 VSS.n11375 VSS.n11352 0.017
R30544 VSS.n11370 VSS.n11355 0.017
R30545 VSS.n11364 VSS.n11358 0.017
R30546 VSS.n11425 VSS.n10830 0.017
R30547 VSS.n13525 VSS.n13524 0.017
R30548 VSS.n13515 VSS.n11427 0.017
R30549 VSS.n13512 VSS.n13458 0.017
R30550 VSS.n13506 VSS.n13464 0.017
R30551 VSS.n13500 VSS.n13468 0.017
R30552 VSS.n13494 VSS.n13471 0.017
R30553 VSS.n13489 VSS.n13474 0.017
R30554 VSS.n13483 VSS.n13477 0.017
R30555 VSS.n13545 VSS.n10740 0.017
R30556 VSS.n13615 VSS.n13614 0.017
R30557 VSS.n13605 VSS.n13547 0.017
R30558 VSS.n13603 VSS.n13549 0.017
R30559 VSS.n13597 VSS.n13555 0.017
R30560 VSS.n13591 VSS.n13559 0.017
R30561 VSS.n13585 VSS.n13562 0.017
R30562 VSS.n13580 VSS.n13565 0.017
R30563 VSS.n13574 VSS.n13568 0.017
R30564 VSS.n13635 VSS.n10650 0.017
R30565 VSS.n13705 VSS.n13704 0.017
R30566 VSS.n13695 VSS.n13637 0.017
R30567 VSS.n13693 VSS.n13639 0.017
R30568 VSS.n13687 VSS.n13645 0.017
R30569 VSS.n13681 VSS.n13649 0.017
R30570 VSS.n13675 VSS.n13652 0.017
R30571 VSS.n13670 VSS.n13655 0.017
R30572 VSS.n13664 VSS.n13658 0.017
R30573 VSS.n13725 VSS.n10560 0.017
R30574 VSS.n13795 VSS.n13794 0.017
R30575 VSS.n13785 VSS.n13727 0.017
R30576 VSS.n13783 VSS.n13729 0.017
R30577 VSS.n13777 VSS.n13735 0.017
R30578 VSS.n13771 VSS.n13739 0.017
R30579 VSS.n13765 VSS.n13742 0.017
R30580 VSS.n13760 VSS.n13745 0.017
R30581 VSS.n13754 VSS.n13748 0.017
R30582 VSS.n13889 VSS.n13888 0.017
R30583 VSS.n13897 VSS.n10517 0.017
R30584 VSS.n13945 VSS.n13944 0.017
R30585 VSS.n13935 VSS.n13899 0.017
R30586 VSS.n13933 VSS.n13901 0.017
R30587 VSS.n13927 VSS.n13907 0.017
R30588 VSS.n13921 VSS.n13911 0.017
R30589 VSS.n13959 VSS.n10491 0.017
R30590 VSS.n13831 VSS.n13829 0.017
R30591 VSS.n7682 VSS.n7676 0.017
R30592 VSS.n7826 VSS.n7825 0.017
R30593 VSS.n7814 VSS.n7685 0.017
R30594 VSS.n7812 VSS.n7691 0.017
R30595 VSS.n7803 VSS.n7802 0.017
R30596 VSS.n7791 VSS.n7704 0.017
R30597 VSS.n7789 VSS.n7710 0.017
R30598 VSS.n7781 VSS.n7780 0.017
R30599 VSS.n7769 VSS.n7723 0.017
R30600 VSS.n7767 VSS.n7729 0.017
R30601 VSS.n7758 VSS.n7757 0.017
R30602 VSS.n7746 VSS.n7742 0.017
R30603 VSS.n7925 VSS.n7924 0.017
R30604 VSS.n7592 VSS.n7590 0.017
R30605 VSS.n7938 VSS.n7584 0.017
R30606 VSS.n7950 VSS.n7949 0.017
R30607 VSS.n7960 VSS.n7959 0.017
R30608 VSS.n7571 VSS.n7569 0.017
R30609 VSS.n7973 VSS.n7563 0.017
R30610 VSS.n7984 VSS.n7983 0.017
R30611 VSS.n7994 VSS.n7993 0.017
R30612 VSS.n7550 VSS.n7548 0.017
R30613 VSS.n8007 VSS.n7542 0.017
R30614 VSS.n8188 VSS.n8187 0.017
R30615 VSS.n8028 VSS.n8025 0.017
R30616 VSS.n8036 VSS.n8030 0.017
R30617 VSS.n8166 VSS.n8165 0.017
R30618 VSS.n8154 VSS.n8039 0.017
R30619 VSS.n8152 VSS.n8045 0.017
R30620 VSS.n8143 VSS.n8142 0.017
R30621 VSS.n8132 VSS.n8058 0.017
R30622 VSS.n8130 VSS.n8064 0.017
R30623 VSS.n8121 VSS.n8120 0.017
R30624 VSS.n8109 VSS.n8077 0.017
R30625 VSS.n8107 VSS.n8083 0.017
R30626 VSS.n8098 VSS.n8097 0.017
R30627 VSS.n8283 VSS.n8282 0.017
R30628 VSS.n7452 VSS.n7450 0.017
R30629 VSS.n8296 VSS.n7444 0.017
R30630 VSS.n8308 VSS.n8307 0.017
R30631 VSS.n8318 VSS.n8317 0.017
R30632 VSS.n7431 VSS.n7429 0.017
R30633 VSS.n8331 VSS.n7423 0.017
R30634 VSS.n8342 VSS.n8341 0.017
R30635 VSS.n8352 VSS.n8351 0.017
R30636 VSS.n7410 VSS.n7408 0.017
R30637 VSS.n8365 VSS.n7402 0.017
R30638 VSS.n8546 VSS.n8545 0.017
R30639 VSS.n8386 VSS.n8383 0.017
R30640 VSS.n8394 VSS.n8388 0.017
R30641 VSS.n8524 VSS.n8523 0.017
R30642 VSS.n8512 VSS.n8397 0.017
R30643 VSS.n8510 VSS.n8403 0.017
R30644 VSS.n8501 VSS.n8500 0.017
R30645 VSS.n8490 VSS.n8416 0.017
R30646 VSS.n8488 VSS.n8422 0.017
R30647 VSS.n8479 VSS.n8478 0.017
R30648 VSS.n8467 VSS.n8435 0.017
R30649 VSS.n8465 VSS.n8441 0.017
R30650 VSS.n8456 VSS.n8455 0.017
R30651 VSS.n8641 VSS.n8640 0.017
R30652 VSS.n7312 VSS.n7310 0.017
R30653 VSS.n8654 VSS.n7304 0.017
R30654 VSS.n8666 VSS.n8665 0.017
R30655 VSS.n8676 VSS.n8675 0.017
R30656 VSS.n7291 VSS.n7289 0.017
R30657 VSS.n8689 VSS.n7283 0.017
R30658 VSS.n8700 VSS.n8699 0.017
R30659 VSS.n8710 VSS.n8709 0.017
R30660 VSS.n7270 VSS.n7268 0.017
R30661 VSS.n8723 VSS.n7262 0.017
R30662 VSS.n8768 VSS.n8767 0.017
R30663 VSS.n8744 VSS.n8741 0.017
R30664 VSS.n8747 VSS.n8746 0.017
R30665 VSS.n8928 VSS.n6902 0.017
R30666 VSS.n8919 VSS.n8918 0.017
R30667 VSS.n8907 VSS.n6914 0.017
R30668 VSS.n8905 VSS.n6920 0.017
R30669 VSS.n8897 VSS.n8896 0.017
R30670 VSS.n8885 VSS.n6933 0.017
R30671 VSS.n8883 VSS.n6939 0.017
R30672 VSS.n8874 VSS.n8873 0.017
R30673 VSS.n8862 VSS.n6952 0.017
R30674 VSS.n8860 VSS.n6958 0.017
R30675 VSS.n7072 VSS.n7064 0.017
R30676 VSS.n7084 VSS.n7083 0.017
R30677 VSS.n7094 VSS.n7093 0.017
R30678 VSS.n7051 VSS.n7049 0.017
R30679 VSS.n7107 VSS.n7043 0.017
R30680 VSS.n7119 VSS.n7118 0.017
R30681 VSS.n7128 VSS.n7127 0.017
R30682 VSS.n7030 VSS.n7028 0.017
R30683 VSS.n7141 VSS.n7022 0.017
R30684 VSS.n7153 VSS.n7152 0.017
R30685 VSS.n7163 VSS.n7162 0.017
R30686 VSS.n7008 VSS.n7006 0.017
R30687 VSS.n9733 VSS.n9678 0.017
R30688 VSS.n9802 VSS.n9801 0.017
R30689 VSS.n9792 VSS.n9735 0.017
R30690 VSS.n9790 VSS.n9737 0.017
R30691 VSS.n9784 VSS.n9743 0.017
R30692 VSS.n9778 VSS.n9747 0.017
R30693 VSS.n9772 VSS.n9751 0.017
R30694 VSS.n9766 VSS.n9754 0.017
R30695 VSS.n9761 VSS.n9757 0.017
R30696 VSS.n9823 VSS.n9588 0.017
R30697 VSS.n9892 VSS.n9891 0.017
R30698 VSS.n9882 VSS.n9825 0.017
R30699 VSS.n9880 VSS.n9827 0.017
R30700 VSS.n9874 VSS.n9833 0.017
R30701 VSS.n9868 VSS.n9837 0.017
R30702 VSS.n9862 VSS.n9841 0.017
R30703 VSS.n9856 VSS.n9844 0.017
R30704 VSS.n9851 VSS.n9847 0.017
R30705 VSS.n9913 VSS.n9498 0.017
R30706 VSS.n9982 VSS.n9981 0.017
R30707 VSS.n9972 VSS.n9915 0.017
R30708 VSS.n9970 VSS.n9917 0.017
R30709 VSS.n9964 VSS.n9923 0.017
R30710 VSS.n9958 VSS.n9927 0.017
R30711 VSS.n9952 VSS.n9931 0.017
R30712 VSS.n9946 VSS.n9934 0.017
R30713 VSS.n9941 VSS.n9937 0.017
R30714 VSS.n10003 VSS.n9408 0.017
R30715 VSS.n10072 VSS.n10071 0.017
R30716 VSS.n10062 VSS.n10005 0.017
R30717 VSS.n10060 VSS.n10007 0.017
R30718 VSS.n10054 VSS.n10013 0.017
R30719 VSS.n10048 VSS.n10017 0.017
R30720 VSS.n10042 VSS.n10021 0.017
R30721 VSS.n10036 VSS.n10024 0.017
R30722 VSS.n10031 VSS.n10027 0.017
R30723 VSS.n10093 VSS.n9318 0.017
R30724 VSS.n10162 VSS.n10161 0.017
R30725 VSS.n10152 VSS.n10095 0.017
R30726 VSS.n10150 VSS.n10097 0.017
R30727 VSS.n10144 VSS.n10103 0.017
R30728 VSS.n10138 VSS.n10107 0.017
R30729 VSS.n10132 VSS.n10111 0.017
R30730 VSS.n10126 VSS.n10114 0.017
R30731 VSS.n10121 VSS.n10117 0.017
R30732 VSS.n10183 VSS.n9228 0.017
R30733 VSS.n10252 VSS.n10251 0.017
R30734 VSS.n10242 VSS.n10185 0.017
R30735 VSS.n10240 VSS.n10187 0.017
R30736 VSS.n10234 VSS.n10193 0.017
R30737 VSS.n10228 VSS.n10197 0.017
R30738 VSS.n10222 VSS.n10201 0.017
R30739 VSS.n10216 VSS.n10204 0.017
R30740 VSS.n10211 VSS.n10207 0.017
R30741 VSS.n10320 VSS.n10319 0.017
R30742 VSS.n10370 VSS.n8931 0.017
R30743 VSS.n8944 VSS.n8940 0.017
R30744 VSS.n8950 VSS.n8946 0.017
R30745 VSS.n8955 VSS.n8952 0.017
R30746 VSS.n8962 VSS.n8957 0.017
R30747 VSS.n8968 VSS.n8964 0.017
R30748 VSS.n8974 VSS.n8970 0.017
R30749 VSS.n8979 VSS.n8976 0.017
R30750 VSS.n9033 VSS.n8981 0.017
R30751 VSS.n9041 VSS.n9031 0.017
R30752 VSS.n9049 VSS.n9029 0.017
R30753 VSS.n9057 VSS.n9027 0.017
R30754 VSS.n9065 VSS.n9025 0.017
R30755 VSS.n9073 VSS.n9023 0.017
R30756 VSS.n9081 VSS.n9021 0.017
R30757 VSS.n9089 VSS.n9019 0.017
R30758 VSS.n9152 VSS.n9151 0.017
R30759 VSS.n4173 VSS.n4171 0.017
R30760 VSS.n4256 VSS.n4165 0.017
R30761 VSS.n4268 VSS.n4267 0.017
R30762 VSS.n4278 VSS.n4277 0.017
R30763 VSS.n4152 VSS.n4150 0.017
R30764 VSS.n4291 VSS.n4144 0.017
R30765 VSS.n4303 VSS.n4302 0.017
R30766 VSS.n4312 VSS.n4311 0.017
R30767 VSS.n4131 VSS.n4129 0.017
R30768 VSS.n4325 VSS.n4121 0.017
R30769 VSS.n4338 VSS.n4337 0.017
R30770 VSS.n4515 VSS.n4514 0.017
R30771 VSS.n4504 VSS.n4503 0.017
R30772 VSS.n4492 VSS.n4348 0.017
R30773 VSS.n4490 VSS.n4355 0.017
R30774 VSS.n4481 VSS.n4480 0.017
R30775 VSS.n4469 VSS.n4368 0.017
R30776 VSS.n4467 VSS.n4374 0.017
R30777 VSS.n4459 VSS.n4458 0.017
R30778 VSS.n4447 VSS.n4387 0.017
R30779 VSS.n4445 VSS.n4393 0.017
R30780 VSS.n4436 VSS.n4435 0.017
R30781 VSS.n4424 VSS.n4406 0.017
R30782 VSS.n4422 VSS.n4413 0.017
R30783 VSS.n4032 VSS.n4030 0.017
R30784 VSS.n4613 VSS.n4024 0.017
R30785 VSS.n4625 VSS.n4624 0.017
R30786 VSS.n4635 VSS.n4634 0.017
R30787 VSS.n4011 VSS.n4009 0.017
R30788 VSS.n4648 VSS.n4003 0.017
R30789 VSS.n4660 VSS.n4659 0.017
R30790 VSS.n4669 VSS.n4668 0.017
R30791 VSS.n3990 VSS.n3988 0.017
R30792 VSS.n4682 VSS.n3980 0.017
R30793 VSS.n4695 VSS.n4694 0.017
R30794 VSS.n4872 VSS.n4871 0.017
R30795 VSS.n4861 VSS.n4860 0.017
R30796 VSS.n4849 VSS.n4705 0.017
R30797 VSS.n4847 VSS.n4712 0.017
R30798 VSS.n4838 VSS.n4837 0.017
R30799 VSS.n4826 VSS.n4725 0.017
R30800 VSS.n4824 VSS.n4731 0.017
R30801 VSS.n4816 VSS.n4815 0.017
R30802 VSS.n4804 VSS.n4744 0.017
R30803 VSS.n4802 VSS.n4750 0.017
R30804 VSS.n4793 VSS.n4792 0.017
R30805 VSS.n4781 VSS.n4763 0.017
R30806 VSS.n4779 VSS.n4770 0.017
R30807 VSS.n3891 VSS.n3889 0.017
R30808 VSS.n4970 VSS.n3883 0.017
R30809 VSS.n4982 VSS.n4981 0.017
R30810 VSS.n4992 VSS.n4991 0.017
R30811 VSS.n3870 VSS.n3868 0.017
R30812 VSS.n5005 VSS.n3862 0.017
R30813 VSS.n5017 VSS.n5016 0.017
R30814 VSS.n5026 VSS.n5025 0.017
R30815 VSS.n3849 VSS.n3847 0.017
R30816 VSS.n5039 VSS.n3839 0.017
R30817 VSS.n5052 VSS.n5051 0.017
R30818 VSS.n5229 VSS.n5228 0.017
R30819 VSS.n5218 VSS.n5217 0.017
R30820 VSS.n5206 VSS.n5062 0.017
R30821 VSS.n5204 VSS.n5069 0.017
R30822 VSS.n5195 VSS.n5194 0.017
R30823 VSS.n5183 VSS.n5082 0.017
R30824 VSS.n5181 VSS.n5088 0.017
R30825 VSS.n5173 VSS.n5172 0.017
R30826 VSS.n5161 VSS.n5101 0.017
R30827 VSS.n5159 VSS.n5107 0.017
R30828 VSS.n5150 VSS.n5149 0.017
R30829 VSS.n5138 VSS.n5120 0.017
R30830 VSS.n5136 VSS.n5127 0.017
R30831 VSS.n3750 VSS.n3748 0.017
R30832 VSS.n5327 VSS.n3742 0.017
R30833 VSS.n5339 VSS.n5338 0.017
R30834 VSS.n5349 VSS.n5348 0.017
R30835 VSS.n3729 VSS.n3727 0.017
R30836 VSS.n5362 VSS.n3721 0.017
R30837 VSS.n5374 VSS.n5373 0.017
R30838 VSS.n5383 VSS.n5382 0.017
R30839 VSS.n3708 VSS.n3706 0.017
R30840 VSS.n5396 VSS.n3698 0.017
R30841 VSS.n5409 VSS.n5408 0.017
R30842 VSS.n5575 VSS.n5574 0.017
R30843 VSS.n5564 VSS.n5563 0.017
R30844 VSS.n5552 VSS.n5419 0.017
R30845 VSS.n5550 VSS.n5426 0.017
R30846 VSS.n5541 VSS.n5540 0.017
R30847 VSS.n5529 VSS.n5439 0.017
R30848 VSS.n5527 VSS.n5445 0.017
R30849 VSS.n5519 VSS.n5518 0.017
R30850 VSS.n5507 VSS.n5458 0.017
R30851 VSS.n5505 VSS.n5464 0.017
R30852 VSS.n5496 VSS.n5495 0.017
R30853 VSS.n5484 VSS.n5477 0.017
R30854 VSS.n5662 VSS.n3636 0.017
R30855 VSS.n3174 VSS.n3173 0.017
R30856 VSS.n3181 VSS.n3171 0.017
R30857 VSS.n3189 VSS.n3169 0.017
R30858 VSS.n3197 VSS.n3167 0.017
R30859 VSS.n3205 VSS.n3165 0.017
R30860 VSS.n3213 VSS.n3163 0.017
R30861 VSS.n3221 VSS.n3161 0.017
R30862 VSS.n6594 VSS.n6593 0.017
R30863 VSS.n6517 VSS.n3230 0.017
R30864 VSS.n3243 VSS.n3239 0.017
R30865 VSS.n3249 VSS.n3245 0.017
R30866 VSS.n3255 VSS.n3251 0.017
R30867 VSS.n3260 VSS.n3257 0.017
R30868 VSS.n3267 VSS.n3262 0.017
R30869 VSS.n3273 VSS.n3269 0.017
R30870 VSS.n3279 VSS.n3275 0.017
R30871 VSS.n3285 VSS.n3281 0.017
R30872 VSS.n6395 VSS.n3288 0.017
R30873 VSS.n3301 VSS.n3297 0.017
R30874 VSS.n3307 VSS.n3303 0.017
R30875 VSS.n3313 VSS.n3309 0.017
R30876 VSS.n3318 VSS.n3315 0.017
R30877 VSS.n3325 VSS.n3320 0.017
R30878 VSS.n3331 VSS.n3327 0.017
R30879 VSS.n3337 VSS.n3333 0.017
R30880 VSS.n3343 VSS.n3339 0.017
R30881 VSS.n6273 VSS.n3346 0.017
R30882 VSS.n3359 VSS.n3355 0.017
R30883 VSS.n3365 VSS.n3361 0.017
R30884 VSS.n3371 VSS.n3367 0.017
R30885 VSS.n3376 VSS.n3373 0.017
R30886 VSS.n3383 VSS.n3378 0.017
R30887 VSS.n3389 VSS.n3385 0.017
R30888 VSS.n3395 VSS.n3391 0.017
R30889 VSS.n3401 VSS.n3397 0.017
R30890 VSS.n6151 VSS.n3404 0.017
R30891 VSS.n3417 VSS.n3413 0.017
R30892 VSS.n3423 VSS.n3419 0.017
R30893 VSS.n3429 VSS.n3425 0.017
R30894 VSS.n3434 VSS.n3431 0.017
R30895 VSS.n3441 VSS.n3436 0.017
R30896 VSS.n3447 VSS.n3443 0.017
R30897 VSS.n3453 VSS.n3449 0.017
R30898 VSS.n3459 VSS.n3455 0.017
R30899 VSS.n6029 VSS.n3462 0.017
R30900 VSS.n3475 VSS.n3471 0.017
R30901 VSS.n3481 VSS.n3477 0.017
R30902 VSS.n3487 VSS.n3483 0.017
R30903 VSS.n3492 VSS.n3489 0.017
R30904 VSS.n3499 VSS.n3494 0.017
R30905 VSS.n3505 VSS.n3501 0.017
R30906 VSS.n3511 VSS.n3507 0.017
R30907 VSS.n3517 VSS.n3513 0.017
R30908 VSS.n5907 VSS.n3520 0.017
R30909 VSS.n3533 VSS.n3529 0.017
R30910 VSS.n3539 VSS.n3535 0.017
R30911 VSS.n3545 VSS.n3541 0.017
R30912 VSS.n3550 VSS.n3547 0.017
R30913 VSS.n3557 VSS.n3552 0.017
R30914 VSS.n3563 VSS.n3559 0.017
R30915 VSS.n3569 VSS.n3565 0.017
R30916 VSS.n3575 VSS.n3571 0.017
R30917 VSS.n5785 VSS.n3578 0.017
R30918 VSS.n3591 VSS.n3587 0.017
R30919 VSS.n3597 VSS.n3593 0.017
R30920 VSS.n3603 VSS.n3599 0.017
R30921 VSS.n3608 VSS.n3605 0.017
R30922 VSS.n3615 VSS.n3610 0.017
R30923 VSS.n3621 VSS.n3617 0.017
R30924 VSS.n3627 VSS.n3623 0.017
R30925 VSS.n3633 VSS.n3629 0.017
R30926 VSS.n1616 VSS.n1610 0.017
R30927 VSS.n1953 VSS.n1952 0.017
R30928 VSS.n1941 VSS.n1619 0.017
R30929 VSS.n1939 VSS.n1625 0.017
R30930 VSS.n1930 VSS.n1929 0.017
R30931 VSS.n1918 VSS.n1638 0.017
R30932 VSS.n1916 VSS.n1644 0.017
R30933 VSS.n1908 VSS.n1907 0.017
R30934 VSS.n1896 VSS.n1657 0.017
R30935 VSS.n1894 VSS.n1663 0.017
R30936 VSS.n1885 VSS.n1884 0.017
R30937 VSS.n1873 VSS.n1676 0.017
R30938 VSS.n1870 VSS.n1716 0.017
R30939 VSS.n1861 VSS.n1860 0.017
R30940 VSS.n1849 VSS.n1731 0.017
R30941 VSS.n1847 VSS.n1737 0.017
R30942 VSS.n1838 VSS.n1837 0.017
R30943 VSS.n1826 VSS.n1750 0.017
R30944 VSS.n1824 VSS.n1756 0.017
R30945 VSS.n1816 VSS.n1815 0.017
R30946 VSS.n1804 VSS.n1769 0.017
R30947 VSS.n1802 VSS.n1775 0.017
R30948 VSS.n1793 VSS.n1792 0.017
R30949 VSS.n2110 VSS.n2109 0.017
R30950 VSS.n2121 VSS.n2120 0.017
R30951 VSS.n1534 VSS.n1532 0.017
R30952 VSS.n2134 VSS.n1526 0.017
R30953 VSS.n2146 VSS.n2145 0.017
R30954 VSS.n2156 VSS.n2155 0.017
R30955 VSS.n1513 VSS.n1511 0.017
R30956 VSS.n2169 VSS.n1505 0.017
R30957 VSS.n2180 VSS.n2179 0.017
R30958 VSS.n2190 VSS.n2189 0.017
R30959 VSS.n1492 VSS.n1490 0.017
R30960 VSS.n2203 VSS.n1484 0.017
R30961 VSS.n2568 VSS.n2567 0.017
R30962 VSS.n2563 VSS.n2214 0.017
R30963 VSS.n2554 VSS.n2553 0.017
R30964 VSS.n2542 VSS.n2228 0.017
R30965 VSS.n2540 VSS.n2234 0.017
R30966 VSS.n2531 VSS.n2530 0.017
R30967 VSS.n2519 VSS.n2247 0.017
R30968 VSS.n2517 VSS.n2253 0.017
R30969 VSS.n2509 VSS.n2508 0.017
R30970 VSS.n2497 VSS.n2266 0.017
R30971 VSS.n2495 VSS.n2272 0.017
R30972 VSS.n2486 VSS.n2485 0.017
R30973 VSS.n2474 VSS.n2285 0.017
R30974 VSS.n2471 VSS.n2325 0.017
R30975 VSS.n2462 VSS.n2461 0.017
R30976 VSS.n2450 VSS.n2340 0.017
R30977 VSS.n2448 VSS.n2346 0.017
R30978 VSS.n2439 VSS.n2438 0.017
R30979 VSS.n2427 VSS.n2359 0.017
R30980 VSS.n2425 VSS.n2365 0.017
R30981 VSS.n2417 VSS.n2416 0.017
R30982 VSS.n2405 VSS.n2378 0.017
R30983 VSS.n2403 VSS.n2384 0.017
R30984 VSS.n2394 VSS.n1379 0.017
R30985 VSS.n2692 VSS.n2691 0.017
R30986 VSS.n2697 VSS.n1370 0.017
R30987 VSS.n2709 VSS.n2708 0.017
R30988 VSS.n2719 VSS.n2718 0.017
R30989 VSS.n1357 VSS.n1355 0.017
R30990 VSS.n2732 VSS.n1349 0.017
R30991 VSS.n2744 VSS.n2743 0.017
R30992 VSS.n2753 VSS.n2752 0.017
R30993 VSS.n1336 VSS.n1334 0.017
R30994 VSS.n2766 VSS.n1328 0.017
R30995 VSS.n2778 VSS.n2777 0.017
R30996 VSS.n2788 VSS.n2787 0.017
R30997 VSS.n2799 VSS.n1314 0.017
R30998 VSS.n2963 VSS.n2801 0.017
R30999 VSS.n2954 VSS.n2953 0.017
R31000 VSS.n2942 VSS.n2815 0.017
R31001 VSS.n2940 VSS.n2821 0.017
R31002 VSS.n2931 VSS.n2930 0.017
R31003 VSS.n2919 VSS.n2834 0.017
R31004 VSS.n2917 VSS.n2840 0.017
R31005 VSS.n2909 VSS.n2908 0.017
R31006 VSS.n2897 VSS.n2853 0.017
R31007 VSS.n2895 VSS.n2859 0.017
R31008 VSS.n2886 VSS.n2885 0.017
R31009 VSS.n2874 VSS.n2872 0.017
R31010 VSS.n641 VSS.n586 0.017
R31011 VSS.n710 VSS.n709 0.017
R31012 VSS.n700 VSS.n643 0.017
R31013 VSS.n698 VSS.n645 0.017
R31014 VSS.n692 VSS.n651 0.017
R31015 VSS.n686 VSS.n655 0.017
R31016 VSS.n680 VSS.n659 0.017
R31017 VSS.n674 VSS.n662 0.017
R31018 VSS.n669 VSS.n665 0.017
R31019 VSS.n731 VSS.n496 0.017
R31020 VSS.n800 VSS.n799 0.017
R31021 VSS.n790 VSS.n733 0.017
R31022 VSS.n788 VSS.n735 0.017
R31023 VSS.n782 VSS.n741 0.017
R31024 VSS.n776 VSS.n745 0.017
R31025 VSS.n770 VSS.n749 0.017
R31026 VSS.n764 VSS.n752 0.017
R31027 VSS.n759 VSS.n755 0.017
R31028 VSS.n821 VSS.n406 0.017
R31029 VSS.n890 VSS.n889 0.017
R31030 VSS.n880 VSS.n823 0.017
R31031 VSS.n878 VSS.n825 0.017
R31032 VSS.n872 VSS.n831 0.017
R31033 VSS.n866 VSS.n835 0.017
R31034 VSS.n860 VSS.n839 0.017
R31035 VSS.n854 VSS.n842 0.017
R31036 VSS.n849 VSS.n845 0.017
R31037 VSS.n911 VSS.n316 0.017
R31038 VSS.n980 VSS.n979 0.017
R31039 VSS.n970 VSS.n913 0.017
R31040 VSS.n968 VSS.n915 0.017
R31041 VSS.n962 VSS.n921 0.017
R31042 VSS.n956 VSS.n925 0.017
R31043 VSS.n950 VSS.n929 0.017
R31044 VSS.n944 VSS.n932 0.017
R31045 VSS.n939 VSS.n935 0.017
R31046 VSS.n1001 VSS.n226 0.017
R31047 VSS.n1070 VSS.n1069 0.017
R31048 VSS.n1060 VSS.n1003 0.017
R31049 VSS.n1058 VSS.n1005 0.017
R31050 VSS.n1052 VSS.n1011 0.017
R31051 VSS.n1046 VSS.n1015 0.017
R31052 VSS.n1040 VSS.n1019 0.017
R31053 VSS.n1034 VSS.n1022 0.017
R31054 VSS.n1029 VSS.n1025 0.017
R31055 VSS.n1091 VSS.n136 0.017
R31056 VSS.n1160 VSS.n1159 0.017
R31057 VSS.n1150 VSS.n1093 0.017
R31058 VSS.n1148 VSS.n1095 0.017
R31059 VSS.n1142 VSS.n1101 0.017
R31060 VSS.n1136 VSS.n1105 0.017
R31061 VSS.n1130 VSS.n1109 0.017
R31062 VSS.n1124 VSS.n1112 0.017
R31063 VSS.n1119 VSS.n1115 0.017
R31064 VSS.n1181 VSS.n45 0.017
R31065 VSS.n1245 VSS.n1244 0.017
R31066 VSS.n1235 VSS.n1183 0.017
R31067 VSS.n1233 VSS.n1185 0.017
R31068 VSS.n1227 VSS.n1191 0.017
R31069 VSS.n1221 VSS.n1195 0.017
R31070 VSS.n1215 VSS.n1199 0.017
R31071 VSS.n1209 VSS.n1202 0.017
R31072 VSS.n1258 VSS.n5 0.017
R31073 VSS.n1264 VSS.n2 0.017
R31074 VSS.n10451 VSS.n10440 0.016
R31075 VSS.n10476 VSS.n10421 0.016
R31076 VSS.n6605 VSS.n6604 0.016
R31077 VSS.n17668 VSS.n17654 0.016
R31078 VSS.n17645 VSS.n17644 0.016
R31079 VSS.n3128 VSS.n3127 0.016
R31080 VSS.n17520 sky130_asc_cap_mim_m3_1_8/Cout 0.016
R31081 VSS.n17476 sky130_asc_cap_mim_m3_1_6/Cout 0.016
R31082 VSS.n10410 sky130_asc_cap_mim_m3_1_7/Cout 0.016
R31083 VSS.n6892 sky130_asc_cap_mim_m3_1_5/Cout 0.016
R31084 VSS.n3125 sky130_asc_cap_mim_m3_1_9/Cout 0.015
R31085 sky130_asc_pnp_05v5_W3p40L3p40_7_0/Base VSS.n3048 0.015
R31086 VSS.n17483 VSS.n17467 0.015
R31087 VSS.n17548 VSS.n17547 0.014
R31088 VSS.n17508 VSS.n17507 0.014
R31089 VSS.n13988 VSS.n13987 0.014
R31090 VSS.n10395 VSS.n10394 0.014
R31091 VSS.n6630 VSS.n6629 0.014
R31092 VSS.n3107 VSS.n3106 0.014
R31093 VSS.n3080 VSS.n3079 0.014
R31094 VSS.n17578 VSS.n17577 0.014
R31095 VSS.n17605 VSS.n17604 0.014
R31096 VSS.n17625 VSS.n17624 0.014
R31097 VSS.n17623 VSS.n17620 0.014
R31098 VSS.n17618 VSS.n17615 0.014
R31099 VSS.n3126 VSS.n3114 0.014
R31100 VSS.n3129 sky130_asc_cap_mim_m3_1_9/Cout 0.014
R31101 VSS.n10492 VSS.n10490 0.014
R31102 VSS.n6899 VSS.n6898 0.013
R31103 VSS.n17528 VSS.n17527 0.013
R31104 VSS.n17488 VSS.n17487 0.013
R31105 VSS.n13968 VSS.n13967 0.013
R31106 VSS.n10375 VSS.n10374 0.013
R31107 VSS.n6610 VSS.n6609 0.013
R31108 VSS.n3087 VSS.n3086 0.013
R31109 VSS.n3060 VSS.n3059 0.013
R31110 VSS.n17598 VSS.n17597 0.013
R31111 VSS.n17543 VSS.n17542 0.012
R31112 VSS.n17539 VSS.n17538 0.012
R31113 VSS.n17535 VSS.n17534 0.012
R31114 VSS.n17503 VSS.n17502 0.012
R31115 VSS.n17499 VSS.n17498 0.012
R31116 VSS.n17495 VSS.n17494 0.012
R31117 VSS.n13983 VSS.n13982 0.012
R31118 VSS.n13979 VSS.n13978 0.012
R31119 VSS.n13975 VSS.n13974 0.012
R31120 VSS.n10390 VSS.n10389 0.012
R31121 VSS.n10386 VSS.n10385 0.012
R31122 VSS.n10382 VSS.n10381 0.012
R31123 VSS.n6625 VSS.n6624 0.012
R31124 VSS.n6621 VSS.n6620 0.012
R31125 VSS.n6617 VSS.n6616 0.012
R31126 VSS.n3102 VSS.n3101 0.012
R31127 VSS.n3098 VSS.n3097 0.012
R31128 VSS.n3094 VSS.n3093 0.012
R31129 VSS.n3075 VSS.n3074 0.012
R31130 VSS.n3071 VSS.n3070 0.012
R31131 VSS.n3067 VSS.n3066 0.012
R31132 VSS.n17583 VSS.n17582 0.012
R31133 VSS.n17587 VSS.n17586 0.012
R31134 VSS.n17591 VSS.n17590 0.012
R31135 VSS.n17604 VSS.n17603 0.012
R31136 VSS.n17630 VSS.n17629 0.012
R31137 VSS.n14377 VSS.n14375 0.012
R31138 VSS.n14711 VSS.n14710 0.012
R31139 VSS.n14700 VSS.n14699 0.012
R31140 VSS.n14396 VSS.n14384 0.012
R31141 VSS.n14688 VSS.n14687 0.012
R31142 VSS.n14677 VSS.n14676 0.012
R31143 VSS.n14415 VSS.n14403 0.012
R31144 VSS.n14666 VSS.n14665 0.012
R31145 VSS.n14655 VSS.n14654 0.012
R31146 VSS.n14434 VSS.n14422 0.012
R31147 VSS.n14643 VSS.n14642 0.012
R31148 VSS.n14632 VSS.n14631 0.012
R31149 VSS.n14489 VSS.n14475 0.012
R31150 VSS.n14619 VSS.n14618 0.012
R31151 VSS.n14608 VSS.n14607 0.012
R31152 VSS.n14508 VSS.n14496 0.012
R31153 VSS.n14596 VSS.n14595 0.012
R31154 VSS.n14585 VSS.n14584 0.012
R31155 VSS.n14527 VSS.n14515 0.012
R31156 VSS.n14574 VSS.n14573 0.012
R31157 VSS.n14563 VSS.n14562 0.012
R31158 VSS.n14550 VSS.n14534 0.012
R31159 VSS.n14551 VSS.n14307 0.012
R31160 VSS.n14868 VSS.n14867 0.012
R31161 VSS.n14881 VSS.n14880 0.012
R31162 VSS.n14892 VSS.n14291 0.012
R31163 VSS.n14903 VSS.n14285 0.012
R31164 VSS.n14904 VSS.n14277 0.012
R31165 VSS.n14916 VSS.n14915 0.012
R31166 VSS.n14927 VSS.n14270 0.012
R31167 VSS.n14937 VSS.n14264 0.012
R31168 VSS.n14938 VSS.n14256 0.012
R31169 VSS.n14950 VSS.n14949 0.012
R31170 VSS.n14961 VSS.n14249 0.012
R31171 VSS.n14972 VSS.n14243 0.012
R31172 VSS.n15326 VSS.n15325 0.012
R31173 VSS.n14986 VSS.n14973 0.012
R31174 VSS.n15312 VSS.n15311 0.012
R31175 VSS.n15301 VSS.n15300 0.012
R31176 VSS.n15005 VSS.n14993 0.012
R31177 VSS.n15289 VSS.n15288 0.012
R31178 VSS.n15278 VSS.n15277 0.012
R31179 VSS.n15024 VSS.n15012 0.012
R31180 VSS.n15267 VSS.n15266 0.012
R31181 VSS.n15256 VSS.n15255 0.012
R31182 VSS.n15043 VSS.n15031 0.012
R31183 VSS.n15244 VSS.n15243 0.012
R31184 VSS.n15233 VSS.n15232 0.012
R31185 VSS.n15098 VSS.n15084 0.012
R31186 VSS.n15220 VSS.n15219 0.012
R31187 VSS.n15209 VSS.n15208 0.012
R31188 VSS.n15117 VSS.n15105 0.012
R31189 VSS.n15197 VSS.n15196 0.012
R31190 VSS.n15186 VSS.n15185 0.012
R31191 VSS.n15136 VSS.n15124 0.012
R31192 VSS.n15175 VSS.n15174 0.012
R31193 VSS.n15164 VSS.n15163 0.012
R31194 VSS.n15152 VSS.n15143 0.012
R31195 VSS.n15449 VSS.n14138 0.012
R31196 VSS.n15451 VSS.n14135 0.012
R31197 VSS.n15466 VSS.n14129 0.012
R31198 VSS.n15467 VSS.n14121 0.012
R31199 VSS.n15479 VSS.n15478 0.012
R31200 VSS.n15490 VSS.n14114 0.012
R31201 VSS.n15501 VSS.n14108 0.012
R31202 VSS.n15502 VSS.n14100 0.012
R31203 VSS.n15513 VSS.n15512 0.012
R31204 VSS.n15524 VSS.n14093 0.012
R31205 VSS.n15535 VSS.n14087 0.012
R31206 VSS.n15536 VSS.n14079 0.012
R31207 VSS.n15548 VSS.n15547 0.012
R31208 VSS.n15559 VSS.n15558 0.012
R31209 VSS.n15573 VSS.n15560 0.012
R31210 VSS.n15879 VSS.n15878 0.012
R31211 VSS.n15868 VSS.n15867 0.012
R31212 VSS.n15592 VSS.n15580 0.012
R31213 VSS.n15856 VSS.n15855 0.012
R31214 VSS.n15845 VSS.n15844 0.012
R31215 VSS.n15611 VSS.n15599 0.012
R31216 VSS.n15834 VSS.n15833 0.012
R31217 VSS.n15823 VSS.n15822 0.012
R31218 VSS.n15630 VSS.n15618 0.012
R31219 VSS.n15811 VSS.n15810 0.012
R31220 VSS.n15800 VSS.n15799 0.012
R31221 VSS.n15685 VSS.n15671 0.012
R31222 VSS.n15787 VSS.n15786 0.012
R31223 VSS.n15776 VSS.n15775 0.012
R31224 VSS.n15704 VSS.n15692 0.012
R31225 VSS.n15764 VSS.n15763 0.012
R31226 VSS.n15753 VSS.n15752 0.012
R31227 VSS.n15723 VSS.n15711 0.012
R31228 VSS.n15742 VSS.n15741 0.012
R31229 VSS.n15731 VSS.n13995 0.012
R31230 VSS.n14007 VSS.n13996 0.012
R31231 VSS.n16012 VSS.n16011 0.012
R31232 VSS.n16001 VSS.n16000 0.012
R31233 VSS.n16689 VSS.n16688 0.012
R31234 VSS.n16756 VSS.n16755 0.012
R31235 VSS.n16747 VSS.n16746 0.012
R31236 VSS.n16740 VSS.n16692 0.012
R31237 VSS.n16734 VSS.n16698 0.012
R31238 VSS.n16728 VSS.n16702 0.012
R31239 VSS.n16722 VSS.n16706 0.012
R31240 VSS.n16717 VSS.n16709 0.012
R31241 VSS.n16712 VSS.n16592 0.012
R31242 VSS.n16779 VSS.n16778 0.012
R31243 VSS.n16846 VSS.n16845 0.012
R31244 VSS.n16837 VSS.n16836 0.012
R31245 VSS.n16830 VSS.n16782 0.012
R31246 VSS.n16824 VSS.n16788 0.012
R31247 VSS.n16818 VSS.n16792 0.012
R31248 VSS.n16812 VSS.n16796 0.012
R31249 VSS.n16807 VSS.n16799 0.012
R31250 VSS.n16802 VSS.n16502 0.012
R31251 VSS.n16869 VSS.n16868 0.012
R31252 VSS.n16936 VSS.n16935 0.012
R31253 VSS.n16927 VSS.n16926 0.012
R31254 VSS.n16920 VSS.n16872 0.012
R31255 VSS.n16914 VSS.n16878 0.012
R31256 VSS.n16908 VSS.n16882 0.012
R31257 VSS.n16902 VSS.n16886 0.012
R31258 VSS.n16897 VSS.n16889 0.012
R31259 VSS.n16892 VSS.n16412 0.012
R31260 VSS.n16959 VSS.n16958 0.012
R31261 VSS.n17026 VSS.n17025 0.012
R31262 VSS.n17017 VSS.n17016 0.012
R31263 VSS.n17010 VSS.n16962 0.012
R31264 VSS.n17004 VSS.n16968 0.012
R31265 VSS.n16998 VSS.n16972 0.012
R31266 VSS.n16992 VSS.n16976 0.012
R31267 VSS.n16987 VSS.n16979 0.012
R31268 VSS.n16982 VSS.n16322 0.012
R31269 VSS.n17049 VSS.n17048 0.012
R31270 VSS.n17116 VSS.n17115 0.012
R31271 VSS.n17107 VSS.n17106 0.012
R31272 VSS.n17100 VSS.n17052 0.012
R31273 VSS.n17094 VSS.n17058 0.012
R31274 VSS.n17088 VSS.n17062 0.012
R31275 VSS.n17082 VSS.n17066 0.012
R31276 VSS.n17077 VSS.n17069 0.012
R31277 VSS.n17072 VSS.n16232 0.012
R31278 VSS.n17139 VSS.n17138 0.012
R31279 VSS.n17206 VSS.n17205 0.012
R31280 VSS.n17197 VSS.n17196 0.012
R31281 VSS.n17190 VSS.n17142 0.012
R31282 VSS.n17184 VSS.n17148 0.012
R31283 VSS.n17178 VSS.n17152 0.012
R31284 VSS.n17172 VSS.n17156 0.012
R31285 VSS.n17167 VSS.n17159 0.012
R31286 VSS.n17162 VSS.n16142 0.012
R31287 VSS.n17229 VSS.n17228 0.012
R31288 VSS.n17296 VSS.n17295 0.012
R31289 VSS.n17287 VSS.n17286 0.012
R31290 VSS.n17280 VSS.n17232 0.012
R31291 VSS.n17274 VSS.n17238 0.012
R31292 VSS.n17268 VSS.n17242 0.012
R31293 VSS.n17262 VSS.n17246 0.012
R31294 VSS.n17257 VSS.n17249 0.012
R31295 VSS.n17252 VSS.n16052 0.012
R31296 VSS.n17390 VSS.n17389 0.012
R31297 VSS.n17398 VSS.n17397 0.012
R31298 VSS.n17452 VSS.n17451 0.012
R31299 VSS.n17443 VSS.n17442 0.012
R31300 VSS.n17436 VSS.n17401 0.012
R31301 VSS.n17430 VSS.n17407 0.012
R31302 VSS.n17424 VSS.n17411 0.012
R31303 VSS.n17418 VSS.n16025 0.012
R31304 VSS.n17332 VSS.n16026 0.012
R31305 VSS.n12802 VSS.n12718 0.012
R31306 VSS.n12813 VSS.n12712 0.012
R31307 VSS.n12814 VSS.n12704 0.012
R31308 VSS.n12826 VSS.n12825 0.012
R31309 VSS.n12837 VSS.n12697 0.012
R31310 VSS.n12848 VSS.n12691 0.012
R31311 VSS.n12849 VSS.n12683 0.012
R31312 VSS.n12860 VSS.n12859 0.012
R31313 VSS.n12871 VSS.n12676 0.012
R31314 VSS.n12883 VSS.n12668 0.012
R31315 VSS.n12885 VSS.n12661 0.012
R31316 VSS.n13063 VSS.n13062 0.012
R31317 VSS.n13050 VSS.n13049 0.012
R31318 VSS.n13039 VSS.n13038 0.012
R31319 VSS.n12914 VSS.n12902 0.012
R31320 VSS.n13027 VSS.n13026 0.012
R31321 VSS.n13016 VSS.n13015 0.012
R31322 VSS.n12933 VSS.n12921 0.012
R31323 VSS.n13005 VSS.n13004 0.012
R31324 VSS.n12994 VSS.n12993 0.012
R31325 VSS.n12952 VSS.n12940 0.012
R31326 VSS.n12982 VSS.n12981 0.012
R31327 VSS.n12971 VSS.n12970 0.012
R31328 VSS.n12960 VSS.n12959 0.012
R31329 VSS.n13159 VSS.n12577 0.012
R31330 VSS.n13170 VSS.n12571 0.012
R31331 VSS.n13171 VSS.n12563 0.012
R31332 VSS.n13183 VSS.n13182 0.012
R31333 VSS.n13194 VSS.n12556 0.012
R31334 VSS.n13205 VSS.n12550 0.012
R31335 VSS.n13206 VSS.n12542 0.012
R31336 VSS.n13217 VSS.n13216 0.012
R31337 VSS.n13228 VSS.n12535 0.012
R31338 VSS.n13240 VSS.n12527 0.012
R31339 VSS.n13242 VSS.n12520 0.012
R31340 VSS.n13312 VSS.n13311 0.012
R31341 VSS.n13299 VSS.n13298 0.012
R31342 VSS.n13288 VSS.n13287 0.012
R31343 VSS.n13275 VSS.n13259 0.012
R31344 VSS.n13276 VSS.n11429 0.012
R31345 VSS.n11441 VSS.n11430 0.012
R31346 VSS.n13446 VSS.n13445 0.012
R31347 VSS.n13436 VSS.n13435 0.012
R31348 VSS.n11460 VSS.n11448 0.012
R31349 VSS.n13424 VSS.n13423 0.012
R31350 VSS.n13413 VSS.n13412 0.012
R31351 VSS.n11479 VSS.n11467 0.012
R31352 VSS.n13401 VSS.n13400 0.012
R31353 VSS.n11680 VSS.n11668 0.012
R31354 VSS.n11691 VSS.n11662 0.012
R31355 VSS.n11692 VSS.n11654 0.012
R31356 VSS.n11704 VSS.n11703 0.012
R31357 VSS.n11715 VSS.n11647 0.012
R31358 VSS.n11726 VSS.n11641 0.012
R31359 VSS.n11727 VSS.n11633 0.012
R31360 VSS.n11738 VSS.n11737 0.012
R31361 VSS.n11749 VSS.n11626 0.012
R31362 VSS.n11760 VSS.n11620 0.012
R31363 VSS.n11761 VSS.n11611 0.012
R31364 VSS.n11773 VSS.n11772 0.012
R31365 VSS.n11815 VSS.n11814 0.012
R31366 VSS.n11826 VSS.n11596 0.012
R31367 VSS.n11837 VSS.n11590 0.012
R31368 VSS.n11838 VSS.n11582 0.012
R31369 VSS.n11850 VSS.n11849 0.012
R31370 VSS.n11861 VSS.n11575 0.012
R31371 VSS.n11871 VSS.n11569 0.012
R31372 VSS.n11872 VSS.n11561 0.012
R31373 VSS.n11884 VSS.n11883 0.012
R31374 VSS.n11895 VSS.n11554 0.012
R31375 VSS.n11906 VSS.n11548 0.012
R31376 VSS.n12401 VSS.n12400 0.012
R31377 VSS.n11920 VSS.n11907 0.012
R31378 VSS.n12387 VSS.n12386 0.012
R31379 VSS.n12376 VSS.n12375 0.012
R31380 VSS.n11939 VSS.n11927 0.012
R31381 VSS.n12364 VSS.n12363 0.012
R31382 VSS.n12353 VSS.n12352 0.012
R31383 VSS.n11958 VSS.n11946 0.012
R31384 VSS.n12342 VSS.n12341 0.012
R31385 VSS.n12331 VSS.n12330 0.012
R31386 VSS.n11977 VSS.n11965 0.012
R31387 VSS.n12319 VSS.n12318 0.012
R31388 VSS.n12308 VSS.n12307 0.012
R31389 VSS.n11999 VSS.n11985 0.012
R31390 VSS.n12295 VSS.n12294 0.012
R31391 VSS.n12284 VSS.n12283 0.012
R31392 VSS.n12018 VSS.n12006 0.012
R31393 VSS.n12272 VSS.n12271 0.012
R31394 VSS.n12261 VSS.n12260 0.012
R31395 VSS.n12037 VSS.n12025 0.012
R31396 VSS.n12250 VSS.n12249 0.012
R31397 VSS.n12239 VSS.n12238 0.012
R31398 VSS.n12056 VSS.n12044 0.012
R31399 VSS.n12227 VSS.n12226 0.012
R31400 VSS.n12216 VSS.n12215 0.012
R31401 VSS.n11156 VSS.n11155 0.012
R31402 VSS.n11224 VSS.n11223 0.012
R31403 VSS.n11215 VSS.n11214 0.012
R31404 VSS.n11208 VSS.n11159 0.012
R31405 VSS.n11202 VSS.n11165 0.012
R31406 VSS.n11196 VSS.n11169 0.012
R31407 VSS.n11191 VSS.n11172 0.012
R31408 VSS.n11185 VSS.n11175 0.012
R31409 VSS.n11178 VSS.n11059 0.012
R31410 VSS.n11246 VSS.n11245 0.012
R31411 VSS.n11314 VSS.n11313 0.012
R31412 VSS.n11305 VSS.n11304 0.012
R31413 VSS.n11298 VSS.n11249 0.012
R31414 VSS.n11292 VSS.n11255 0.012
R31415 VSS.n11286 VSS.n11259 0.012
R31416 VSS.n11281 VSS.n11262 0.012
R31417 VSS.n11275 VSS.n11265 0.012
R31418 VSS.n11268 VSS.n10969 0.012
R31419 VSS.n11336 VSS.n11335 0.012
R31420 VSS.n11404 VSS.n11403 0.012
R31421 VSS.n11395 VSS.n11394 0.012
R31422 VSS.n11388 VSS.n11339 0.012
R31423 VSS.n11382 VSS.n11345 0.012
R31424 VSS.n11376 VSS.n11349 0.012
R31425 VSS.n11371 VSS.n11352 0.012
R31426 VSS.n11365 VSS.n11355 0.012
R31427 VSS.n11358 VSS.n10879 0.012
R31428 VSS.n11426 VSS.n11425 0.012
R31429 VSS.n13524 VSS.n13523 0.012
R31430 VSS.n13515 VSS.n13514 0.012
R31431 VSS.n13507 VSS.n13458 0.012
R31432 VSS.n13501 VSS.n13464 0.012
R31433 VSS.n13495 VSS.n13468 0.012
R31434 VSS.n13490 VSS.n13471 0.012
R31435 VSS.n13484 VSS.n13474 0.012
R31436 VSS.n13477 VSS.n10789 0.012
R31437 VSS.n13546 VSS.n13545 0.012
R31438 VSS.n13614 VSS.n13613 0.012
R31439 VSS.n13605 VSS.n13604 0.012
R31440 VSS.n13598 VSS.n13549 0.012
R31441 VSS.n13592 VSS.n13555 0.012
R31442 VSS.n13586 VSS.n13559 0.012
R31443 VSS.n13581 VSS.n13562 0.012
R31444 VSS.n13575 VSS.n13565 0.012
R31445 VSS.n13568 VSS.n10699 0.012
R31446 VSS.n13636 VSS.n13635 0.012
R31447 VSS.n13704 VSS.n13703 0.012
R31448 VSS.n13695 VSS.n13694 0.012
R31449 VSS.n13688 VSS.n13639 0.012
R31450 VSS.n13682 VSS.n13645 0.012
R31451 VSS.n13676 VSS.n13649 0.012
R31452 VSS.n13671 VSS.n13652 0.012
R31453 VSS.n13665 VSS.n13655 0.012
R31454 VSS.n13658 VSS.n10609 0.012
R31455 VSS.n13726 VSS.n13725 0.012
R31456 VSS.n13794 VSS.n13793 0.012
R31457 VSS.n13785 VSS.n13784 0.012
R31458 VSS.n13778 VSS.n13729 0.012
R31459 VSS.n13772 VSS.n13735 0.012
R31460 VSS.n13766 VSS.n13739 0.012
R31461 VSS.n13761 VSS.n13742 0.012
R31462 VSS.n13755 VSS.n13745 0.012
R31463 VSS.n13748 VSS.n10519 0.012
R31464 VSS.n13890 VSS.n13889 0.012
R31465 VSS.n13898 VSS.n13897 0.012
R31466 VSS.n13944 VSS.n13943 0.012
R31467 VSS.n13935 VSS.n13934 0.012
R31468 VSS.n13928 VSS.n13901 0.012
R31469 VSS.n13922 VSS.n13907 0.012
R31470 VSS.n13916 VSS.n13911 0.012
R31471 VSS.n13959 VSS.n10492 0.012
R31472 VSS.n13832 VSS.n13831 0.012
R31473 VSS.n7684 VSS.n7682 0.012
R31474 VSS.n7825 VSS.n7824 0.012
R31475 VSS.n7814 VSS.n7813 0.012
R31476 VSS.n7703 VSS.n7691 0.012
R31477 VSS.n7802 VSS.n7801 0.012
R31478 VSS.n7791 VSS.n7790 0.012
R31479 VSS.n7722 VSS.n7710 0.012
R31480 VSS.n7780 VSS.n7779 0.012
R31481 VSS.n7769 VSS.n7768 0.012
R31482 VSS.n7741 VSS.n7729 0.012
R31483 VSS.n7757 VSS.n7756 0.012
R31484 VSS.n7746 VSS.n7745 0.012
R31485 VSS.n7926 VSS.n7925 0.012
R31486 VSS.n7937 VSS.n7590 0.012
R31487 VSS.n7948 VSS.n7584 0.012
R31488 VSS.n7949 VSS.n7576 0.012
R31489 VSS.n7961 VSS.n7960 0.012
R31490 VSS.n7972 VSS.n7569 0.012
R31491 VSS.n7982 VSS.n7563 0.012
R31492 VSS.n7983 VSS.n7555 0.012
R31493 VSS.n7995 VSS.n7994 0.012
R31494 VSS.n8006 VSS.n7548 0.012
R31495 VSS.n8017 VSS.n7542 0.012
R31496 VSS.n8187 VSS.n8186 0.012
R31497 VSS.n8029 VSS.n8028 0.012
R31498 VSS.n8038 VSS.n8036 0.012
R31499 VSS.n8165 VSS.n8164 0.012
R31500 VSS.n8154 VSS.n8153 0.012
R31501 VSS.n8057 VSS.n8045 0.012
R31502 VSS.n8142 VSS.n8141 0.012
R31503 VSS.n8132 VSS.n8131 0.012
R31504 VSS.n8076 VSS.n8064 0.012
R31505 VSS.n8120 VSS.n8119 0.012
R31506 VSS.n8109 VSS.n8108 0.012
R31507 VSS.n8094 VSS.n8083 0.012
R31508 VSS.n8097 VSS.n8096 0.012
R31509 VSS.n8284 VSS.n8283 0.012
R31510 VSS.n8295 VSS.n7450 0.012
R31511 VSS.n8306 VSS.n7444 0.012
R31512 VSS.n8307 VSS.n7436 0.012
R31513 VSS.n8319 VSS.n8318 0.012
R31514 VSS.n8330 VSS.n7429 0.012
R31515 VSS.n8340 VSS.n7423 0.012
R31516 VSS.n8341 VSS.n7415 0.012
R31517 VSS.n8353 VSS.n8352 0.012
R31518 VSS.n8364 VSS.n7408 0.012
R31519 VSS.n8375 VSS.n7402 0.012
R31520 VSS.n8545 VSS.n8544 0.012
R31521 VSS.n8387 VSS.n8386 0.012
R31522 VSS.n8396 VSS.n8394 0.012
R31523 VSS.n8523 VSS.n8522 0.012
R31524 VSS.n8512 VSS.n8511 0.012
R31525 VSS.n8415 VSS.n8403 0.012
R31526 VSS.n8500 VSS.n8499 0.012
R31527 VSS.n8490 VSS.n8489 0.012
R31528 VSS.n8434 VSS.n8422 0.012
R31529 VSS.n8478 VSS.n8477 0.012
R31530 VSS.n8467 VSS.n8466 0.012
R31531 VSS.n8452 VSS.n8441 0.012
R31532 VSS.n8455 VSS.n8454 0.012
R31533 VSS.n8642 VSS.n8641 0.012
R31534 VSS.n8653 VSS.n7310 0.012
R31535 VSS.n8664 VSS.n7304 0.012
R31536 VSS.n8665 VSS.n7296 0.012
R31537 VSS.n8677 VSS.n8676 0.012
R31538 VSS.n8688 VSS.n7289 0.012
R31539 VSS.n8698 VSS.n7283 0.012
R31540 VSS.n8699 VSS.n7275 0.012
R31541 VSS.n8711 VSS.n8710 0.012
R31542 VSS.n8722 VSS.n7268 0.012
R31543 VSS.n8733 VSS.n7262 0.012
R31544 VSS.n8767 VSS.n8766 0.012
R31545 VSS.n8745 VSS.n8744 0.012
R31546 VSS.n8746 VSS.n6901 0.012
R31547 VSS.n6913 VSS.n6902 0.012
R31548 VSS.n8918 VSS.n8917 0.012
R31549 VSS.n8907 VSS.n8906 0.012
R31550 VSS.n6932 VSS.n6920 0.012
R31551 VSS.n8896 VSS.n8895 0.012
R31552 VSS.n8885 VSS.n8884 0.012
R31553 VSS.n6951 VSS.n6939 0.012
R31554 VSS.n8873 VSS.n8872 0.012
R31555 VSS.n8862 VSS.n8861 0.012
R31556 VSS.n7070 VSS.n6958 0.012
R31557 VSS.n7082 VSS.n7064 0.012
R31558 VSS.n7083 VSS.n7056 0.012
R31559 VSS.n7095 VSS.n7094 0.012
R31560 VSS.n7106 VSS.n7049 0.012
R31561 VSS.n7117 VSS.n7043 0.012
R31562 VSS.n7118 VSS.n7035 0.012
R31563 VSS.n7129 VSS.n7128 0.012
R31564 VSS.n7140 VSS.n7028 0.012
R31565 VSS.n7151 VSS.n7022 0.012
R31566 VSS.n7152 VSS.n7014 0.012
R31567 VSS.n7164 VSS.n7163 0.012
R31568 VSS.n7176 VSS.n7006 0.012
R31569 VSS.n9734 VSS.n9733 0.012
R31570 VSS.n9801 VSS.n9800 0.012
R31571 VSS.n9792 VSS.n9791 0.012
R31572 VSS.n9785 VSS.n9737 0.012
R31573 VSS.n9779 VSS.n9743 0.012
R31574 VSS.n9773 VSS.n9747 0.012
R31575 VSS.n9767 VSS.n9751 0.012
R31576 VSS.n9762 VSS.n9754 0.012
R31577 VSS.n9757 VSS.n9637 0.012
R31578 VSS.n9824 VSS.n9823 0.012
R31579 VSS.n9891 VSS.n9890 0.012
R31580 VSS.n9882 VSS.n9881 0.012
R31581 VSS.n9875 VSS.n9827 0.012
R31582 VSS.n9869 VSS.n9833 0.012
R31583 VSS.n9863 VSS.n9837 0.012
R31584 VSS.n9857 VSS.n9841 0.012
R31585 VSS.n9852 VSS.n9844 0.012
R31586 VSS.n9847 VSS.n9547 0.012
R31587 VSS.n9914 VSS.n9913 0.012
R31588 VSS.n9981 VSS.n9980 0.012
R31589 VSS.n9972 VSS.n9971 0.012
R31590 VSS.n9965 VSS.n9917 0.012
R31591 VSS.n9959 VSS.n9923 0.012
R31592 VSS.n9953 VSS.n9927 0.012
R31593 VSS.n9947 VSS.n9931 0.012
R31594 VSS.n9942 VSS.n9934 0.012
R31595 VSS.n9937 VSS.n9457 0.012
R31596 VSS.n10004 VSS.n10003 0.012
R31597 VSS.n10071 VSS.n10070 0.012
R31598 VSS.n10062 VSS.n10061 0.012
R31599 VSS.n10055 VSS.n10007 0.012
R31600 VSS.n10049 VSS.n10013 0.012
R31601 VSS.n10043 VSS.n10017 0.012
R31602 VSS.n10037 VSS.n10021 0.012
R31603 VSS.n10032 VSS.n10024 0.012
R31604 VSS.n10027 VSS.n9367 0.012
R31605 VSS.n10094 VSS.n10093 0.012
R31606 VSS.n10161 VSS.n10160 0.012
R31607 VSS.n10152 VSS.n10151 0.012
R31608 VSS.n10145 VSS.n10097 0.012
R31609 VSS.n10139 VSS.n10103 0.012
R31610 VSS.n10133 VSS.n10107 0.012
R31611 VSS.n10127 VSS.n10111 0.012
R31612 VSS.n10122 VSS.n10114 0.012
R31613 VSS.n10117 VSS.n9277 0.012
R31614 VSS.n10184 VSS.n10183 0.012
R31615 VSS.n10251 VSS.n10250 0.012
R31616 VSS.n10242 VSS.n10241 0.012
R31617 VSS.n10235 VSS.n10187 0.012
R31618 VSS.n10229 VSS.n10193 0.012
R31619 VSS.n10223 VSS.n10197 0.012
R31620 VSS.n10217 VSS.n10201 0.012
R31621 VSS.n10212 VSS.n10204 0.012
R31622 VSS.n10207 VSS.n9187 0.012
R31623 VSS.n10319 VSS.n8930 0.012
R31624 VSS.n8939 VSS.n8931 0.012
R31625 VSS.n8945 VSS.n8944 0.012
R31626 VSS.n8951 VSS.n8950 0.012
R31627 VSS.n8956 VSS.n8955 0.012
R31628 VSS.n8963 VSS.n8962 0.012
R31629 VSS.n8969 VSS.n8968 0.012
R31630 VSS.n8975 VSS.n8974 0.012
R31631 VSS.n8980 VSS.n8979 0.012
R31632 VSS.n9040 VSS.n9033 0.012
R31633 VSS.n9048 VSS.n9031 0.012
R31634 VSS.n9056 VSS.n9029 0.012
R31635 VSS.n9064 VSS.n9027 0.012
R31636 VSS.n9072 VSS.n9025 0.012
R31637 VSS.n9080 VSS.n9023 0.012
R31638 VSS.n9088 VSS.n9021 0.012
R31639 VSS.n9096 VSS.n9019 0.012
R31640 VSS.n9151 VSS.n9150 0.012
R31641 VSS.n4255 VSS.n4171 0.012
R31642 VSS.n4266 VSS.n4165 0.012
R31643 VSS.n4267 VSS.n4157 0.012
R31644 VSS.n4279 VSS.n4278 0.012
R31645 VSS.n4290 VSS.n4150 0.012
R31646 VSS.n4301 VSS.n4144 0.012
R31647 VSS.n4302 VSS.n4136 0.012
R31648 VSS.n4313 VSS.n4312 0.012
R31649 VSS.n4324 VSS.n4129 0.012
R31650 VSS.n4336 VSS.n4121 0.012
R31651 VSS.n4338 VSS.n4114 0.012
R31652 VSS.n4516 VSS.n4515 0.012
R31653 VSS.n4503 VSS.n4502 0.012
R31654 VSS.n4492 VSS.n4491 0.012
R31655 VSS.n4367 VSS.n4355 0.012
R31656 VSS.n4480 VSS.n4479 0.012
R31657 VSS.n4469 VSS.n4468 0.012
R31658 VSS.n4386 VSS.n4374 0.012
R31659 VSS.n4458 VSS.n4457 0.012
R31660 VSS.n4447 VSS.n4446 0.012
R31661 VSS.n4405 VSS.n4393 0.012
R31662 VSS.n4435 VSS.n4434 0.012
R31663 VSS.n4424 VSS.n4423 0.012
R31664 VSS.n4413 VSS.n4412 0.012
R31665 VSS.n4612 VSS.n4030 0.012
R31666 VSS.n4623 VSS.n4024 0.012
R31667 VSS.n4624 VSS.n4016 0.012
R31668 VSS.n4636 VSS.n4635 0.012
R31669 VSS.n4647 VSS.n4009 0.012
R31670 VSS.n4658 VSS.n4003 0.012
R31671 VSS.n4659 VSS.n3995 0.012
R31672 VSS.n4670 VSS.n4669 0.012
R31673 VSS.n4681 VSS.n3988 0.012
R31674 VSS.n4693 VSS.n3980 0.012
R31675 VSS.n4695 VSS.n3973 0.012
R31676 VSS.n4873 VSS.n4872 0.012
R31677 VSS.n4860 VSS.n4859 0.012
R31678 VSS.n4849 VSS.n4848 0.012
R31679 VSS.n4724 VSS.n4712 0.012
R31680 VSS.n4837 VSS.n4836 0.012
R31681 VSS.n4826 VSS.n4825 0.012
R31682 VSS.n4743 VSS.n4731 0.012
R31683 VSS.n4815 VSS.n4814 0.012
R31684 VSS.n4804 VSS.n4803 0.012
R31685 VSS.n4762 VSS.n4750 0.012
R31686 VSS.n4792 VSS.n4791 0.012
R31687 VSS.n4781 VSS.n4780 0.012
R31688 VSS.n4770 VSS.n4769 0.012
R31689 VSS.n4969 VSS.n3889 0.012
R31690 VSS.n4980 VSS.n3883 0.012
R31691 VSS.n4981 VSS.n3875 0.012
R31692 VSS.n4993 VSS.n4992 0.012
R31693 VSS.n5004 VSS.n3868 0.012
R31694 VSS.n5015 VSS.n3862 0.012
R31695 VSS.n5016 VSS.n3854 0.012
R31696 VSS.n5027 VSS.n5026 0.012
R31697 VSS.n5038 VSS.n3847 0.012
R31698 VSS.n5050 VSS.n3839 0.012
R31699 VSS.n5052 VSS.n3832 0.012
R31700 VSS.n5230 VSS.n5229 0.012
R31701 VSS.n5217 VSS.n5216 0.012
R31702 VSS.n5206 VSS.n5205 0.012
R31703 VSS.n5081 VSS.n5069 0.012
R31704 VSS.n5194 VSS.n5193 0.012
R31705 VSS.n5183 VSS.n5182 0.012
R31706 VSS.n5100 VSS.n5088 0.012
R31707 VSS.n5172 VSS.n5171 0.012
R31708 VSS.n5161 VSS.n5160 0.012
R31709 VSS.n5119 VSS.n5107 0.012
R31710 VSS.n5149 VSS.n5148 0.012
R31711 VSS.n5138 VSS.n5137 0.012
R31712 VSS.n5127 VSS.n5126 0.012
R31713 VSS.n5326 VSS.n3748 0.012
R31714 VSS.n5337 VSS.n3742 0.012
R31715 VSS.n5338 VSS.n3734 0.012
R31716 VSS.n5350 VSS.n5349 0.012
R31717 VSS.n5361 VSS.n3727 0.012
R31718 VSS.n5372 VSS.n3721 0.012
R31719 VSS.n5373 VSS.n3713 0.012
R31720 VSS.n5384 VSS.n5383 0.012
R31721 VSS.n5395 VSS.n3706 0.012
R31722 VSS.n5407 VSS.n3698 0.012
R31723 VSS.n5409 VSS.n3691 0.012
R31724 VSS.n5576 VSS.n5575 0.012
R31725 VSS.n5563 VSS.n5562 0.012
R31726 VSS.n5552 VSS.n5551 0.012
R31727 VSS.n5438 VSS.n5426 0.012
R31728 VSS.n5540 VSS.n5539 0.012
R31729 VSS.n5529 VSS.n5528 0.012
R31730 VSS.n5457 VSS.n5445 0.012
R31731 VSS.n5518 VSS.n5517 0.012
R31732 VSS.n5507 VSS.n5506 0.012
R31733 VSS.n5476 VSS.n5464 0.012
R31734 VSS.n5495 VSS.n5494 0.012
R31735 VSS.n5484 VSS.n3635 0.012
R31736 VSS.n3646 VSS.n3636 0.012
R31737 VSS.n6604 VSS.n3137 0.012
R31738 VSS.n3180 VSS.n3173 0.012
R31739 VSS.n3188 VSS.n3171 0.012
R31740 VSS.n3196 VSS.n3169 0.012
R31741 VSS.n3204 VSS.n3167 0.012
R31742 VSS.n3212 VSS.n3165 0.012
R31743 VSS.n3220 VSS.n3163 0.012
R31744 VSS.n3228 VSS.n3161 0.012
R31745 VSS.n6593 VSS.n6592 0.012
R31746 VSS.n3238 VSS.n3230 0.012
R31747 VSS.n3244 VSS.n3243 0.012
R31748 VSS.n3250 VSS.n3249 0.012
R31749 VSS.n3256 VSS.n3255 0.012
R31750 VSS.n3261 VSS.n3260 0.012
R31751 VSS.n3268 VSS.n3267 0.012
R31752 VSS.n3274 VSS.n3273 0.012
R31753 VSS.n3280 VSS.n3279 0.012
R31754 VSS.n3286 VSS.n3285 0.012
R31755 VSS.n3296 VSS.n3288 0.012
R31756 VSS.n3302 VSS.n3301 0.012
R31757 VSS.n3308 VSS.n3307 0.012
R31758 VSS.n3314 VSS.n3313 0.012
R31759 VSS.n3319 VSS.n3318 0.012
R31760 VSS.n3326 VSS.n3325 0.012
R31761 VSS.n3332 VSS.n3331 0.012
R31762 VSS.n3338 VSS.n3337 0.012
R31763 VSS.n3344 VSS.n3343 0.012
R31764 VSS.n3354 VSS.n3346 0.012
R31765 VSS.n3360 VSS.n3359 0.012
R31766 VSS.n3366 VSS.n3365 0.012
R31767 VSS.n3372 VSS.n3371 0.012
R31768 VSS.n3377 VSS.n3376 0.012
R31769 VSS.n3384 VSS.n3383 0.012
R31770 VSS.n3390 VSS.n3389 0.012
R31771 VSS.n3396 VSS.n3395 0.012
R31772 VSS.n3402 VSS.n3401 0.012
R31773 VSS.n3412 VSS.n3404 0.012
R31774 VSS.n3418 VSS.n3417 0.012
R31775 VSS.n3424 VSS.n3423 0.012
R31776 VSS.n3430 VSS.n3429 0.012
R31777 VSS.n3435 VSS.n3434 0.012
R31778 VSS.n3442 VSS.n3441 0.012
R31779 VSS.n3448 VSS.n3447 0.012
R31780 VSS.n3454 VSS.n3453 0.012
R31781 VSS.n3460 VSS.n3459 0.012
R31782 VSS.n3470 VSS.n3462 0.012
R31783 VSS.n3476 VSS.n3475 0.012
R31784 VSS.n3482 VSS.n3481 0.012
R31785 VSS.n3488 VSS.n3487 0.012
R31786 VSS.n3493 VSS.n3492 0.012
R31787 VSS.n3500 VSS.n3499 0.012
R31788 VSS.n3506 VSS.n3505 0.012
R31789 VSS.n3512 VSS.n3511 0.012
R31790 VSS.n3518 VSS.n3517 0.012
R31791 VSS.n3528 VSS.n3520 0.012
R31792 VSS.n3534 VSS.n3533 0.012
R31793 VSS.n3540 VSS.n3539 0.012
R31794 VSS.n3546 VSS.n3545 0.012
R31795 VSS.n3551 VSS.n3550 0.012
R31796 VSS.n3558 VSS.n3557 0.012
R31797 VSS.n3564 VSS.n3563 0.012
R31798 VSS.n3570 VSS.n3569 0.012
R31799 VSS.n3576 VSS.n3575 0.012
R31800 VSS.n3586 VSS.n3578 0.012
R31801 VSS.n3592 VSS.n3591 0.012
R31802 VSS.n3598 VSS.n3597 0.012
R31803 VSS.n3604 VSS.n3603 0.012
R31804 VSS.n3609 VSS.n3608 0.012
R31805 VSS.n3616 VSS.n3615 0.012
R31806 VSS.n3622 VSS.n3621 0.012
R31807 VSS.n3628 VSS.n3627 0.012
R31808 VSS.n3634 VSS.n3633 0.012
R31809 VSS.n1618 VSS.n1616 0.012
R31810 VSS.n1952 VSS.n1951 0.012
R31811 VSS.n1941 VSS.n1940 0.012
R31812 VSS.n1637 VSS.n1625 0.012
R31813 VSS.n1929 VSS.n1928 0.012
R31814 VSS.n1918 VSS.n1917 0.012
R31815 VSS.n1656 VSS.n1644 0.012
R31816 VSS.n1907 VSS.n1906 0.012
R31817 VSS.n1896 VSS.n1895 0.012
R31818 VSS.n1675 VSS.n1663 0.012
R31819 VSS.n1884 VSS.n1883 0.012
R31820 VSS.n1873 VSS.n1872 0.012
R31821 VSS.n1730 VSS.n1716 0.012
R31822 VSS.n1860 VSS.n1859 0.012
R31823 VSS.n1849 VSS.n1848 0.012
R31824 VSS.n1749 VSS.n1737 0.012
R31825 VSS.n1837 VSS.n1836 0.012
R31826 VSS.n1826 VSS.n1825 0.012
R31827 VSS.n1768 VSS.n1756 0.012
R31828 VSS.n1815 VSS.n1814 0.012
R31829 VSS.n1804 VSS.n1803 0.012
R31830 VSS.n1791 VSS.n1775 0.012
R31831 VSS.n1792 VSS.n1548 0.012
R31832 VSS.n2109 VSS.n2108 0.012
R31833 VSS.n2122 VSS.n2121 0.012
R31834 VSS.n2133 VSS.n1532 0.012
R31835 VSS.n2144 VSS.n1526 0.012
R31836 VSS.n2145 VSS.n1518 0.012
R31837 VSS.n2157 VSS.n2156 0.012
R31838 VSS.n2168 VSS.n1511 0.012
R31839 VSS.n2178 VSS.n1505 0.012
R31840 VSS.n2179 VSS.n1497 0.012
R31841 VSS.n2191 VSS.n2190 0.012
R31842 VSS.n2202 VSS.n1490 0.012
R31843 VSS.n2213 VSS.n1484 0.012
R31844 VSS.n2567 VSS.n2566 0.012
R31845 VSS.n2227 VSS.n2214 0.012
R31846 VSS.n2553 VSS.n2552 0.012
R31847 VSS.n2542 VSS.n2541 0.012
R31848 VSS.n2246 VSS.n2234 0.012
R31849 VSS.n2530 VSS.n2529 0.012
R31850 VSS.n2519 VSS.n2518 0.012
R31851 VSS.n2265 VSS.n2253 0.012
R31852 VSS.n2508 VSS.n2507 0.012
R31853 VSS.n2497 VSS.n2496 0.012
R31854 VSS.n2284 VSS.n2272 0.012
R31855 VSS.n2485 VSS.n2484 0.012
R31856 VSS.n2474 VSS.n2473 0.012
R31857 VSS.n2339 VSS.n2325 0.012
R31858 VSS.n2461 VSS.n2460 0.012
R31859 VSS.n2450 VSS.n2449 0.012
R31860 VSS.n2358 VSS.n2346 0.012
R31861 VSS.n2438 VSS.n2437 0.012
R31862 VSS.n2427 VSS.n2426 0.012
R31863 VSS.n2377 VSS.n2365 0.012
R31864 VSS.n2416 VSS.n2415 0.012
R31865 VSS.n2405 VSS.n2404 0.012
R31866 VSS.n2393 VSS.n2384 0.012
R31867 VSS.n2690 VSS.n1379 0.012
R31868 VSS.n2692 VSS.n1376 0.012
R31869 VSS.n2707 VSS.n1370 0.012
R31870 VSS.n2708 VSS.n1362 0.012
R31871 VSS.n2720 VSS.n2719 0.012
R31872 VSS.n2731 VSS.n1355 0.012
R31873 VSS.n2742 VSS.n1349 0.012
R31874 VSS.n2743 VSS.n1341 0.012
R31875 VSS.n2754 VSS.n2753 0.012
R31876 VSS.n2765 VSS.n1334 0.012
R31877 VSS.n2776 VSS.n1328 0.012
R31878 VSS.n2777 VSS.n1320 0.012
R31879 VSS.n2789 VSS.n2788 0.012
R31880 VSS.n2800 VSS.n2799 0.012
R31881 VSS.n2814 VSS.n2801 0.012
R31882 VSS.n2953 VSS.n2952 0.012
R31883 VSS.n2942 VSS.n2941 0.012
R31884 VSS.n2833 VSS.n2821 0.012
R31885 VSS.n2930 VSS.n2929 0.012
R31886 VSS.n2919 VSS.n2918 0.012
R31887 VSS.n2852 VSS.n2840 0.012
R31888 VSS.n2908 VSS.n2907 0.012
R31889 VSS.n2897 VSS.n2896 0.012
R31890 VSS.n2871 VSS.n2859 0.012
R31891 VSS.n2885 VSS.n2884 0.012
R31892 VSS.n2874 VSS.n2873 0.012
R31893 VSS.n642 VSS.n641 0.012
R31894 VSS.n709 VSS.n708 0.012
R31895 VSS.n700 VSS.n699 0.012
R31896 VSS.n693 VSS.n645 0.012
R31897 VSS.n687 VSS.n651 0.012
R31898 VSS.n681 VSS.n655 0.012
R31899 VSS.n675 VSS.n659 0.012
R31900 VSS.n670 VSS.n662 0.012
R31901 VSS.n665 VSS.n545 0.012
R31902 VSS.n732 VSS.n731 0.012
R31903 VSS.n799 VSS.n798 0.012
R31904 VSS.n790 VSS.n789 0.012
R31905 VSS.n783 VSS.n735 0.012
R31906 VSS.n777 VSS.n741 0.012
R31907 VSS.n771 VSS.n745 0.012
R31908 VSS.n765 VSS.n749 0.012
R31909 VSS.n760 VSS.n752 0.012
R31910 VSS.n755 VSS.n455 0.012
R31911 VSS.n822 VSS.n821 0.012
R31912 VSS.n889 VSS.n888 0.012
R31913 VSS.n880 VSS.n879 0.012
R31914 VSS.n873 VSS.n825 0.012
R31915 VSS.n867 VSS.n831 0.012
R31916 VSS.n861 VSS.n835 0.012
R31917 VSS.n855 VSS.n839 0.012
R31918 VSS.n850 VSS.n842 0.012
R31919 VSS.n845 VSS.n365 0.012
R31920 VSS.n912 VSS.n911 0.012
R31921 VSS.n979 VSS.n978 0.012
R31922 VSS.n970 VSS.n969 0.012
R31923 VSS.n963 VSS.n915 0.012
R31924 VSS.n957 VSS.n921 0.012
R31925 VSS.n951 VSS.n925 0.012
R31926 VSS.n945 VSS.n929 0.012
R31927 VSS.n940 VSS.n932 0.012
R31928 VSS.n935 VSS.n275 0.012
R31929 VSS.n1002 VSS.n1001 0.012
R31930 VSS.n1069 VSS.n1068 0.012
R31931 VSS.n1060 VSS.n1059 0.012
R31932 VSS.n1053 VSS.n1005 0.012
R31933 VSS.n1047 VSS.n1011 0.012
R31934 VSS.n1041 VSS.n1015 0.012
R31935 VSS.n1035 VSS.n1019 0.012
R31936 VSS.n1030 VSS.n1022 0.012
R31937 VSS.n1025 VSS.n185 0.012
R31938 VSS.n1092 VSS.n1091 0.012
R31939 VSS.n1159 VSS.n1158 0.012
R31940 VSS.n1150 VSS.n1149 0.012
R31941 VSS.n1143 VSS.n1095 0.012
R31942 VSS.n1137 VSS.n1101 0.012
R31943 VSS.n1131 VSS.n1105 0.012
R31944 VSS.n1125 VSS.n1109 0.012
R31945 VSS.n1120 VSS.n1112 0.012
R31946 VSS.n1115 VSS.n95 0.012
R31947 VSS.n1182 VSS.n1181 0.012
R31948 VSS.n1244 VSS.n1243 0.012
R31949 VSS.n1235 VSS.n1234 0.012
R31950 VSS.n1228 VSS.n1185 0.012
R31951 VSS.n1222 VSS.n1191 0.012
R31952 VSS.n1216 VSS.n1195 0.012
R31953 VSS.n1210 VSS.n1199 0.012
R31954 VSS.n1205 VSS.n1202 0.012
R31955 VSS.n1259 VSS.n1258 0.012
R31956 VSS.n1260 VSS.n2 0.012
R31957 VSS.n1265 VSS.n1264 0.012
R31958 VSS.n3050 VSS.n3049 0.012
R31959 VSS.n17593 VSS.n17592 0.011
R31960 VSS.n17589 VSS.n17588 0.011
R31961 VSS.n17585 VSS.n17584 0.011
R31962 VSS.n3065 VSS.n3064 0.011
R31963 VSS.n3069 VSS.n3068 0.011
R31964 VSS.n3073 VSS.n3072 0.011
R31965 VSS.n3092 VSS.n3091 0.011
R31966 VSS.n3096 VSS.n3095 0.011
R31967 VSS.n3100 VSS.n3099 0.011
R31968 VSS.n6615 VSS.n6614 0.011
R31969 VSS.n6619 VSS.n6618 0.011
R31970 VSS.n6623 VSS.n6622 0.011
R31971 VSS.n10380 VSS.n10379 0.011
R31972 VSS.n10384 VSS.n10383 0.011
R31973 VSS.n10388 VSS.n10387 0.011
R31974 VSS.n13973 VSS.n13972 0.011
R31975 VSS.n13977 VSS.n13976 0.011
R31976 VSS.n13981 VSS.n13980 0.011
R31977 VSS.n17493 VSS.n17492 0.011
R31978 VSS.n17497 VSS.n17496 0.011
R31979 VSS.n17501 VSS.n17500 0.011
R31980 VSS.n17533 VSS.n17532 0.011
R31981 VSS.n17537 VSS.n17536 0.011
R31982 VSS.n17541 VSS.n17540 0.011
R31983 VSS.n17711 VSS.n17639 0.011
R31984 VSS.n17637 VSS.n17635 0.011
R31985 VSS.n17633 VSS.n17631 0.011
R31986 VSS.n10415 VSS.n10414 0.011
R31987 VSS.n3131 VSS.n3113 0.011
R31988 VSS.n17484 VSS.n13994 0.01
R31989 VSS.n17530 VSS.n17529 0.01
R31990 VSS.n17490 VSS.n17489 0.01
R31991 VSS.n13970 VSS.n13969 0.01
R31992 VSS.n10377 VSS.n10376 0.01
R31993 VSS.n6612 VSS.n6611 0.01
R31994 VSS.n3089 VSS.n3088 0.01
R31995 VSS.n3062 VSS.n3061 0.01
R31996 VSS.n17596 VSS.n17595 0.01
R31997 VSS.n13963 VSS.n10400 0.01
R31998 VSS.n10446 VSS.n10441 0.01
R31999 VSS.n10471 VSS.n10423 0.01
R32000 VSS.n17674 VSS.n17652 0.01
R32001 VSS.n17689 VSS.n17688 0.01
R32002 VSS.n17575 VSS.n17573 0.009
R32003 VSS.n17571 VSS.n17570 0.009
R32004 VSS.n17568 VSS.n17567 0.009
R32005 VSS.n17565 VSS.n17564 0.009
R32006 VSS.n17562 VSS.n17561 0.009
R32007 VSS.n17559 VSS.n17558 0.009
R32008 VSS.n17556 VSS.n17555 0.009
R32009 VSS.n17553 VSS.n17552 0.009
R32010 VSS.n13963 VSS.n13962 0.009
R32011 VSS.n17540 VSS.n17539 0.009
R32012 VSS.n17536 VSS.n17535 0.009
R32013 VSS.n17532 VSS.n17531 0.009
R32014 VSS.n17500 VSS.n17499 0.009
R32015 VSS.n17496 VSS.n17495 0.009
R32016 VSS.n17492 VSS.n17491 0.009
R32017 VSS.n13980 VSS.n13979 0.009
R32018 VSS.n13976 VSS.n13975 0.009
R32019 VSS.n13972 VSS.n13971 0.009
R32020 VSS.n10387 VSS.n10386 0.009
R32021 VSS.n10383 VSS.n10382 0.009
R32022 VSS.n10379 VSS.n10378 0.009
R32023 VSS.n6622 VSS.n6621 0.009
R32024 VSS.n6618 VSS.n6617 0.009
R32025 VSS.n6614 VSS.n6613 0.009
R32026 VSS.n3099 VSS.n3098 0.009
R32027 VSS.n3095 VSS.n3094 0.009
R32028 VSS.n3091 VSS.n3090 0.009
R32029 VSS.n3072 VSS.n3071 0.009
R32030 VSS.n3068 VSS.n3067 0.009
R32031 VSS.n3064 VSS.n3063 0.009
R32032 VSS.n17586 VSS.n17585 0.009
R32033 VSS.n17590 VSS.n17589 0.009
R32034 VSS.n17594 VSS.n17593 0.009
R32035 VSS.n17633 VSS.n17632 0.009
R32036 VSS.n17637 VSS.n17636 0.009
R32037 VSS.n17711 VSS.n17710 0.009
R32038 VSS.n3130 VSS.n3129 0.008
R32039 VSS.n3126 VSS.n3125 0.007
R32040 VSS.n10402 VSS.n10401 0.007
R32041 VSS.n17546 VSS.n17545 0.007
R32042 VSS.n17544 VSS.n17543 0.007
R32043 VSS.n17506 VSS.n17505 0.007
R32044 VSS.n17504 VSS.n17503 0.007
R32045 VSS.n13986 VSS.n13985 0.007
R32046 VSS.n13984 VSS.n13983 0.007
R32047 VSS.n10393 VSS.n10392 0.007
R32048 VSS.n10391 VSS.n10390 0.007
R32049 VSS.n6628 VSS.n6627 0.007
R32050 VSS.n6626 VSS.n6625 0.007
R32051 VSS.n3105 VSS.n3104 0.007
R32052 VSS.n3103 VSS.n3102 0.007
R32053 VSS.n3078 VSS.n3077 0.007
R32054 VSS.n3076 VSS.n3075 0.007
R32055 VSS.n17580 VSS.n17579 0.007
R32056 VSS.n17582 VSS.n17581 0.007
R32057 VSS.n17614 VSS.n17613 0.007
R32058 VSS.n17629 VSS.n17628 0.007
R32059 VSS.n17709 VSS.n17708 0.007
R32060 VSS.n17542 VSS.n17541 0.007
R32061 VSS.n17538 VSS.n17537 0.007
R32062 VSS.n17534 VSS.n17533 0.007
R32063 VSS.n17502 VSS.n17501 0.007
R32064 VSS.n17498 VSS.n17497 0.007
R32065 VSS.n17494 VSS.n17493 0.007
R32066 VSS.n13982 VSS.n13981 0.007
R32067 VSS.n13978 VSS.n13977 0.007
R32068 VSS.n13974 VSS.n13973 0.007
R32069 VSS.n10389 VSS.n10388 0.007
R32070 VSS.n10385 VSS.n10384 0.007
R32071 VSS.n10381 VSS.n10380 0.007
R32072 VSS.n6624 VSS.n6623 0.007
R32073 VSS.n6620 VSS.n6619 0.007
R32074 VSS.n6616 VSS.n6615 0.007
R32075 VSS.n3101 VSS.n3100 0.007
R32076 VSS.n3097 VSS.n3096 0.007
R32077 VSS.n3093 VSS.n3092 0.007
R32078 VSS.n3074 VSS.n3073 0.007
R32079 VSS.n3070 VSS.n3069 0.007
R32080 VSS.n3066 VSS.n3065 0.007
R32081 VSS.n17584 VSS.n17583 0.007
R32082 VSS.n17588 VSS.n17587 0.007
R32083 VSS.n17592 VSS.n17591 0.007
R32084 VSS.n17603 VSS.n17602 0.007
R32085 VSS.n17622 VSS.n17621 0.007
R32086 VSS.n17617 VSS.n17616 0.007
R32087 VSS.n17631 VSS.n17630 0.007
R32088 VSS.n17635 VSS.n17634 0.007
R32089 VSS.n17639 VSS.n17638 0.007
R32090 VSS.n17707 VSS.n17706 0.006
R32091 VSS.n17575 VSS.n17574 0.005
R32092 VSS.n17572 VSS.n17571 0.005
R32093 VSS.n17569 VSS.n17568 0.005
R32094 VSS.n17566 VSS.n17565 0.005
R32095 VSS.n17563 VSS.n17562 0.005
R32096 VSS.n17560 VSS.n17559 0.005
R32097 VSS.n17557 VSS.n17556 0.005
R32098 VSS.n17554 VSS.n17553 0.005
R32099 VSS.n10442 VSS.n10427 0.005
R32100 VSS.n10466 VSS.n10425 0.005
R32101 VSS.n17676 VSS.n17649 0.005
R32102 VSS.n17683 VSS.n17682 0.005
R32103 VSS.n10416 VSS.n10402 0.004
R32104 VSS.n17418 VSS.n16024 0.003
R32105 VSS.n3133 VSS.n3132 0.002
R32106 VSS.n17468 VSS.n13994 0.002
R32107 VSS.n6896 VSS.n6883 0.002
R32108 VSS.n17609 VSS.n17608 0.001
R32109 VSS.n3130 VSS.n3114 0.001
R32110 VSS.n6605 VSS.n3136 0.001
R32111 VSS.n3049 sky130_asc_pnp_05v5_W3p40L3p40_7_0/Base 0.001
R32112 VSS.n17712 VSS.n17609 0.001
R32113 VSS.n3125 VSS.n3124 0.001
R32114 VSS.n17545 VSS.n17511 0.001
R32115 VSS.n17527 VSS.n17526 0.001
R32116 VSS.n17547 VSS.n17510 0.001
R32117 VSS.n17505 VSS.n13991 0.001
R32118 VSS.n17487 VSS.n17486 0.001
R32119 VSS.n17507 VSS.n13990 0.001
R32120 VSS.n13985 VSS.n10398 0.001
R32121 VSS.n13967 VSS.n13966 0.001
R32122 VSS.n13987 VSS.n10397 0.001
R32123 VSS.n10392 VSS.n6633 0.001
R32124 VSS.n10374 VSS.n10373 0.001
R32125 VSS.n10394 VSS.n6632 0.001
R32126 VSS.n6627 VSS.n3110 0.001
R32127 VSS.n6609 VSS.n6608 0.001
R32128 VSS.n6629 VSS.n3109 0.001
R32129 VSS.n3104 VSS.n3083 0.001
R32130 VSS.n3086 VSS.n3085 0.001
R32131 VSS.n3106 VSS.n3082 0.001
R32132 VSS.n3077 VSS.n3056 0.001
R32133 VSS.n3059 VSS.n3058 0.001
R32134 VSS.n3079 VSS.n3055 0.001
R32135 VSS.n17580 VSS.n3053 0.001
R32136 VSS.n17599 VSS.n17598 0.001
R32137 VSS.n17578 VSS.n3054 0.001
R32138 VSS.n17627 VSS.n17626 0.001
R32139 VSS.n17706 VSS.n17705 0.001
R32140 VSS.n17613 VSS.n17611 0.001
R32141 VSS.t30 VSS.n16035 0.001
R32142 VSS.n17460 VSS.n16035 0.001
R32143 VSS.n17305 VSS.n16074 0.001
R32144 VSS.t54 VSS.n16074 0.001
R32145 VSS.n17215 VSS.n16164 0.001
R32146 VSS.t50 VSS.n16164 0.001
R32147 VSS.n17125 VSS.n16254 0.001
R32148 VSS.t42 VSS.n16254 0.001
R32149 VSS.n17035 VSS.n16344 0.001
R32150 VSS.t68 VSS.n16344 0.001
R32151 VSS.n16945 VSS.n16434 0.001
R32152 VSS.t74 VSS.n16434 0.001
R32153 VSS.n16855 VSS.n16524 0.001
R32154 VSS.t90 VSS.n16524 0.001
R32155 VSS.n16765 VSS.n16614 0.001
R32156 VSS.t28 VSS.n16614 0.001
R32157 VSS.n11232 VSS.n11081 0.001
R32158 VSS.t58 VSS.n11081 0.001
R32159 VSS.n11322 VSS.n10991 0.001
R32160 VSS.t32 VSS.n10991 0.001
R32161 VSS.n11412 VSS.n10901 0.001
R32162 VSS.t92 VSS.n10901 0.001
R32163 VSS.n13532 VSS.n10811 0.001
R32164 VSS.t88 VSS.n10811 0.001
R32165 VSS.n13622 VSS.n10721 0.001
R32166 VSS.t72 VSS.n10721 0.001
R32167 VSS.n13712 VSS.n10631 0.001
R32168 VSS.t78 VSS.n10631 0.001
R32169 VSS.n13802 VSS.n10541 0.001
R32170 VSS.t82 VSS.n10541 0.001
R32171 VSS.t62 VSS.n10496 0.001
R32172 VSS.n13952 VSS.n10496 0.001
R32173 VSS.n10260 VSS.n9209 0.001
R32174 VSS.t34 VSS.n9209 0.001
R32175 VSS.n10170 VSS.n9299 0.001
R32176 VSS.t26 VSS.n9299 0.001
R32177 VSS.n10080 VSS.n9389 0.001
R32178 VSS.t52 VSS.n9389 0.001
R32179 VSS.n9990 VSS.n9479 0.001
R32180 VSS.t56 VSS.n9479 0.001
R32181 VSS.n9900 VSS.n9569 0.001
R32182 VSS.t80 VSS.n9569 0.001
R32183 VSS.n9810 VSS.n9659 0.001
R32184 VSS.t18 VSS.n9659 0.001
R32185 VSS.n9178 VSS.n8935 0.001
R32186 VSS.t38 VSS.n9178 0.001
R32187 VSS.n5733 VSS.n3582 0.001
R32188 VSS.t46 VSS.n5733 0.001
R32189 VSS.n5855 VSS.n3524 0.001
R32190 VSS.t70 VSS.n5855 0.001
R32191 VSS.n5977 VSS.n3466 0.001
R32192 VSS.t66 VSS.n5977 0.001
R32193 VSS.n6099 VSS.n3408 0.001
R32194 VSS.t64 VSS.n6099 0.001
R32195 VSS.n6221 VSS.n3350 0.001
R32196 VSS.t84 VSS.n6221 0.001
R32197 VSS.n6343 VSS.n3292 0.001
R32198 VSS.t86 VSS.n6343 0.001
R32199 VSS.n6465 VSS.n3234 0.001
R32200 VSS.t24 VSS.n6465 0.001
R32201 VSS.n6598 VSS.n3145 0.001
R32202 VSS.n3145 VSS.t44 0.001
R32203 VSS.n1252 VSS.n26 0.001
R32204 VSS.t60 VSS.n26 0.001
R32205 VSS.n1168 VSS.n117 0.001
R32206 VSS.t48 VSS.n117 0.001
R32207 VSS.n1078 VSS.n207 0.001
R32208 VSS.t76 VSS.n207 0.001
R32209 VSS.n988 VSS.n297 0.001
R32210 VSS.t22 VSS.n297 0.001
R32211 VSS.n898 VSS.n387 0.001
R32212 VSS.t16 VSS.n387 0.001
R32213 VSS.n808 VSS.n477 0.001
R32214 VSS.t36 VSS.n477 0.001
R32215 VSS.n718 VSS.n567 0.001
R32216 VSS.t40 VSS.n567 0.001
R32217 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n54 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t14 247.724
R32218 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n24 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t67 212.91
R32219 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n85 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n84 195.413
R32220 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n84 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n83 195.413
R32221 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n83 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n82 195.413
R32222 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n82 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n80 195.413
R32223 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n80 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n79 195.413
R32224 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n79 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n78 195.413
R32225 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n78 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n77 195.413
R32226 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n77 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n76 195.413
R32227 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n76 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n75 195.413
R32228 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n75 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n74 195.413
R32229 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n74 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n73 195.413
R32230 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n73 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n72 195.413
R32231 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n72 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n71 195.413
R32232 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n71 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n70 195.413
R32233 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n70 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n69 195.413
R32234 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n69 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n68 195.413
R32235 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n66 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n65 195.413
R32236 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n65 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n64 195.413
R32237 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n64 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n63 195.413
R32238 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n63 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n62 195.413
R32239 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n62 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n61 195.413
R32240 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n61 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n60 195.413
R32241 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n60 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n59 195.413
R32242 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n59 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n58 195.413
R32243 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n58 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n57 195.413
R32244 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n57 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n56 195.413
R32245 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n56 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n55 195.413
R32246 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n55 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n54 195.413
R32247 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n19 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t68 180.68
R32248 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n67 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n66 168.533
R32249 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n33 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t65 154.653
R32250 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n30 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t64 154.653
R32251 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n22 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t66 154.653
R32252 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n27 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t63 154.653
R32253 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n21 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t69 154.653
R32254 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n23 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t62 154.653
R32255 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n20 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t70 154.653
R32256 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n26 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n24 118.858
R32257 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n39 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n38 85.333
R32258 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n38 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n37 85.333
R32259 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n37 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n36 85.333
R32260 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n36 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n35 85.333
R32261 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n35 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n32 85.333
R32262 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n32 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n29 85.333
R32263 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n29 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n26 85.333
R32264 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n28 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n27 78.084
R32265 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n39 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n19 76
R32266 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n38 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n20 76
R32267 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n37 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n21 76
R32268 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n36 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n22 76
R32269 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n35 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n34 76
R32270 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n32 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n31 76
R32271 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n29 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n28 76
R32272 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n26 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n25 76
R32273 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n67 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n40 57.196
R32274 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n24 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n23 56.845
R32275 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n85 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t48 52.312
R32276 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n31 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n30 51.092
R32277 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n84 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n0 47.884
R32278 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n80 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n6 47.884
R32279 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n79 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n7 47.884
R32280 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n78 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n8 47.884
R32281 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n77 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n9 47.884
R32282 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n76 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n10 47.884
R32283 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n75 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n11 47.884
R32284 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n74 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n12 47.884
R32285 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n73 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n13 47.884
R32286 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n72 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n14 47.884
R32287 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n71 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n15 47.884
R32288 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n70 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n16 47.884
R32289 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n69 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n17 47.884
R32290 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n68 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n18 47.884
R32291 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n66 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n41 47.884
R32292 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n65 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n42 47.884
R32293 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n64 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n43 47.884
R32294 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n63 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n44 47.884
R32295 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n62 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n45 47.884
R32296 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n61 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n46 47.884
R32297 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n60 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n47 47.884
R32298 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n59 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n48 47.884
R32299 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n58 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n49 47.884
R32300 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n57 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n50 47.884
R32301 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n56 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n51 47.884
R32302 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n55 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n52 47.884
R32303 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n54 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n53 47.884
R32304 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n82 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n81 47.882
R32305 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n83 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n5 46.86
R32306 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n40 sky130_asc_nfet_01v8_lvt_9_2/GATE 37.973
R32307 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n40 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n39 30.293
R32308 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n68 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n67 26.88
R32309 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n34 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n33 24.1
R32310 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n5 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n3 16.93
R32311 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n3 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n2 11.022
R32312 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n2 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t61 4.85
R32313 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n1 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t0 4.85
R32314 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n0 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t20 4.428
R32315 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n0 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t32 4.428
R32316 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n4 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t58 4.428
R32317 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n4 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t59 4.428
R32318 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n6 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t54 4.428
R32319 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n6 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t55 4.428
R32320 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n7 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t56 4.428
R32321 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n7 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t57 4.428
R32322 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n8 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t43 4.428
R32323 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n8 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t44 4.428
R32324 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n9 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t26 4.428
R32325 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n9 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t46 4.428
R32326 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n10 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t53 4.428
R32327 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n10 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t29 4.428
R32328 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n11 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t40 4.428
R32329 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n11 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t19 4.428
R32330 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n12 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t41 4.428
R32331 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n12 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t22 4.428
R32332 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n13 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t23 4.428
R32333 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n13 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t34 4.428
R32334 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n14 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t2 4.428
R32335 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n14 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t36 4.428
R32336 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n15 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t42 4.428
R32337 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n15 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t50 4.428
R32338 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n16 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t51 4.428
R32339 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n16 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t35 4.428
R32340 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n17 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t52 4.428
R32341 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n17 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t38 4.428
R32342 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n18 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t45 4.428
R32343 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n18 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t16 4.428
R32344 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n41 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t27 4.428
R32345 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n41 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t47 4.428
R32346 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n42 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t30 4.428
R32347 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n42 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t31 4.428
R32348 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n43 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t8 4.428
R32349 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n43 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t9 4.428
R32350 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n44 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t12 4.428
R32351 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n44 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t13 4.428
R32352 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n45 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t24 4.428
R32353 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n45 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t3 4.428
R32354 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n46 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t4 4.428
R32355 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n46 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t5 4.428
R32356 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n47 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t6 4.428
R32357 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n47 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t15 4.428
R32358 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n48 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t25 4.428
R32359 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n48 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t37 4.428
R32360 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n49 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t28 4.428
R32361 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n49 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t39 4.428
R32362 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n50 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t7 4.428
R32363 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n50 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t17 4.428
R32364 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n51 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t18 4.428
R32365 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n51 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t21 4.428
R32366 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n52 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t33 4.428
R32367 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n52 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t1 4.428
R32368 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n53 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t10 4.428
R32369 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n53 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t11 4.428
R32370 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n81 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t60 4.428
R32371 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n81 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t49 4.428
R32372 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n5 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n4 1.024
R32373 sky130_asc_pfet_01v8_lvt_60_1/DRAIN sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n85 0.853
R32374 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n3 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n1 0.38
R32375 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n2 sky130_asc_res_xhigh_po_2p85_1_20/Rin 0.018
R32376 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n1 sky130_asc_res_xhigh_po_2p85_1_18/Rin 0.018
R32377 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n6 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n5 321.976
R32378 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n14 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n13 321.976
R32379 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n8 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n7 195.413
R32380 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n7 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n6 195.413
R32381 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n15 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n14 195.413
R32382 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n16 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n15 189.16
R32383 sky130_asc_nfet_01v8_lvt_9_1/SOURCE sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n17 188.733
R32384 sky130_asc_nfet_01v8_lvt_9_1/SOURCE sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t8 137.314
R32385 sky130_asc_nfet_01v8_lvt_9_2/SOURCE sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t15 137.313
R32386 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n9 sky130_asc_nfet_01v8_lvt_9_2/SOURCE 136.106
R32387 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n6 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n4 126.563
R32388 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n7 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n3 126.563
R32389 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n8 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n2 126.563
R32390 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n14 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n12 126.563
R32391 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n15 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n11 126.563
R32392 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n17 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n0 124.681
R32393 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n1 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t18 119.662
R32394 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n1 sky130_asc_nfet_01v8_lvt_1_1/DRAIN 85.76
R32395 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n10 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n1 60.656
R32396 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n9 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n8 52.906
R32397 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n10 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n9 21.029
R32398 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n16 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n10 7.192
R32399 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n17 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n16 5.513
R32400 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n5 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t14 4.35
R32401 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n5 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t10 4.35
R32402 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n4 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t12 4.35
R32403 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n4 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t13 4.35
R32404 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n3 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t9 4.35
R32405 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n3 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t11 4.35
R32406 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n2 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t17 4.35
R32407 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n2 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t16 4.35
R32408 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n13 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t5 4.35
R32409 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n13 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t0 4.35
R32410 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n12 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t3 4.35
R32411 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n12 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t4 4.35
R32412 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n11 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t1 4.35
R32413 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n11 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t2 4.35
R32414 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n0 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t6 4.35
R32415 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n0 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t7 4.35
R32416 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n47 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t3 243.258
R32417 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n54 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n53 242.276
R32418 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n28 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t23 222.22
R32419 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n49 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n48 195.413
R32420 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n48 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n47 195.413
R32421 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n56 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n55 195.413
R32422 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n55 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n54 195.413
R32423 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n50 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n49 170.24
R32424 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n26 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t21 166.1
R32425 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n4 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t15 166.1
R32426 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n35 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t26 166.1
R32427 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n9 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t9 166.1
R32428 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n2 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t13 166.1
R32429 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n32 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t25 166.1
R32430 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n12 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t17 166.1
R32431 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n29 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t24 166.1
R32432 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n15 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t19 166.1
R32433 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n18 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t11 166.099
R32434 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n24 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t22 164.092
R32435 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n31 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n28 122.204
R32436 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n10 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n9 100.256
R32437 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n19 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n18 95.28
R32438 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n43 sky130_asc_nfet_01v8_lvt_9_2/DRAIN 91.306
R32439 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n30 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n29 88.688
R32440 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n38 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n37 85.333
R32441 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n37 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n34 85.333
R32442 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n34 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n31 85.333
R32443 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n6 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n3 85.333
R32444 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n8 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n6 85.333
R32445 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n11 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n8 85.333
R32446 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n14 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n11 85.333
R32447 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n17 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n14 85.333
R32448 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n19 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n17 85.333
R32449 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n39 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n38 81.066
R32450 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n38 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n27 76
R32451 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n37 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n36 76
R32452 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n34 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n33 76
R32453 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n31 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n30 76
R32454 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n3 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n2 76
R32455 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n6 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n5 76
R32456 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n8 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n7 76
R32457 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n11 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n10 76
R32458 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n14 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n13 76
R32459 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n17 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n16 76
R32460 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n13 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n12 73.264
R32461 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n52 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n51 66.158
R32462 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n33 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n32 61.696
R32463 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n56 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t14 52.311
R32464 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n55 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n0 47.884
R32465 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n54 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n1 47.884
R32466 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n16 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n15 46.272
R32467 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n3 sky130_asc_pfet_01v8_lvt_6_1/GATE 46.08
R32468 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n43 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n42 43.495
R32469 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n49 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n44 43.495
R32470 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n48 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n45 43.495
R32471 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n47 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n46 43.495
R32472 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n21 sky130_asc_pfet_01v8_lvt_6_0/GATE 43.093
R32473 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n52 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n19 40.473
R32474 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n36 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n35 34.704
R32475 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n50 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n43 25.173
R32476 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n51 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n41 18.097
R32477 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n25 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n24 9.3
R32478 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n27 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n26 7.712
R32479 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n5 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n4 7.712
R32480 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n53 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t12 5.448
R32481 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n0 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t16 4.428
R32482 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n0 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t10 4.428
R32483 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n1 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t18 4.428
R32484 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n1 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t20 4.428
R32485 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n42 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t2 4.35
R32486 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n42 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t0 4.35
R32487 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n44 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t1 4.35
R32488 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n44 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t4 4.35
R32489 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n45 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t5 4.35
R32490 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n45 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t6 4.35
R32491 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n46 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t7 4.35
R32492 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n46 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t8 4.35
R32493 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n41 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n40 3.774
R32494 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n51 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n50 3.772
R32495 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n53 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n52 3.054
R32496 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n22 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n21 2.986
R32497 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n40 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n39 2.986
R32498 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n24 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n23 2.008
R32499 sky130_asc_pfet_01v8_lvt_6_1/DRAIN sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n56 0.853
R32500 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n25 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n22 0.64
R32501 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n40 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n25 0.64
R32502 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n41 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n20 0.039
R32503 vbg.n29 vbg.t1 247.724
R32504 vbg.n175 vbg.n174 195.413
R32505 vbg.n174 vbg.n173 195.413
R32506 vbg.n173 vbg.n172 195.413
R32507 vbg.n172 vbg.n171 195.413
R32508 vbg.n169 vbg.n168 195.413
R32509 vbg.n168 vbg.n167 195.413
R32510 vbg.n167 vbg.n166 195.413
R32511 vbg.n166 vbg.n165 195.413
R32512 vbg.n165 vbg.n164 195.413
R32513 vbg.n164 vbg.n163 195.413
R32514 vbg.n163 vbg.n162 195.413
R32515 vbg.n162 vbg.n161 195.413
R32516 vbg.n161 vbg.n160 195.413
R32517 vbg.n160 vbg.n159 195.413
R32518 vbg.n159 vbg.n158 195.413
R32519 vbg.n158 vbg.n157 195.413
R32520 vbg.n157 vbg.n40 195.413
R32521 vbg.n40 vbg.n39 195.413
R32522 vbg.n39 vbg.n38 195.413
R32523 vbg.n38 vbg.n37 195.413
R32524 vbg.n37 vbg.n36 195.413
R32525 vbg.n36 vbg.n35 195.413
R32526 vbg.n35 vbg.n34 195.413
R32527 vbg.n34 vbg.n33 195.413
R32528 vbg.n33 vbg.n32 195.413
R32529 vbg.n32 vbg.n31 195.413
R32530 vbg.n31 vbg.n30 195.413
R32531 vbg.n30 vbg.n29 195.413
R32532 vbg.n170 vbg.n169 147.626
R32533 vbg.n170 vbg.n4 88.562
R32534 vbg.n175 vbg.t42 52.312
R32535 vbg.n174 vbg.n0 47.884
R32536 vbg.n173 vbg.n1 47.884
R32537 vbg.n172 vbg.n2 47.884
R32538 vbg.n171 vbg.n3 47.884
R32539 vbg.n169 vbg.n5 47.884
R32540 vbg.n168 vbg.n6 47.884
R32541 vbg.n167 vbg.n7 47.884
R32542 vbg.n166 vbg.n8 47.884
R32543 vbg.n165 vbg.n9 47.884
R32544 vbg.n164 vbg.n10 47.884
R32545 vbg.n163 vbg.n11 47.884
R32546 vbg.n162 vbg.n12 47.884
R32547 vbg.n161 vbg.n13 47.884
R32548 vbg.n160 vbg.n14 47.884
R32549 vbg.n159 vbg.n15 47.884
R32550 vbg.n158 vbg.n16 47.884
R32551 vbg.n40 vbg.n17 47.884
R32552 vbg.n39 vbg.n18 47.884
R32553 vbg.n38 vbg.n19 47.884
R32554 vbg.n37 vbg.n20 47.884
R32555 vbg.n36 vbg.n21 47.884
R32556 vbg.n35 vbg.n22 47.884
R32557 vbg.n34 vbg.n23 47.884
R32558 vbg.n33 vbg.n24 47.884
R32559 vbg.n32 vbg.n25 47.884
R32560 vbg.n31 vbg.n26 47.884
R32561 vbg.n30 vbg.n27 47.884
R32562 vbg.n29 vbg.n28 47.884
R32563 vbg.n171 vbg.n170 47.786
R32564 vbg.n157 vbg.n156 44.423
R32565 vbg.n58 vbg 30.4
R32566 vbg.n103 vbg.n102 13.176
R32567 vbg.n148 vbg.n147 9.3
R32568 vbg.n141 vbg.n140 9.3
R32569 vbg.n134 vbg.n133 9.3
R32570 vbg.n127 vbg.n126 9.3
R32571 vbg.n120 vbg.n119 9.3
R32572 vbg.n113 vbg.n112 9.3
R32573 vbg.n106 vbg.n105 9.3
R32574 vbg.n99 vbg.n98 9.3
R32575 vbg.n92 vbg.n91 9.3
R32576 vbg.n86 vbg.n85 9.3
R32577 vbg.n80 vbg.n79 9.3
R32578 vbg.n75 vbg.n74 9.3
R32579 vbg.n70 vbg.n69 9.3
R32580 vbg.n65 vbg.n64 9.3
R32581 vbg.n62 vbg.n61 9.3
R32582 vbg.n67 vbg.n66 9.3
R32583 vbg.n72 vbg.n71 9.3
R32584 vbg.n77 vbg.n76 9.3
R32585 vbg.n82 vbg.n81 9.3
R32586 vbg.n84 vbg.n83 9.3
R32587 vbg.n88 vbg.n87 9.3
R32588 vbg.n90 vbg.n89 9.3
R32589 vbg.n94 vbg.n93 9.3
R32590 vbg.n97 vbg.n96 9.3
R32591 vbg.n101 vbg.n100 9.3
R32592 vbg.n104 vbg.n103 9.3
R32593 vbg.n109 vbg.n108 9.3
R32594 vbg.n111 vbg.n110 9.3
R32595 vbg.n116 vbg.n115 9.3
R32596 vbg.n118 vbg.n117 9.3
R32597 vbg.n123 vbg.n122 9.3
R32598 vbg.n125 vbg.n124 9.3
R32599 vbg.n130 vbg.n129 9.3
R32600 vbg.n132 vbg.n131 9.3
R32601 vbg.n137 vbg.n136 9.3
R32602 vbg.n139 vbg.n138 9.3
R32603 vbg.n144 vbg.n143 9.3
R32604 vbg.n146 vbg.n145 9.3
R32605 vbg.n151 vbg.n150 9.3
R32606 vbg.n153 vbg.n152 9.3
R32607 vbg.n56 vbg.n52 8.897
R32608 vbg.n56 vbg.n50 8.886
R32609 vbg.n56 vbg.n48 8.875
R32610 vbg.n56 vbg.n46 8.864
R32611 vbg.n56 vbg.n44 8.854
R32612 vbg.n56 vbg.n43 8.843
R32613 vbg.n156 vbg.n57 5.418
R32614 vbg.n55 vbg.n54 5.38
R32615 vbg.n57 vbg.n42 5.38
R32616 vbg.n4 vbg.t60 4.85
R32617 vbg.n156 vbg.n155 4.84
R32618 vbg.n56 vbg.t40 4.428
R32619 vbg.n56 vbg.t41 4.428
R32620 vbg.n0 vbg.t43 4.428
R32621 vbg.n0 vbg.t17 4.428
R32622 vbg.n1 vbg.t45 4.428
R32623 vbg.n1 vbg.t22 4.428
R32624 vbg.n2 vbg.t52 4.428
R32625 vbg.n2 vbg.t55 4.428
R32626 vbg.n3 vbg.t44 4.428
R32627 vbg.n3 vbg.t57 4.428
R32628 vbg.n5 vbg.t50 4.428
R32629 vbg.n5 vbg.t51 4.428
R32630 vbg.n6 vbg.t36 4.428
R32631 vbg.n6 vbg.t37 4.428
R32632 vbg.n7 vbg.t54 4.428
R32633 vbg.n7 vbg.t39 4.428
R32634 vbg.n8 vbg.t49 4.428
R32635 vbg.n8 vbg.t14 4.428
R32636 vbg.n9 vbg.t30 4.428
R32637 vbg.n9 vbg.t18 4.428
R32638 vbg.n10 vbg.t33 4.428
R32639 vbg.n10 vbg.t34 4.428
R32640 vbg.n11 vbg.t8 4.428
R32641 vbg.n11 vbg.t20 4.428
R32642 vbg.n12 vbg.t10 4.428
R32643 vbg.n12 vbg.t24 4.428
R32644 vbg.n13 vbg.t25 4.428
R32645 vbg.n13 vbg.t2 4.428
R32646 vbg.n14 vbg.t46 4.428
R32647 vbg.n14 vbg.t47 4.428
R32648 vbg.n15 vbg.t48 4.428
R32649 vbg.n15 vbg.t26 4.428
R32650 vbg.n16 vbg.t27 4.428
R32651 vbg.n16 vbg.t38 4.428
R32652 vbg.n17 vbg.t15 4.428
R32653 vbg.n17 vbg.t16 4.428
R32654 vbg.n18 vbg.t31 4.428
R32655 vbg.n18 vbg.t21 4.428
R32656 vbg.n19 vbg.t35 4.428
R32657 vbg.n19 vbg.t0 4.428
R32658 vbg.n20 vbg.t9 4.428
R32659 vbg.n20 vbg.t56 4.428
R32660 vbg.n21 vbg.t11 4.428
R32661 vbg.n21 vbg.t12 4.428
R32662 vbg.n22 vbg.t58 4.428
R32663 vbg.n22 vbg.t3 4.428
R32664 vbg.n23 vbg.t53 4.428
R32665 vbg.n23 vbg.t5 4.428
R32666 vbg.n24 vbg.t13 4.428
R32667 vbg.n24 vbg.t28 4.428
R32668 vbg.n25 vbg.t29 4.428
R32669 vbg.n25 vbg.t4 4.428
R32670 vbg.n26 vbg.t32 4.428
R32671 vbg.n26 vbg.t6 4.428
R32672 vbg.n27 vbg.t7 4.428
R32673 vbg.n27 vbg.t19 4.428
R32674 vbg.n28 vbg.t59 4.428
R32675 vbg.n28 vbg.t23 4.428
R32676 vbg.n57 vbg.n56 1.844
R32677 vbg.n56 vbg.n55 1.844
R32678 vbg vbg.n175 0.853
R32679 vbg.n54 vbg.n53 0.752
R32680 vbg.n42 vbg.n41 0.752
R32681 vbg.n59 vbg.n58 0.19
R32682 vbg.n104 vbg.n101 0.19
R32683 vbg.n96 vbg.n95 0.189
R32684 vbg.n108 vbg.n107 0.189
R32685 vbg.n115 vbg.n114 0.178
R32686 vbg.n122 vbg.n121 0.166
R32687 vbg.n46 vbg.n45 0.155
R32688 vbg.n129 vbg.n128 0.155
R32689 vbg.n48 vbg.n47 0.144
R32690 vbg.n136 vbg.n135 0.144
R32691 vbg.n63 vbg.n62 0.144
R32692 vbg.n68 vbg.n67 0.144
R32693 vbg.n73 vbg.n72 0.144
R32694 vbg.n78 vbg.n77 0.144
R32695 vbg.n84 vbg.n82 0.144
R32696 vbg.n90 vbg.n88 0.144
R32697 vbg.n97 vbg.n94 0.144
R32698 vbg.n111 vbg.n109 0.144
R32699 vbg.n118 vbg.n116 0.144
R32700 vbg.n125 vbg.n123 0.144
R32701 vbg.n132 vbg.n130 0.144
R32702 vbg.n139 vbg.n137 0.144
R32703 vbg.n146 vbg.n144 0.144
R32704 vbg.n153 vbg.n151 0.144
R32705 vbg.n50 vbg.n49 0.133
R32706 vbg.n143 vbg.n142 0.133
R32707 vbg.n52 vbg.n51 0.121
R32708 vbg.n150 vbg.n149 0.121
R32709 vbg.n99 vbg.n97 0.043
R32710 vbg.n109 vbg.n106 0.043
R32711 vbg.n62 vbg.n60 0.04
R32712 vbg.n154 vbg.n153 0.04
R32713 vbg.n92 vbg.n90 0.038
R32714 vbg.n116 vbg.n113 0.038
R32715 vbg.n67 vbg.n65 0.035
R32716 vbg.n148 vbg.n146 0.035
R32717 vbg.n86 vbg.n84 0.032
R32718 vbg.n123 vbg.n120 0.032
R32719 vbg.n72 vbg.n70 0.029
R32720 vbg.n141 vbg.n139 0.029
R32721 vbg.n80 vbg.n78 0.027
R32722 vbg.n130 vbg.n127 0.027
R32723 vbg.n77 vbg.n75 0.024
R32724 vbg.n134 vbg.n132 0.024
R32725 vbg.n75 vbg.n73 0.021
R32726 vbg.n137 vbg.n134 0.021
R32727 vbg.n82 vbg.n80 0.019
R32728 vbg.n127 vbg.n125 0.019
R32729 vbg.n4 sky130_asc_res_xhigh_po_2p85_1_8/Rin 0.018
R32730 vbg.n70 vbg.n68 0.016
R32731 vbg.n144 vbg.n141 0.016
R32732 vbg.n88 vbg.n86 0.013
R32733 vbg.n120 vbg.n118 0.013
R32734 vbg.n65 vbg.n63 0.01
R32735 vbg.n151 vbg.n148 0.01
R32736 vbg.n94 vbg.n92 0.008
R32737 vbg.n113 vbg.n111 0.008
R32738 vbg.n60 vbg.n59 0.005
R32739 vbg.n155 vbg.n154 0.005
R32740 vbg.n101 vbg.n99 0.002
R32741 vbg.n106 vbg.n104 0.002
R32742 sky130_asc_nfet_01v8_lvt_1_0/GATE sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t12 352.424
R32743 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n34 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t14 297.811
R32744 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n109 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n108 239.836
R32745 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n115 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n114 195.413
R32746 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n114 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n112 195.413
R32747 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n112 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n111 195.413
R32748 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n111 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n110 195.413
R32749 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n110 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n109 195.413
R32750 sky130_asc_nfet_01v8_lvt_1_0/DRAIN sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t13 176.798
R32751 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n35 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n34 103.039
R32752 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n34 sky130_asc_nfet_01v8_lvt_1_1/GATE 54.613
R32753 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n115 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t4 52.312
R32754 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n112 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n12 47.884
R32755 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n111 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n13 47.884
R32756 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n110 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n14 47.884
R32757 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n109 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n15 47.884
R32758 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n114 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n113 47.882
R32759 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n38 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n35 45.105
R32760 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n35 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n33 32.292
R32761 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n33 sky130_asc_nfet_01v8_lvt_1_0/DRAIN 15.217
R32762 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n33 sky130_asc_nfet_01v8_lvt_1_0/GATE 14.46
R32763 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n69 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n68 13.176
R32764 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n7 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n103 9.3
R32765 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n3 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n98 9.3
R32766 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n92 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n91 9.3
R32767 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n1 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n85 9.3
R32768 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n5 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n80 9.3
R32769 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n9 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n75 9.3
R32770 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n11 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n70 9.3
R32771 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n10 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n66 9.3
R32772 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n8 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n61 9.3
R32773 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n4 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n57 9.3
R32774 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n0 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n53 9.3
R32775 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n49 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n48 9.3
R32776 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n2 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n44 9.3
R32777 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n6 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n41 9.3
R32778 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n107 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n106 9.3
R32779 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n7 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n105 9.3
R32780 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n102 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n101 9.3
R32781 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n3 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n100 9.3
R32782 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n97 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n96 9.3
R32783 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n95 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n94 9.3
R32784 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n90 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n89 9.3
R32785 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n88 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n87 9.3
R32786 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n1 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n84 9.3
R32787 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n83 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n82 9.3
R32788 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n5 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n79 9.3
R32789 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n78 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n77 9.3
R32790 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n9 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n74 9.3
R32791 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n73 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n72 9.3
R32792 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n11 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n69 9.3
R32793 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n10 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n67 9.3
R32794 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n65 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n64 9.3
R32795 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n8 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n62 9.3
R32796 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n60 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n59 9.3
R32797 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n4 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n58 9.3
R32798 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n56 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n55 9.3
R32799 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n0 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n54 9.3
R32800 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n51 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n50 9.3
R32801 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n46 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n45 9.3
R32802 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n43 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n42 9.3
R32803 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n40 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n39 9.3
R32804 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n31 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n20 8.907
R32805 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n31 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n22 8.897
R32806 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n31 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n24 8.885
R32807 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n31 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n26 8.875
R32808 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n31 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n28 8.864
R32809 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n31 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n29 8.854
R32810 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n31 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n30 8.843
R32811 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n108 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n32 5.417
R32812 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n32 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n17 5.38
R32813 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n108 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n107 4.885
R32814 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n12 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t2 4.428
R32815 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n12 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t0 4.428
R32816 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n13 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t3 4.428
R32817 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n13 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t6 4.428
R32818 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n14 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t7 4.428
R32819 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n14 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t5 4.428
R32820 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n15 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t9 4.428
R32821 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n15 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t1 4.428
R32822 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n31 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t8 4.428
R32823 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n113 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t10 4.428
R32824 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n113 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t11 4.428
R32825 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n37 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n36 4.141
R32826 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n38 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n37 3.915
R32827 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n32 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n31 1.844
R32828 sky130_asc_pfet_01v8_lvt_12_1/DRAIN sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n115 0.853
R32829 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n19 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n18 0.752
R32830 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n17 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n16 0.752
R32831 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n11 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n10 0.19
R32832 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n64 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n63 0.189
R32833 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n72 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n71 0.189
R32834 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n77 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n76 0.177
R32835 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n82 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n81 0.166
R32836 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n87 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n86 0.155
R32837 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n28 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n27 0.155
R32838 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n26 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n25 0.144
R32839 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n94 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n93 0.144
R32840 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n6 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n40 0.144
R32841 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n2 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n43 0.144
R32842 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n47 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n46 0.144
R32843 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n52 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n51 0.144
R32844 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n56 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n0 0.144
R32845 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n60 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n4 0.144
R32846 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n65 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n8 0.144
R32847 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n9 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n73 0.144
R32848 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n5 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n78 0.144
R32849 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n1 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n83 0.144
R32850 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n90 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n88 0.144
R32851 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n97 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n95 0.144
R32852 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n102 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n3 0.144
R32853 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n107 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n7 0.144
R32854 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n100 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n99 0.132
R32855 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n24 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n23 0.132
R32856 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n22 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n21 0.121
R32857 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n105 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n104 0.121
R32858 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n20 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n19 0.109
R32859 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n73 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n11 0.045
R32860 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n10 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n65 0.045
R32861 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n51 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n49 0.024
R32862 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n92 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n90 0.024
R32863 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n49 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n47 0.021
R32864 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n95 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n92 0.021
R32865 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n40 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n38 0.224
R32866 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n78 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n9 0.046
R32867 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n8 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n60 0.046
R32868 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n88 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n1 0.046
R32869 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n0 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n52 0.046
R32870 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n7 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n102 0.045
R32871 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n43 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n6 0.045
R32872 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n83 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n5 0.045
R32873 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n4 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n56 0.045
R32874 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n3 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n97 0.045
R32875 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n46 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n2 0.045
R32876 sky130_asc_res_xhigh_po_2p85_1_21/Rout sky130_asc_res_xhigh_po_2p85_2_1/Rin 16.781
R32877 sky130_asc_res_xhigh_po_2p85_2_1/Rin sky130_asc_res_xhigh_po_2p85_1_21/Rout.t0 4.85
R32878 a_15392_9587.t0 a_15392_9587.t1 7.619
R32879 sky130_asc_res_xhigh_po_2p85_1_19/Rin sky130_asc_res_xhigh_po_2p85_1_20/Rout 49.324
R32880 sky130_asc_res_xhigh_po_2p85_1_20/Rout sky130_asc_res_xhigh_po_2p85_1_19/Rin.t0 4.85
R32881 a_39402_28387.t0 a_39402_28387.t1 7.619
R32882 sky130_asc_res_xhigh_po_2p85_1_17/Rout sky130_asc_res_xhigh_po_2p85_1_16/Rin 11.801
R32883 sky130_asc_res_xhigh_po_2p85_1_16/Rin sky130_asc_res_xhigh_po_2p85_1_17/Rout.t0 4.85
R32884 a_41264_17107.t0 a_41264_17107.t1 7.619
R32885 sky130_asc_res_xhigh_po_2p85_1_15/Rout sky130_asc_res_xhigh_po_2p85_1_14/Rin 38.745
R32886 sky130_asc_res_xhigh_po_2p85_1_14/Rin sky130_asc_res_xhigh_po_2p85_1_14/Rin.t0 4.85
R32887 a_37148_9587.t0 a_37148_9587.t1 7.619
R32888 sky130_asc_res_xhigh_po_2p85_1_2/Rin sky130_asc_res_xhigh_po_2p85_1_3/Rout 35.865
R32889 sky130_asc_res_xhigh_po_2p85_1_3/Rout sky130_asc_res_xhigh_po_2p85_1_2/Rin.t0 4.85
R32890 sky130_asc_res_xhigh_po_2p85_1_1/Rout sky130_asc_res_xhigh_po_2p85_1_0/Rin 239.877
R32891 sky130_asc_res_xhigh_po_2p85_1_0/Rin sky130_asc_res_xhigh_po_2p85_1_0/Rin.t0 4.871
R32892 sky130_asc_res_xhigh_po_2p85_1_29/Rout sky130_asc_res_xhigh_po_2p85_1_28/Rin 20.304
R32893 sky130_asc_res_xhigh_po_2p85_1_28/Rin sky130_asc_res_xhigh_po_2p85_1_29/Rout.t0 4.85
R32894 sky130_asc_res_xhigh_po_2p85_1_26/Rin sky130_asc_res_xhigh_po_2p85_1_27/Rout 21.953
R32895 sky130_asc_res_xhigh_po_2p85_1_27/Rout sky130_asc_res_xhigh_po_2p85_1_26/Rin.t0 4.85
R32896 a_27838_5827.t0 a_27838_5827.t1 7.619
R32897 sky130_asc_res_xhigh_po_2p85_1_24/Rin sky130_asc_res_xhigh_po_2p85_1_25/Rout 66.68
R32898 sky130_asc_res_xhigh_po_2p85_1_25/Rout sky130_asc_res_xhigh_po_2p85_1_24/Rin.t0 4.85
R32899 sky130_asc_res_xhigh_po_2p85_1_9/Rout sky130_asc_res_xhigh_po_2p85_2_0/Rin 62.118
R32900 sky130_asc_res_xhigh_po_2p85_2_0/Rin sky130_asc_res_xhigh_po_2p85_1_9/Rout.t0 4.85
R32901 a_15392_13347.t0 a_15392_13347.t1 7.619
R32902 sky130_asc_res_xhigh_po_2p85_1_3/Rin sky130_asc_res_xhigh_po_2p85_1_4/Rout 11.802
R32903 sky130_asc_res_xhigh_po_2p85_1_4/Rout sky130_asc_res_xhigh_po_2p85_1_4/Rout.t0 4.868
R32904 sky130_asc_res_xhigh_po_2p85_1_15/Rin sky130_asc_res_xhigh_po_2p85_1_16/Rout 36.059
R32905 sky130_asc_res_xhigh_po_2p85_1_16/Rout sky130_asc_res_xhigh_po_2p85_1_16/Rout.t0 4.871
R32906 sky130_asc_res_xhigh_po_2p85_1_13/Rin sky130_asc_res_xhigh_po_2p85_1_14/Rout 34.118
R32907 sky130_asc_res_xhigh_po_2p85_1_14/Rout sky130_asc_res_xhigh_po_2p85_1_14/Rout.t0 4.868
R32908 sky130_asc_res_xhigh_po_2p85_1_12/Rout sky130_asc_res_xhigh_po_2p85_1_11/Rin 24.949
R32909 sky130_asc_res_xhigh_po_2p85_1_11/Rin sky130_asc_res_xhigh_po_2p85_1_12/Rout.t0 4.85
R32910 sky130_asc_res_xhigh_po_2p85_1_18/Rout sky130_asc_res_xhigh_po_2p85_1_17/Rin 48.898
R32911 sky130_asc_res_xhigh_po_2p85_1_17/Rin sky130_asc_res_xhigh_po_2p85_1_18/Rout.t0 4.85
R32912 sky130_asc_res_xhigh_po_2p85_1_22/Rin sky130_asc_res_xhigh_po_2p85_1_23/Rout 39.244
R32913 sky130_asc_res_xhigh_po_2p85_1_23/Rout sky130_asc_res_xhigh_po_2p85_1_22/Rin.t0 4.85
R32914 sky130_asc_res_xhigh_po_2p85_1_10/Rin sky130_asc_res_xhigh_po_2p85_1_11/Rout 45.745
R32915 sky130_asc_res_xhigh_po_2p85_1_11/Rout sky130_asc_res_xhigh_po_2p85_1_10/Rin.t0 4.85
R32916 a_22350_5827.t0 a_22350_5827.t1 7.619
R32917 a_41754_24627.t0 a_41754_24627.t1 7.619
R32918 sky130_asc_res_xhigh_po_2p85_1_30/Rout sky130_asc_res_xhigh_po_2p85_1_29/Rin 16.826
R32919 sky130_asc_res_xhigh_po_2p85_1_29/Rin sky130_asc_res_xhigh_po_2p85_1_30/Rout.t0 4.85
R32920 a_28916_9587.t0 a_28916_9587.t1 7.619
R32921 sky130_asc_res_xhigh_po_2p85_1_7/Rout sky130_asc_res_xhigh_po_2p85_1_6/Rin 62.403
R32922 sky130_asc_res_xhigh_po_2p85_1_6/Rin sky130_asc_res_xhigh_po_2p85_1_7/Rout.t0 4.85
R32923 a_15392_17107.t0 a_15392_17107.t1 7.619
R32924 sky130_asc_res_xhigh_po_2p85_1_23/Rin sky130_asc_res_xhigh_po_2p85_1_24/Rout 71.046
R32925 sky130_asc_res_xhigh_po_2p85_1_24/Rout sky130_asc_res_xhigh_po_2p85_1_24/Rout.t0 4.85
R32926 sky130_asc_res_xhigh_po_2p85_1_4/Rin sky130_asc_res_xhigh_po_2p85_1_5/Rout 25.102
R32927 sky130_asc_res_xhigh_po_2p85_1_5/Rout sky130_asc_res_xhigh_po_2p85_1_5/Rout.t0 4.868
R32928 a_12648_17107.t0 a_12648_17107.t1 7.619
R32929 sky130_asc_res_xhigh_po_2p85_1_13/Rout sky130_asc_res_xhigh_po_2p85_1_12/Rin 52.669
R32930 sky130_asc_res_xhigh_po_2p85_1_12/Rin sky130_asc_res_xhigh_po_2p85_1_12/Rin.t0 4.85
R32931 a_39892_9587.t0 a_39892_9587.t1 7.619
R32932 sky130_asc_res_xhigh_po_2p85_1_2/Rout sky130_asc_res_xhigh_po_2p85_1_1/Rin 45.771
R32933 sky130_asc_res_xhigh_po_2p85_1_1/Rin sky130_asc_res_xhigh_po_2p85_1_2/Rout.t0 4.85
R32934 a_31660_9587.t0 a_31660_9587.t1 7.619
R32935 porst.n0 porst.t4 180.68
R32936 porst.n17 porst.t8 154.653
R32937 porst.n14 porst.t7 154.653
R32938 porst.n3 porst.t0 154.653
R32939 porst.n11 porst.t6 154.653
R32940 porst.n2 porst.t3 154.653
R32941 porst.n8 porst.t5 154.653
R32942 porst.n1 porst.t1 154.653
R32943 porst.n4 porst.t2 154.652
R32944 porst.n9 porst.n8 105.076
R32945 porst.n23 porst.n22 85.333
R32946 porst.n22 porst.n21 85.333
R32947 porst.n21 porst.n20 85.333
R32948 porst.n20 porst.n19 85.333
R32949 porst.n19 porst.n16 85.333
R32950 porst.n16 porst.n13 85.333
R32951 porst.n13 porst.n10 85.333
R32952 porst.n10 porst.n7 85.333
R32953 porst.n7 porst.n5 85.333
R32954 porst.n5 porst.n4 78.892
R32955 porst.n12 porst.n11 78.084
R32956 porst.n23 porst.n0 76
R32957 porst.n22 porst.n1 76
R32958 porst.n21 porst.n2 76
R32959 porst.n20 porst.n3 76
R32960 porst.n19 porst.n18 76
R32961 porst.n16 porst.n15 76
R32962 porst.n13 porst.n12 76
R32963 porst.n10 porst.n9 76
R32964 porst.n7 porst.n6 76
R32965 porst porst.n23 68.266
R32966 porst.n5 porst 52.391
R32967 porst.n15 porst.n14 51.092
R32968 porst.n18 porst.n17 24.1
R32969 sky130_asc_res_xhigh_po_2p85_1_22/Rout sky130_asc_res_xhigh_po_2p85_1_21/Rin 62.827
R32970 sky130_asc_res_xhigh_po_2p85_1_21/Rin sky130_asc_res_xhigh_po_2p85_1_22/Rout.t0 4.85
R32971 sky130_asc_res_xhigh_po_2p85_1_26/Rout sky130_asc_res_xhigh_po_2p85_1_25/Rin 32.359
R32972 sky130_asc_res_xhigh_po_2p85_1_25/Rin sky130_asc_res_xhigh_po_2p85_1_26/Rout.t0 4.85
R32973 sky130_asc_res_xhigh_po_2p85_1_6/Rout sky130_asc_res_xhigh_po_2p85_1_5/Rin 16.835
R32974 sky130_asc_res_xhigh_po_2p85_1_5/Rin sky130_asc_res_xhigh_po_2p85_1_6/Rout.t0 4.85
C0 sky130_asc_res_xhigh_po_2p85_1_9/Rin sky130_asc_res_xhigh_po_2p85_1_12/Rin 0.16fF
C1 VDD a_25584_13347# 0.38fF
C2 sky130_asc_res_xhigh_po_2p85_1_29/Rout sky130_asc_res_xhigh_po_2p85_1_28/Rout 0.23fF
C3 sky130_asc_res_xhigh_po_2p85_1_18/Rout sky130_asc_res_xhigh_po_2p85_1_7/Rin 0.17fF
C4 vbg sky130_asc_pfet_01v8_lvt_60_1/DRAIN 0.25fF
C5 sky130_asc_pfet_01v8_lvt_60_0/GATE sky130_asc_pfet_01v8_lvt_6_1/DRAIN 5.75fF
C6 sky130_asc_res_xhigh_po_2p85_1_0/Rin a_12648_13347# 0.02fF
C7 vbg sky130_asc_res_xhigh_po_2p85_1_0/Rin 0.12fF
C8 sky130_asc_res_xhigh_po_2p85_1_22/Rin sky130_asc_res_xhigh_po_2p85_1_22/Rout 0.44fF
C9 vbg a_41754_20867# 0.02fF
C10 sky130_asc_res_xhigh_po_2p85_1_14/Rin sky130_asc_res_xhigh_po_2p85_1_12/Rin 0.60fF
C11 sky130_asc_res_xhigh_po_2p85_1_9/Rin sky130_asc_res_xhigh_po_2p85_1_24/Rin 0.05fF
C12 VDD sky130_asc_pfet_01v8_lvt_6_1/DRAIN 11.33fF
C13 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_res_xhigh_po_2p85_1_29/Rout 0.02fF
C14 sky130_asc_nfet_01v8_lvt_1_0/DRAIN a_8728_24627# 0.41fF
C15 sky130_asc_res_xhigh_po_2p85_1_24/Rout a_19606_5827# 0.00fF
C16 sky130_asc_pfet_01v8_lvt_60_1/DRAIN sky130_asc_res_xhigh_po_2p85_1_0/Rin 0.28fF
C17 sky130_asc_res_xhigh_po_2p85_1_24/Rout a_25094_5827# 0.02fF
C18 sky130_asc_pfet_01v8_lvt_60_0/GATE sky130_asc_nfet_01v8_lvt_1_0/DRAIN 9.76fF
C19 VDD a_12648_9587# 0.25fF
C20 sky130_asc_res_xhigh_po_2p85_1_0/Rin a_9904_13347# 0.02fF
C21 sky130_asc_res_xhigh_po_2p85_1_30/Rout sky130_asc_res_xhigh_po_2p85_1_12/Rin 0.01fF
C22 sky130_asc_res_xhigh_po_2p85_1_22/Rin sky130_asc_res_xhigh_po_2p85_1_26/Rout 0.04fF
C23 sky130_asc_res_xhigh_po_2p85_1_9/Rin sky130_asc_res_xhigh_po_2p85_1_22/Rout 0.12fF
C24 sky130_asc_res_xhigh_po_2p85_1_10/Rin sky130_asc_res_xhigh_po_2p85_1_12/Rin 1.06fF
C25 sky130_asc_res_xhigh_po_2p85_1_22/Rin sky130_asc_res_xhigh_po_2p85_1_26/Rin 0.08fF
C26 sky130_asc_res_xhigh_po_2p85_1_2/Rin sky130_asc_res_xhigh_po_2p85_1_24/Rin 0.08fF
C27 VDD sky130_asc_res_xhigh_po_2p85_1_24/Rout 0.67fF
C28 VDD a_41754_35907# 0.39fF
C29 VDD sky130_asc_nfet_01v8_lvt_1_0/DRAIN 10.14fF
C30 sky130_asc_pfet_01v8_lvt_60_0/GATE vbg 38.82fF
C31 sky130_asc_res_xhigh_po_2p85_1_22/Rout sky130_asc_res_xhigh_po_2p85_1_24/Rin 0.47fF
C32 sky130_asc_res_xhigh_po_2p85_1_9/Rin sky130_asc_res_xhigh_po_2p85_1_30/Rout 0.02fF
C33 sky130_asc_res_xhigh_po_2p85_1_9/Rin sky130_asc_res_xhigh_po_2p85_1_10/Rin 0.22fF
C34 VDD a_12648_13347# 0.38fF
C35 sky130_asc_res_xhigh_po_2p85_1_24/Rout a_16849_5827# 0.00fF
C36 sky130_asc_res_xhigh_po_2p85_1_5/Rout a_9904_13347# 0.03fF
C37 VDD vbg 22.63fF
C38 sky130_asc_res_xhigh_po_2p85_1_0/Rin sky130_asc_res_xhigh_po_2p85_1_5/Rout 0.29fF
C39 VDD a_9904_9587# 0.38fF
C40 sky130_asc_res_xhigh_po_2p85_1_0/Rin a_9904_5827# 0.01fF
C41 sky130_asc_pfet_01v8_lvt_60_0/GATE sky130_asc_pfet_01v8_lvt_60_1/DRAIN 39.11fF
C42 sky130_asc_res_xhigh_po_2p85_1_22/Rin sky130_asc_res_xhigh_po_2p85_1_28/Rout 0.13fF
C43 sky130_asc_res_xhigh_po_2p85_1_17/Rout sky130_asc_res_xhigh_po_2p85_1_16/Rout 0.23fF
C44 a_12648_13347# sky130_asc_res_xhigh_po_2p85_1_9/Rout 0.29fF
C45 sky130_asc_pfet_01v8_lvt_60_0/GATE sky130_asc_res_xhigh_po_2p85_1_0/Rin 0.04fF
C46 sky130_asc_res_xhigh_po_2p85_1_10/Rin sky130_asc_res_xhigh_po_2p85_1_14/Rin 0.27fF
C47 VDD a_34404_9587# 0.25fF
C48 sky130_asc_res_xhigh_po_2p85_1_4/Rout sky130_asc_res_xhigh_po_2p85_1_2/Rout 0.12fF
C49 sky130_asc_res_xhigh_po_2p85_1_24/Rin sky130_asc_res_xhigh_po_2p85_1_26/Rout 0.45fF
C50 VDD sky130_asc_pfet_01v8_lvt_60_1/DRAIN 24.33fF
C51 sky130_asc_res_xhigh_po_2p85_1_24/Rin sky130_asc_res_xhigh_po_2p85_1_26/Rin 0.09fF
C52 sky130_asc_res_xhigh_po_2p85_1_6/Rout sky130_asc_res_xhigh_po_2p85_1_5/Rout 0.22fF
C53 VDD a_9904_13347# 0.38fF
C54 VDD sky130_asc_res_xhigh_po_2p85_1_0/Rin 4.38fF
C55 VDD a_41754_20867# 0.39fF
C56 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_res_xhigh_po_2p85_1_22/Rin 0.89fF
C57 porst sky130_asc_res_xhigh_po_2p85_1_6/Rout 0.04fF
C58 VDD sky130_asc_res_xhigh_po_2p85_1_16/Rout 0.50fF
C59 sky130_asc_pfet_01v8_lvt_60_0/GATE sky130_asc_res_xhigh_po_2p85_1_6/Rout 0.07fF
C60 porst sky130_asc_res_xhigh_po_2p85_1_5/Rout 0.18fF
C61 sky130_asc_pfet_01v8_lvt_60_0/GATE sky130_asc_res_xhigh_po_2p85_1_5/Rout 0.09fF
C62 VDD a_26159_9587# 0.25fF
C63 sky130_asc_res_xhigh_po_2p85_1_16/Rout sky130_asc_res_xhigh_po_2p85_1_12/Rout 0.21fF
C64 sky130_asc_pfet_01v8_lvt_60_0/GATE a_8728_24627# 0.20fF
C65 sky130_asc_res_xhigh_po_2p85_1_0/Rin sky130_asc_res_xhigh_po_2p85_1_9/Rout 0.00fF
C66 VDD sky130_asc_res_xhigh_po_2p85_1_6/Rout 0.43fF
C67 sky130_asc_pfet_01v8_lvt_60_0/GATE porst 3.26fF
C68 sky130_asc_res_xhigh_po_2p85_1_24/Rin sky130_asc_res_xhigh_po_2p85_1_28/Rout 0.13fF
C69 VDD sky130_asc_res_xhigh_po_2p85_1_5/Rout 0.55fF
C70 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_res_xhigh_po_2p85_1_12/Rin 0.01fF
C71 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_asc_res_xhigh_po_2p85_1_19/Rin 0.56fF
C72 VDD sky130_asc_res_xhigh_po_2p85_1_17/Rout 0.42fF
C73 sky130_asc_res_xhigh_po_2p85_1_12/Rin sky130_asc_res_xhigh_po_2p85_1_14/Rout 0.56fF
C74 VDD a_9904_5827# 0.42fF
C75 VDD a_8728_24627# 0.45fF
C76 sky130_asc_pfet_01v8_lvt_60_1/DRAIN a_42146_28387# 0.02fF
C77 VDD a_19606_5827# 0.42fF
C78 VDD a_25094_5827# 0.30fF
C79 VDD porst 0.50fF
C80 VDD sky130_asc_pfet_01v8_lvt_60_0/GATE 215.62fF
C81 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_res_xhigh_po_2p85_1_9/Rin 0.12fF
C82 VDD a_30582_5827# 0.42fF
C83 sky130_asc_res_xhigh_po_2p85_1_9/Rin sky130_asc_res_xhigh_po_2p85_1_14/Rout 0.04fF
C84 vbg sky130_asc_res_xhigh_po_2p85_1_18/Rout 0.37fF
C85 a_12648_9587# sky130_asc_res_xhigh_po_2p85_1_21/Rout 0.29fF
C86 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_res_xhigh_po_2p85_1_24/Rin 0.76fF
C87 sky130_asc_res_xhigh_po_2p85_1_22/Rin a_25584_13347# 0.02fF
C88 sky130_asc_res_xhigh_po_2p85_1_26/Rout sky130_asc_res_xhigh_po_2p85_1_26/Rin 0.83fF
C89 sky130_asc_res_xhigh_po_2p85_1_2/Rout sky130_asc_res_xhigh_po_2p85_1_24/Rin 0.00fF
C90 sky130_asc_res_xhigh_po_2p85_1_24/Rout sky130_asc_res_xhigh_po_2p85_1_21/Rout 0.08fF
C91 sky130_asc_res_xhigh_po_2p85_1_14/Rin sky130_asc_res_xhigh_po_2p85_1_14/Rout 0.23fF
C92 VDD sky130_asc_res_xhigh_po_2p85_1_12/Rout 1.07fF
C93 sky130_asc_res_xhigh_po_2p85_1_16/Rout a_37148_5827# 0.28fF
C94 VDD a_16849_5827# 0.42fF
C95 sky130_asc_pfet_01v8_lvt_60_1/DRAIN sky130_asc_res_xhigh_po_2p85_1_18/Rout 0.23fF
C96 VDD sky130_asc_res_xhigh_po_2p85_1_9/Rout 0.92fF
C97 VDD a_33326_5827# 0.42fF
C98 sky130_asc_res_xhigh_po_2p85_1_18/Rout sky130_asc_res_xhigh_po_2p85_1_0/Rin 0.34fF
C99 sky130_asc_res_xhigh_po_2p85_1_7/Rin sky130_asc_res_xhigh_po_2p85_1_7/Rout 1.09fF
C100 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_res_xhigh_po_2p85_1_22/Rout 0.68fF
C101 sky130_asc_res_xhigh_po_2p85_1_28/Rout sky130_asc_res_xhigh_po_2p85_1_26/Rout 0.17fF
C102 sky130_asc_res_xhigh_po_2p85_1_2/Rin sky130_asc_res_xhigh_po_2p85_1_2/Rout 0.56fF
C103 sky130_asc_res_xhigh_po_2p85_1_28/Rout sky130_asc_res_xhigh_po_2p85_1_26/Rin 1.66fF
C104 sky130_asc_res_xhigh_po_2p85_1_12/Rout a_33326_5827# 0.06fF
C105 a_26159_9587# sky130_asc_res_xhigh_po_2p85_1_29/Rout 0.28fF
C106 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_res_xhigh_po_2p85_1_30/Rout 0.79fF
C107 sky130_asc_res_xhigh_po_2p85_1_4/Rout a_9904_9587# 0.02fF
C108 sky130_asc_res_xhigh_po_2p85_1_10/Rin sky130_asc_res_xhigh_po_2p85_1_14/Rout 0.25fF
C109 VDD a_42146_28387# 0.49fF
C110 sky130_asc_res_xhigh_po_2p85_1_16/Rout a_39892_5827# 0.02fF
C111 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_asc_res_xhigh_po_2p85_1_7/Rin 3.54fF
C112 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_res_xhigh_po_2p85_1_7/Rout 1.32fF
C113 sky130_asc_res_xhigh_po_2p85_1_22/Rin sky130_asc_res_xhigh_po_2p85_1_24/Rout 0.56fF
C114 sky130_asc_res_xhigh_po_2p85_1_18/Rout sky130_asc_res_xhigh_po_2p85_1_17/Rout 0.24fF
C115 VDD a_37148_5827# 0.30fF
C116 sky130_asc_res_xhigh_po_2p85_1_29/Rout a_30582_5827# 0.02fF
C117 a_9904_13347# sky130_asc_res_xhigh_po_2p85_1_4/Rout 0.01fF
C118 sky130_asc_res_xhigh_po_2p85_1_0/Rin sky130_asc_res_xhigh_po_2p85_1_4/Rout 0.93fF
C119 sky130_asc_res_xhigh_po_2p85_1_12/Rout a_37148_5827# 0.43fF
C120 a_25584_13347# sky130_asc_res_xhigh_po_2p85_1_22/Rout 0.01fF
C121 VDD sky130_asc_res_xhigh_po_2p85_1_29/Rout 0.47fF
C122 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_asc_pfet_01v8_lvt_60_2/DRAIN 0.15fF
C123 sky130_asc_res_xhigh_po_2p85_1_19/Rin sky130_asc_pfet_01v8_lvt_6_1/DRAIN 0.19fF
C124 VDD sky130_asc_res_xhigh_po_2p85_1_18/Rout 0.69fF
C125 sky130_asc_res_xhigh_po_2p85_1_24/Rin a_12648_9587# 0.41fF
C126 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_res_xhigh_po_2p85_1_7/Rin 0.22fF
C127 sky130_asc_res_xhigh_po_2p85_1_9/Rin sky130_asc_res_xhigh_po_2p85_1_24/Rout 1.30fF
C128 sky130_asc_res_xhigh_po_2p85_1_5/Rout sky130_asc_res_xhigh_po_2p85_1_4/Rout 0.23fF
C129 VDD a_39892_5827# 0.42fF
C130 a_12648_13347# sky130_asc_res_xhigh_po_2p85_1_9/Rin 0.28fF
C131 sky130_asc_res_xhigh_po_2p85_1_0/Rin sky130_asc_res_xhigh_po_2p85_1_22/Rin 0.02fF
C132 sky130_asc_res_xhigh_po_2p85_1_24/Rin sky130_asc_res_xhigh_po_2p85_1_24/Rout 0.29fF
C133 a_34404_9587# sky130_asc_res_xhigh_po_2p85_1_12/Rin 0.55fF
C134 VDD sky130_asc_res_xhigh_po_2p85_1_21/Rout 0.52fF
C135 sky130_asc_res_xhigh_po_2p85_1_19/Rin a_41754_35907# 0.02fF
C136 sky130_asc_nfet_01v8_lvt_1_1/DRAIN sky130_asc_res_xhigh_po_2p85_1_19/Rout 0.04fF
C137 sky130_asc_res_xhigh_po_2p85_1_22/Rout a_12648_9587# 0.30fF
C138 sky130_asc_res_xhigh_po_2p85_1_9/Rin a_34404_9587# 0.01fF
C139 a_9904_9587# sky130_asc_res_xhigh_po_2p85_1_24/Rin 0.28fF
C140 sky130_asc_nfet_01v8_lvt_1_1/DRAIN sky130_asc_res_xhigh_po_2p85_1_7/Rin 0.06fF
C141 sky130_asc_res_xhigh_po_2p85_1_2/Rin sky130_asc_res_xhigh_po_2p85_1_24/Rout 0.08fF
C142 VDD sky130_asc_res_xhigh_po_2p85_1_4/Rout 0.42fF
C143 a_42146_28387# sky130_asc_res_xhigh_po_2p85_1_18/Rout 0.01fF
C144 sky130_asc_res_xhigh_po_2p85_1_22/Rout sky130_asc_res_xhigh_po_2p85_1_24/Rout 0.00fF
C145 sky130_asc_res_xhigh_po_2p85_1_16/Rout sky130_asc_res_xhigh_po_2p85_1_12/Rin 0.22fF
C146 vbg sky130_asc_res_xhigh_po_2p85_1_19/Rin 0.41fF
C147 sky130_asc_res_xhigh_po_2p85_1_2/Rin a_12648_13347# 0.02fF
C148 sky130_asc_res_xhigh_po_2p85_1_0/Rin sky130_asc_res_xhigh_po_2p85_1_9/Rin 0.02fF
C149 sky130_asc_res_xhigh_po_2p85_1_22/Rin a_25094_5827# 0.02fF
C150 a_34404_9587# sky130_asc_res_xhigh_po_2p85_1_14/Rin 0.28fF
C151 sky130_asc_res_xhigh_po_2p85_1_2/Rin a_9904_9587# 0.43fF
C152 a_41264_13347# sky130_asc_res_xhigh_po_2p85_1_16/Rout 0.01fF
C153 sky130_asc_res_xhigh_po_2p85_1_9/Rin a_26159_9587# 0.02fF
C154 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_asc_pfet_01v8_lvt_6_1/DRAIN 0.03fF
C155 sky130_asc_nfet_01v8_lvt_1_1/DRAIN sky130_asc_pfet_01v8_lvt_60_2/DRAIN 2.29fF
C156 sky130_asc_res_xhigh_po_2p85_1_19/Rin sky130_asc_pfet_01v8_lvt_60_1/DRAIN 2.17fF
C157 VDD sky130_asc_res_xhigh_po_2p85_1_22/Rin 0.60fF
C158 sky130_asc_pfet_01v8_lvt_6_1/DRAIN sky130_asc_res_xhigh_po_2p85_1_7/Rin 0.02fF
C159 sky130_asc_nfet_01v8_lvt_1_0/DRAIN sky130_asc_res_xhigh_po_2p85_1_7/Rout 0.02fF
C160 sky130_asc_res_xhigh_po_2p85_1_24/Rout sky130_asc_res_xhigh_po_2p85_1_26/Rout 0.37fF
C161 sky130_asc_res_xhigh_po_2p85_1_16/Rout sky130_asc_res_xhigh_po_2p85_1_14/Rin 1.72fF
C162 sky130_asc_res_xhigh_po_2p85_1_24/Rout sky130_asc_res_xhigh_po_2p85_1_26/Rin 0.12fF
C163 sky130_asc_res_xhigh_po_2p85_1_12/Rin a_30582_5827# 0.49fF
C164 a_9904_13347# sky130_asc_res_xhigh_po_2p85_1_2/Rin 0.81fF
C165 sky130_asc_res_xhigh_po_2p85_1_0/Rin sky130_asc_res_xhigh_po_2p85_1_2/Rin 0.17fF
C166 sky130_asc_res_xhigh_po_2p85_1_17/Rout a_41264_13347# 0.02fF
C167 sky130_asc_res_xhigh_po_2p85_1_10/Rin a_34404_9587# 0.36fF
C168 sky130_asc_res_xhigh_po_2p85_1_0/Rin sky130_asc_res_xhigh_po_2p85_1_22/Rout 0.00fF
C169 sky130_asc_res_xhigh_po_2p85_1_22/Rin sky130_asc_res_xhigh_po_2p85_1_9/Rout 0.20fF
C170 VDD sky130_asc_res_xhigh_po_2p85_1_12/Rin 4.31fF
C171 sky130_asc_res_xhigh_po_2p85_1_24/Rin a_19606_5827# 0.48fF
C172 sky130_asc_res_xhigh_po_2p85_1_19/Rout a_41754_35907# 0.01fF
C173 sky130_asc_nfet_01v8_lvt_1_0/DRAIN sky130_asc_res_xhigh_po_2p85_1_19/Rout 0.00fF
C174 sky130_asc_res_xhigh_po_2p85_1_12/Rin sky130_asc_res_xhigh_po_2p85_1_12/Rout 0.23fF
C175 sky130_asc_pfet_01v8_lvt_6_1/DRAIN sky130_asc_pfet_01v8_lvt_60_2/DRAIN 2.05fF
C176 VDD sky130_asc_res_xhigh_po_2p85_1_9/Rin 0.74fF
C177 sky130_asc_nfet_01v8_lvt_1_0/DRAIN sky130_asc_res_xhigh_po_2p85_1_7/Rin 0.03fF
C178 sky130_asc_res_xhigh_po_2p85_1_24/Rout sky130_asc_res_xhigh_po_2p85_1_28/Rout 0.03fF
C179 VDD a_41264_13347# 0.38fF
C180 a_26159_9587# sky130_asc_res_xhigh_po_2p85_1_30/Rout 0.28fF
C181 sky130_asc_pfet_01v8_lvt_60_0/GATE sky130_asc_res_xhigh_po_2p85_1_19/Rin 0.52fF
C182 vbg sky130_asc_res_xhigh_po_2p85_1_19/Rout 0.98fF
C183 VDD sky130_asc_res_xhigh_po_2p85_1_24/Rin 6.29fF
C184 sky130_asc_res_xhigh_po_2p85_1_12/Rin a_33326_5827# 0.01fF
C185 vbg sky130_asc_res_xhigh_po_2p85_1_7/Rin 0.25fF
C186 sky130_asc_res_xhigh_po_2p85_1_9/Rin sky130_asc_res_xhigh_po_2p85_1_9/Rout 0.38fF
C187 VDD sky130_asc_res_xhigh_po_2p85_1_14/Rin 0.33fF
C188 VDD sky130_asc_res_xhigh_po_2p85_1_19/Rin 0.79fF
C189 sky130_asc_res_xhigh_po_2p85_1_9/Rout sky130_asc_res_xhigh_po_2p85_1_24/Rin 0.52fF
C190 sky130_asc_res_xhigh_po_2p85_1_14/Rin sky130_asc_res_xhigh_po_2p85_1_12/Rout 0.30fF
C191 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_res_xhigh_po_2p85_1_24/Rout 0.07fF
C192 sky130_asc_nfet_01v8_lvt_1_0/DRAIN sky130_asc_pfet_01v8_lvt_60_2/DRAIN 0.42fF
C193 sky130_asc_nfet_01v8_lvt_1_1/DRAIN sky130_asc_pfet_01v8_lvt_6_1/DRAIN 2.87fF
C194 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_asc_pfet_01v8_lvt_60_1/DRAIN 0.14fF
C195 VDD sky130_asc_res_xhigh_po_2p85_1_2/Rin 0.49fF
C196 sky130_asc_res_xhigh_po_2p85_1_7/Rout sky130_asc_res_xhigh_po_2p85_1_6/Rout 0.25fF
C197 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_asc_res_xhigh_po_2p85_1_0/Rin 4.48fF
C198 sky130_asc_pfet_01v8_lvt_60_1/DRAIN sky130_asc_res_xhigh_po_2p85_1_7/Rin 0.05fF
C199 VDD sky130_asc_res_xhigh_po_2p85_1_22/Rout 1.35fF
C200 a_8728_24627# sky130_asc_res_xhigh_po_2p85_1_7/Rout 0.04fF
C201 sky130_asc_res_xhigh_po_2p85_1_7/Rin sky130_asc_res_xhigh_po_2p85_1_0/Rin 0.03fF
C202 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_asc_res_xhigh_po_2p85_1_16/Rout 0.19fF
C203 sky130_asc_res_xhigh_po_2p85_1_7/Rin a_41754_20867# 0.01fF
C204 a_19606_5827# sky130_asc_res_xhigh_po_2p85_1_26/Rout 0.28fF
C205 VDD sky130_asc_res_xhigh_po_2p85_1_30/Rout 0.25fF
C206 a_12648_13347# sky130_asc_res_xhigh_po_2p85_1_2/Rout 0.01fF
C207 sky130_asc_pfet_01v8_lvt_60_0/GATE sky130_asc_res_xhigh_po_2p85_1_7/Rout 0.15fF
C208 VDD sky130_asc_res_xhigh_po_2p85_1_10/Rin 1.17fF
C209 a_19606_5827# sky130_asc_res_xhigh_po_2p85_1_26/Rin 0.34fF
C210 sky130_asc_res_xhigh_po_2p85_1_26/Rout a_25094_5827# 0.94fF
C211 a_25094_5827# sky130_asc_res_xhigh_po_2p85_1_26/Rin 0.54fF
C212 sky130_asc_res_xhigh_po_2p85_1_9/Rout sky130_asc_res_xhigh_po_2p85_1_22/Rout 0.90fF
C213 sky130_asc_res_xhigh_po_2p85_1_2/Rout a_9904_9587# 0.01fF
C214 a_34404_9587# sky130_asc_res_xhigh_po_2p85_1_14/Rout 0.31fF
C215 sky130_asc_res_xhigh_po_2p85_1_10/Rin sky130_asc_res_xhigh_po_2p85_1_12/Rout 0.45fF
C216 sky130_asc_nfet_01v8_lvt_1_0/DRAIN sky130_asc_nfet_01v8_lvt_1_1/DRAIN 1.11fF
C217 VDD sky130_asc_res_xhigh_po_2p85_1_7/Rout 0.60fF
C218 sky130_asc_pfet_01v8_lvt_60_1/DRAIN sky130_asc_pfet_01v8_lvt_60_2/DRAIN 0.34fF
C219 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_asc_res_xhigh_po_2p85_1_17/Rout 0.08fF
C220 VDD sky130_asc_res_xhigh_po_2p85_1_26/Rout 2.43fF
C221 VDD sky130_asc_res_xhigh_po_2p85_1_26/Rin 0.63fF
C222 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_res_xhigh_po_2p85_1_0/Rin 0.22fF
C223 sky130_asc_res_xhigh_po_2p85_1_9/Rin sky130_asc_res_xhigh_po_2p85_1_29/Rout 0.04fF
C224 sky130_asc_res_xhigh_po_2p85_1_10/Rin a_33326_5827# 0.06fF
C225 sky130_asc_res_xhigh_po_2p85_1_7/Rin a_8728_24627# 0.04fF
C226 sky130_asc_pfet_01v8_lvt_60_0/GATE sky130_asc_res_xhigh_po_2p85_1_19/Rout 1.16fF
C227 sky130_asc_res_xhigh_po_2p85_1_14/Rin a_37148_5827# 0.47fF
C228 sky130_asc_res_xhigh_po_2p85_1_28/Rout a_19606_5827# 0.19fF
C229 a_9904_13347# sky130_asc_res_xhigh_po_2p85_1_2/Rout 0.32fF
C230 sky130_asc_pfet_01v8_lvt_60_0/GATE sky130_asc_res_xhigh_po_2p85_1_7/Rin 0.19fF
C231 sky130_asc_res_xhigh_po_2p85_1_0/Rin sky130_asc_res_xhigh_po_2p85_1_2/Rout 3.59fF
C232 a_16849_5827# sky130_asc_res_xhigh_po_2p85_1_26/Rin 0.28fF
C233 sky130_asc_res_xhigh_po_2p85_1_28/Rout a_25094_5827# 0.17fF
C234 sky130_asc_pfet_01v8_lvt_60_2/DRAIN a_26159_9587# 0.48fF
C235 sky130_asc_res_xhigh_po_2p85_1_28/Rout a_30582_5827# 0.01fF
C236 VDD sky130_asc_res_xhigh_po_2p85_1_19/Rout 6.54fF
C237 VDD sky130_asc_res_xhigh_po_2p85_1_7/Rin 2.16fF
C238 sky130_asc_nfet_01v8_lvt_1_1/DRAIN sky130_asc_pfet_01v8_lvt_60_1/DRAIN 2.32fF
C239 VDD sky130_asc_res_xhigh_po_2p85_1_28/Rout 0.62fF
C240 sky130_asc_res_xhigh_po_2p85_1_19/Rin sky130_asc_res_xhigh_po_2p85_1_18/Rout 0.01fF
C241 sky130_asc_nfet_01v8_lvt_1_1/DRAIN sky130_asc_res_xhigh_po_2p85_1_0/Rin 0.03fF
C242 sky130_asc_res_xhigh_po_2p85_1_9/Rin sky130_asc_res_xhigh_po_2p85_1_21/Rout 0.09fF
C243 sky130_asc_res_xhigh_po_2p85_1_10/Rin a_37148_5827# 0.01fF
C244 sky130_asc_pfet_01v8_lvt_60_0/GATE sky130_asc_pfet_01v8_lvt_60_2/DRAIN 44.86fF
C245 a_16849_5827# sky130_asc_res_xhigh_po_2p85_1_28/Rout 0.45fF
C246 sky130_asc_res_xhigh_po_2p85_1_14/Rin a_39892_5827# 0.01fF
C247 a_12648_9587# sky130_asc_res_xhigh_po_2p85_1_24/Rout 0.08fF
C248 sky130_asc_res_xhigh_po_2p85_1_2/Rout a_9904_5827# 0.02fF
C249 sky130_asc_res_xhigh_po_2p85_1_24/Rin sky130_asc_res_xhigh_po_2p85_1_21/Rout 0.00fF
C250 sky130_asc_res_xhigh_po_2p85_1_0/Rin a_25584_13347# 0.02fF
C251 sky130_asc_res_xhigh_po_2p85_1_14/Rout a_30582_5827# 0.28fF
C252 sky130_asc_res_xhigh_po_2p85_1_30/Rout sky130_asc_res_xhigh_po_2p85_1_29/Rout 0.28fF
C253 VDD sky130_asc_pfet_01v8_lvt_60_2/DRAIN 44.20fF
C254 VDD sky130_asc_res_xhigh_po_2p85_1_14/Rout 0.61fF
C255 sky130_asc_pfet_01v8_lvt_60_1/DRAIN sky130_asc_pfet_01v8_lvt_6_1/DRAIN 4.55fF
C256 VDD sky130_asc_res_xhigh_po_2p85_1_2/Rout 0.57fF
C257 sky130_asc_pfet_01v8_lvt_6_1/DRAIN sky130_asc_res_xhigh_po_2p85_1_0/Rin 0.22fF
C258 sky130_asc_pfet_01v8_lvt_60_0/GATE sky130_asc_nfet_01v8_lvt_1_1/DRAIN 3.13fF
C259 sky130_asc_res_xhigh_po_2p85_1_22/Rout sky130_asc_res_xhigh_po_2p85_1_21/Rout 0.23fF
C260 sky130_asc_pfet_01v8_lvt_60_2/DRAIN sky130_asc_res_xhigh_po_2p85_1_9/Rout 1.43fF
C261 a_9904_9587# sky130_asc_res_xhigh_po_2p85_1_24/Rout 0.28fF
C262 sky130_asc_res_xhigh_po_2p85_1_2/Rin sky130_asc_res_xhigh_po_2p85_1_4/Rout 0.24fF
C263 sky130_asc_res_xhigh_po_2p85_1_9/Rin sky130_asc_res_xhigh_po_2p85_1_22/Rin 0.03fF
C264 sky130_asc_res_xhigh_po_2p85_1_14/Rout a_33326_5827# 0.04fF
C265 VDD sky130_asc_nfet_01v8_lvt_1_1/DRAIN 4.10fF
C266 sky130_asc_res_xhigh_po_2p85_1_19/Rout sky130_asc_res_xhigh_po_2p85_1_18/Rout 0.17fF
C267 a_39892_5827# VSS 2.80fF
C268 a_37148_5827# VSS 2.39fF
C269 a_33326_5827# VSS 2.77fF
C270 a_30582_5827# VSS 2.42fF
C271 sky130_asc_res_xhigh_po_2p85_1_26/Rin VSS 5.55fF
C272 a_25094_5827# VSS 2.41fF
C273 sky130_asc_res_xhigh_po_2p85_1_26/Rout VSS 5.62fF
C274 a_19606_5827# VSS 2.41fF
C275 sky130_asc_res_xhigh_po_2p85_1_28/Rout VSS 4.31fF
C276 a_16849_5827# VSS 2.44fF
C277 a_9904_5827# VSS 2.95fF
C278 sky130_asc_res_xhigh_po_2p85_1_12/Rout VSS 5.09fF
C279 sky130_asc_res_xhigh_po_2p85_1_14/Rout VSS 8.32fF $ **FLOATING
C280 sky130_asc_res_xhigh_po_2p85_1_29/Rout VSS 5.60fF
C281 sky130_asc_res_xhigh_po_2p85_1_21/Rout VSS 5.31fF
C282 sky130_asc_res_xhigh_po_2p85_1_24/Rout VSS 10.20fF $ **FLOATING
C283 sky130_asc_res_xhigh_po_2p85_1_12/Rin VSS 8.07fF $ **FLOATING
C284 sky130_asc_res_xhigh_po_2p85_1_14/Rin VSS 6.34fF $ **FLOATING
C285 a_34404_9587# VSS 2.40fF
C286 sky130_asc_res_xhigh_po_2p85_1_10/Rin VSS 6.39fF
C287 sky130_asc_res_xhigh_po_2p85_1_30/Rout VSS 3.95fF
C288 a_26159_9587# VSS 2.43fF
C289 a_12648_9587# VSS 2.56fF
C290 sky130_asc_res_xhigh_po_2p85_1_24/Rin VSS 9.38fF
C291 a_9904_9587# VSS 2.57fF
C292 sky130_asc_res_xhigh_po_2p85_1_16/Rout VSS 6.25fF $ **FLOATING
C293 a_41264_13347# VSS 2.80fF
C294 sky130_asc_res_xhigh_po_2p85_1_22/Rout VSS 10.11fF
C295 sky130_asc_res_xhigh_po_2p85_1_9/Rout VSS 9.21fF
C296 sky130_asc_res_xhigh_po_2p85_1_2/Rout VSS 8.40fF
C297 sky130_asc_res_xhigh_po_2p85_1_4/Rout VSS 4.03fF $ **FLOATING
C298 a_25584_13347# VSS 2.80fF
C299 sky130_asc_res_xhigh_po_2p85_1_22/Rin VSS 7.25fF
C300 sky130_asc_res_xhigh_po_2p85_1_9/Rin VSS 12.34fF
C301 a_12648_13347# VSS 2.42fF
C302 sky130_asc_res_xhigh_po_2p85_1_2/Rin VSS 7.01fF
C303 a_9904_13347# VSS 2.42fF
C304 sky130_asc_res_xhigh_po_2p85_1_17/Rout VSS 4.73fF
C305 sky130_asc_res_xhigh_po_2p85_1_5/Rout VSS 6.07fF $ **FLOATING
C306 sky130_asc_res_xhigh_po_2p85_1_6/Rout VSS 4.29fF
C307 porst VSS 13.37fF
C308 a_41754_20867# VSS 2.80fF
C309 sky130_asc_res_xhigh_po_2p85_1_0/Rin VSS 31.35fF $ **FLOATING
C310 sky130_asc_res_xhigh_po_2p85_1_7/Rout VSS 9.80fF
C311 a_8728_24627# VSS 2.32fF
C312 sky130_asc_res_xhigh_po_2p85_1_7/Rin VSS 14.46fF
C313 sky130_asc_res_xhigh_po_2p85_1_18/Rout VSS 8.50fF
C314 a_42146_28387# VSS 2.80fF
C315 sky130_asc_pfet_01v8_lvt_60_2/DRAIN VSS 135.58fF
C316 sky130_asc_pfet_01v8_lvt_6_1/DRAIN VSS 12.48fF $ **FLOATING
C317 sky130_asc_pfet_01v8_lvt_60_1/DRAIN VSS 14.82fF $ **FLOATING
C318 a_41754_35907# VSS 2.80fF
C319 sky130_asc_res_xhigh_po_2p85_1_19/Rin VSS 7.37fF
C320 sky130_asc_res_xhigh_po_2p85_1_19/Rout VSS 130.83fF
C321 sky130_asc_nfet_01v8_lvt_1_1/DRAIN VSS 7.22fF $ **FLOATING
C322 sky130_asc_nfet_01v8_lvt_1_0/DRAIN VSS 20.11fF $ **FLOATING
C323 vbg VSS 11.99fF
C324 sky130_asc_pfet_01v8_lvt_60_0/GATE VSS 148.50fF $ **FLOATING
C325 VDD VSS 988.47fF
C326 sky130_asc_res_xhigh_po_2p85_1_5/Rin VSS 1.33fF $ **FLOATING
C327 sky130_asc_res_xhigh_po_2p85_1_6/Rout.t0 VSS 0.12fF
C328 sky130_asc_res_xhigh_po_2p85_1_25/Rin VSS 2.51fF $ **FLOATING
C329 sky130_asc_res_xhigh_po_2p85_1_26/Rout.t0 VSS 0.20fF
C330 sky130_asc_res_xhigh_po_2p85_1_21/Rin VSS 3.12fF $ **FLOATING
C331 sky130_asc_res_xhigh_po_2p85_1_22/Rout.t0 VSS 0.23fF
C332 porst.t4 VSS 1.27fF
C333 porst.n0 VSS 0.20fF $ **FLOATING
C334 porst.t1 VSS 1.25fF
C335 porst.n1 VSS 0.35fF $ **FLOATING
C336 porst.t3 VSS 1.25fF
C337 porst.n2 VSS 0.36fF $ **FLOATING
C338 porst.t0 VSS 1.25fF
C339 porst.n3 VSS 0.35fF $ **FLOATING
C340 porst.t2 VSS 1.25fF
C341 porst.n4 VSS 0.33fF $ **FLOATING
C342 porst.n5 VSS 0.26fF $ **FLOATING
C343 porst.n6 VSS 0.07fF $ **FLOATING
C344 porst.n7 VSS 0.10fF $ **FLOATING
C345 porst.t5 VSS 1.25fF
C346 porst.n8 VSS 0.28fF $ **FLOATING
C347 porst.n9 VSS 0.07fF $ **FLOATING
C348 porst.n10 VSS 0.10fF $ **FLOATING
C349 porst.t6 VSS 1.25fF
C350 porst.n11 VSS 0.28fF $ **FLOATING
C351 porst.n12 VSS 0.07fF $ **FLOATING
C352 porst.n13 VSS 0.10fF $ **FLOATING
C353 porst.t7 VSS 1.25fF
C354 porst.n14 VSS 0.28fF $ **FLOATING
C355 porst.n15 VSS 0.07fF $ **FLOATING
C356 porst.n16 VSS 0.10fF $ **FLOATING
C357 porst.t8 VSS 1.25fF
C358 porst.n17 VSS 0.28fF $ **FLOATING
C359 porst.n18 VSS 0.07fF $ **FLOATING
C360 porst.n19 VSS 0.10fF $ **FLOATING
C361 porst.n20 VSS 0.10fF $ **FLOATING
C362 porst.n21 VSS 0.10fF $ **FLOATING
C363 porst.n22 VSS 0.10fF $ **FLOATING
C364 porst.n23 VSS 0.09fF $ **FLOATING
C365 a_31660_9587.t1 VSS 0.84fF
C366 a_31660_9587.t0 VSS 1.57fF
C367 sky130_asc_res_xhigh_po_2p85_1_1/Rin VSS 3.72fF $ **FLOATING
C368 sky130_asc_res_xhigh_po_2p85_1_2/Rout.t0 VSS 0.29fF
C369 a_39892_9587.t1 VSS 0.97fF
C370 a_39892_9587.t0 VSS 1.83fF
C371 sky130_asc_res_xhigh_po_2p85_1_13/Rout VSS 4.23fF
C372 sky130_asc_res_xhigh_po_2p85_1_12/Rin.t0 VSS 0.29fF
C373 a_12648_17107.t1 VSS 0.84fF
C374 a_12648_17107.t0 VSS 1.57fF
C375 sky130_asc_res_xhigh_po_2p85_1_4/Rin VSS 2.07fF
C376 sky130_asc_res_xhigh_po_2p85_1_5/Rout.t0 VSS 0.17fF
C377 sky130_asc_res_xhigh_po_2p85_1_23/Rin VSS 3.50fF
C378 sky130_asc_res_xhigh_po_2p85_1_24/Rout.t0 VSS 0.23fF
C379 a_15392_17107.t1 VSS 1.10fF
C380 a_15392_17107.t0 VSS 2.05fF
C381 sky130_asc_res_xhigh_po_2p85_1_6/Rin VSS 3.07fF $ **FLOATING
C382 sky130_asc_res_xhigh_po_2p85_1_7/Rout.t0 VSS 0.22fF
C383 a_28916_9587.t1 VSS 0.83fF
C384 a_28916_9587.t0 VSS 1.56fF
C385 sky130_asc_res_xhigh_po_2p85_1_29/Rin VSS 1.22fF $ **FLOATING
C386 sky130_asc_res_xhigh_po_2p85_1_30/Rout.t0 VSS 0.11fF
C387 a_41754_24627.t1 VSS 0.98fF
C388 a_41754_24627.t0 VSS 1.83fF
C389 a_22350_5827.t1 VSS 0.84fF
C390 a_22350_5827.t0 VSS 1.56fF
C391 sky130_asc_res_xhigh_po_2p85_1_11/Rout VSS 1.98fF $ **FLOATING
C392 sky130_asc_res_xhigh_po_2p85_1_10/Rin.t0 VSS 0.15fF
C393 sky130_asc_res_xhigh_po_2p85_1_23/Rout VSS 2.23fF $ **FLOATING
C394 sky130_asc_res_xhigh_po_2p85_1_22/Rin.t0 VSS 0.18fF
C395 sky130_asc_res_xhigh_po_2p85_1_17/Rin VSS 2.66fF $ **FLOATING
C396 sky130_asc_res_xhigh_po_2p85_1_18/Rout.t0 VSS 0.20fF
C397 sky130_asc_res_xhigh_po_2p85_1_11/Rin VSS 1.57fF $ **FLOATING
C398 sky130_asc_res_xhigh_po_2p85_1_12/Rout.t0 VSS 0.13fF
C399 sky130_asc_res_xhigh_po_2p85_1_13/Rin VSS 2.87fF
C400 sky130_asc_res_xhigh_po_2p85_1_14/Rout.t0 VSS 0.22fF
C401 sky130_asc_res_xhigh_po_2p85_1_15/Rin VSS 2.13fF
C402 sky130_asc_res_xhigh_po_2p85_1_16/Rout.t0 VSS 0.17fF
C403 sky130_asc_res_xhigh_po_2p85_1_3/Rin VSS 1.39fF
C404 sky130_asc_res_xhigh_po_2p85_1_4/Rout.t0 VSS 0.12fF
C405 a_15392_13347.t1 VSS 1.10fF
C406 a_15392_13347.t0 VSS 2.05fF
C407 sky130_asc_res_xhigh_po_2p85_2_0/Rin VSS 2.88fF $ **FLOATING
C408 sky130_asc_res_xhigh_po_2p85_1_9/Rout.t0 VSS 0.21fF
C409 sky130_asc_res_xhigh_po_2p85_1_25/Rout VSS 4.88fF $ **FLOATING
C410 sky130_asc_res_xhigh_po_2p85_1_24/Rin.t0 VSS 0.35fF
C411 a_27838_5827.t1 VSS 0.84fF
C412 a_27838_5827.t0 VSS 1.58fF
C413 sky130_asc_res_xhigh_po_2p85_1_27/Rout VSS 1.64fF $ **FLOATING
C414 sky130_asc_res_xhigh_po_2p85_1_26/Rin.t0 VSS 0.12fF
C415 sky130_asc_res_xhigh_po_2p85_1_28/Rin VSS 1.71fF $ **FLOATING
C416 sky130_asc_res_xhigh_po_2p85_1_29/Rout.t0 VSS 0.15fF
C417 sky130_asc_res_xhigh_po_2p85_1_1/Rout VSS 14.86fF
C418 sky130_asc_res_xhigh_po_2p85_1_0/Rin.t0 VSS 0.65fF
C419 sky130_asc_res_xhigh_po_2p85_1_3/Rout VSS 2.17fF $ **FLOATING
C420 sky130_asc_res_xhigh_po_2p85_1_2/Rin.t0 VSS 0.17fF
C421 a_37148_9587.t1 VSS 0.84fF
C422 a_37148_9587.t0 VSS 1.56fF
C423 sky130_asc_res_xhigh_po_2p85_1_15/Rout VSS 2.16fF
C424 sky130_asc_res_xhigh_po_2p85_1_14/Rin.t0 VSS 0.16fF
C425 a_41264_17107.t1 VSS 0.97fF
C426 a_41264_17107.t0 VSS 1.83fF
C427 sky130_asc_res_xhigh_po_2p85_1_16/Rin VSS 1.44fF $ **FLOATING
C428 sky130_asc_res_xhigh_po_2p85_1_17/Rout.t0 VSS 0.13fF
C429 a_39402_28387.t1 VSS 0.84fF
C430 a_39402_28387.t0 VSS 1.56fF
C431 sky130_asc_res_xhigh_po_2p85_1_20/Rout VSS 2.96fF $ **FLOATING
C432 sky130_asc_res_xhigh_po_2p85_1_19/Rin.t0 VSS 0.23fF
C433 a_15392_9587.t1 VSS 1.15fF
C434 a_15392_9587.t0 VSS 2.15fF
C435 sky130_asc_res_xhigh_po_2p85_2_1/Rin VSS 1.63fF $ **FLOATING
C436 sky130_asc_res_xhigh_po_2p85_1_21/Rout.t0 VSS 0.14fF
C437 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n0 VSS 0.02fF $ **FLOATING
C438 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n1 VSS 0.02fF $ **FLOATING
C439 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n2 VSS 0.02fF $ **FLOATING
C440 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n3 VSS 0.02fF $ **FLOATING
C441 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n4 VSS 0.02fF $ **FLOATING
C442 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n5 VSS 0.02fF $ **FLOATING
C443 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n6 VSS 0.02fF $ **FLOATING
C444 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n7 VSS 0.02fF $ **FLOATING
C445 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n8 VSS 0.02fF $ **FLOATING
C446 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n9 VSS 0.02fF $ **FLOATING
C447 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n10 VSS 0.02fF $ **FLOATING
C448 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n11 VSS 0.02fF $ **FLOATING
C449 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t4 VSS 1.83fF
C450 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t2 VSS 0.21fF
C451 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t0 VSS 0.21fF
C452 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n12 VSS 1.57fF $ **FLOATING
C453 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t3 VSS 0.21fF
C454 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t6 VSS 0.21fF
C455 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n13 VSS 1.57fF $ **FLOATING
C456 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t7 VSS 0.21fF
C457 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t5 VSS 0.21fF
C458 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n14 VSS 1.57fF $ **FLOATING
C459 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t9 VSS 0.21fF
C460 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t1 VSS 0.21fF
C461 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n15 VSS 1.57fF $ **FLOATING
C462 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n16 VSS 0.00fF $ **FLOATING
C463 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n17 VSS 0.01fF $ **FLOATING
C464 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t8 VSS 0.21fF
C465 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n18 VSS 0.00fF $ **FLOATING
C466 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n19 VSS 0.00fF $ **FLOATING
C467 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n20 VSS 0.01fF $ **FLOATING
C468 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n21 VSS 0.00fF $ **FLOATING
C469 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n22 VSS 0.01fF $ **FLOATING
C470 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n23 VSS 0.00fF $ **FLOATING
C471 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n24 VSS 0.01fF $ **FLOATING
C472 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n25 VSS 0.00fF $ **FLOATING
C473 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n26 VSS 0.01fF $ **FLOATING
C474 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n27 VSS 0.00fF $ **FLOATING
C475 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n28 VSS 0.01fF $ **FLOATING
C476 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n29 VSS 0.01fF $ **FLOATING
C477 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n30 VSS 0.01fF $ **FLOATING
C478 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n31 VSS 0.63fF $ **FLOATING
C479 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n32 VSS 0.00fF $ **FLOATING
C480 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t13 VSS 1.33fF
C481 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t12 VSS 3.77fF
C482 sky130_asc_nfet_01v8_lvt_1_0/GATE VSS 0.60fF $ **FLOATING
C483 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n33 VSS 1.22fF $ **FLOATING
C484 sky130_asc_nfet_01v8_lvt_1_1/GATE VSS 0.13fF $ **FLOATING
C485 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t14 VSS 3.69fF
C486 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n34 VSS 3.15fF $ **FLOATING
C487 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n35 VSS 6.09fF $ **FLOATING
C488 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n36 VSS 0.01fF $ **FLOATING
C489 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n37 VSS 0.01fF $ **FLOATING
C490 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n38 VSS 1.61fF $ **FLOATING
C491 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n39 VSS 0.01fF $ **FLOATING
C492 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n40 VSS 0.03fF $ **FLOATING
C493 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n41 VSS 0.00fF $ **FLOATING
C494 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n42 VSS 0.01fF $ **FLOATING
C495 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n43 VSS 0.02fF $ **FLOATING
C496 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n44 VSS 0.00fF $ **FLOATING
C497 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n45 VSS 0.01fF $ **FLOATING
C498 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n46 VSS 0.02fF $ **FLOATING
C499 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n47 VSS 0.02fF $ **FLOATING
C500 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n48 VSS 0.00fF $ **FLOATING
C501 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n49 VSS 0.00fF $ **FLOATING
C502 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n50 VSS 0.01fF $ **FLOATING
C503 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n51 VSS 0.02fF $ **FLOATING
C504 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n52 VSS 0.02fF $ **FLOATING
C505 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n53 VSS 0.00fF $ **FLOATING
C506 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n54 VSS 0.01fF $ **FLOATING
C507 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n55 VSS 0.01fF $ **FLOATING
C508 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n56 VSS 0.02fF $ **FLOATING
C509 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n57 VSS 0.00fF $ **FLOATING
C510 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n58 VSS 0.01fF $ **FLOATING
C511 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n59 VSS 0.01fF $ **FLOATING
C512 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n60 VSS 0.02fF $ **FLOATING
C513 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n61 VSS 0.00fF $ **FLOATING
C514 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n62 VSS 0.01fF $ **FLOATING
C515 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n63 VSS 0.01fF $ **FLOATING
C516 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n64 VSS 0.01fF $ **FLOATING
C517 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n65 VSS 0.02fF $ **FLOATING
C518 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n66 VSS 0.00fF $ **FLOATING
C519 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n67 VSS 0.01fF $ **FLOATING
C520 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n68 VSS 0.01fF $ **FLOATING
C521 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n69 VSS 0.01fF $ **FLOATING
C522 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n70 VSS 0.00fF $ **FLOATING
C523 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n71 VSS 0.01fF $ **FLOATING
C524 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n72 VSS 0.01fF $ **FLOATING
C525 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n73 VSS 0.02fF $ **FLOATING
C526 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n74 VSS 0.01fF $ **FLOATING
C527 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n75 VSS 0.00fF $ **FLOATING
C528 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n76 VSS 0.01fF $ **FLOATING
C529 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n77 VSS 0.01fF $ **FLOATING
C530 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n78 VSS 0.02fF $ **FLOATING
C531 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n79 VSS 0.01fF $ **FLOATING
C532 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n80 VSS 0.00fF $ **FLOATING
C533 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n81 VSS 0.01fF $ **FLOATING
C534 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n82 VSS 0.01fF $ **FLOATING
C535 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n83 VSS 0.02fF $ **FLOATING
C536 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n84 VSS 0.01fF $ **FLOATING
C537 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n85 VSS 0.00fF $ **FLOATING
C538 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n86 VSS 0.01fF $ **FLOATING
C539 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n87 VSS 0.00fF $ **FLOATING
C540 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n88 VSS 0.02fF $ **FLOATING
C541 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n89 VSS 0.01fF $ **FLOATING
C542 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n90 VSS 0.02fF $ **FLOATING
C543 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n91 VSS 0.00fF $ **FLOATING
C544 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n92 VSS 0.00fF $ **FLOATING
C545 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n93 VSS 0.01fF $ **FLOATING
C546 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n94 VSS 0.00fF $ **FLOATING
C547 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n95 VSS 0.02fF $ **FLOATING
C548 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n96 VSS 0.01fF $ **FLOATING
C549 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n97 VSS 0.02fF $ **FLOATING
C550 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n98 VSS 0.00fF $ **FLOATING
C551 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n99 VSS 0.01fF $ **FLOATING
C552 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n100 VSS 0.00fF $ **FLOATING
C553 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n101 VSS 0.01fF $ **FLOATING
C554 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n102 VSS 0.02fF $ **FLOATING
C555 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n103 VSS 0.00fF $ **FLOATING
C556 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n104 VSS 0.01fF $ **FLOATING
C557 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n105 VSS 0.00fF $ **FLOATING
C558 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n106 VSS 0.01fF $ **FLOATING
C559 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n107 VSS 0.07fF $ **FLOATING
C560 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n108 VSS 0.34fF $ **FLOATING
C561 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n109 VSS 0.72fF $ **FLOATING
C562 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n110 VSS 0.65fF $ **FLOATING
C563 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n111 VSS 0.65fF $ **FLOATING
C564 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n112 VSS 0.65fF $ **FLOATING
C565 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t10 VSS 0.21fF
C566 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.t11 VSS 0.21fF
C567 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n113 VSS 1.57fF $ **FLOATING
C568 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n114 VSS 0.65fF $ **FLOATING
C569 sky130_asc_nfet_01v8_lvt_1_0/DRAIN.n115 VSS 0.49fF $ **FLOATING
C570 sky130_asc_pfet_01v8_lvt_12_1/DRAIN VSS 0.04fF $ **FLOATING
C571 vbg.t42 VSS 1.37fF
C572 vbg.t43 VSS 0.16fF
C573 vbg.t17 VSS 0.16fF
C574 vbg.n0 VSS 1.17fF $ **FLOATING
C575 vbg.t45 VSS 0.16fF
C576 vbg.t22 VSS 0.16fF
C577 vbg.n1 VSS 1.17fF $ **FLOATING
C578 vbg.t52 VSS 0.16fF
C579 vbg.t55 VSS 0.16fF
C580 vbg.n2 VSS 1.17fF $ **FLOATING
C581 vbg.t44 VSS 0.16fF
C582 vbg.t57 VSS 0.16fF
C583 vbg.n3 VSS 1.17fF $ **FLOATING
C584 vbg.t60 VSS 0.51fF
C585 sky130_asc_res_xhigh_po_2p85_1_8/Rin VSS 0.86fF $ **FLOATING
C586 vbg.n4 VSS 6.91fF $ **FLOATING
C587 vbg.t50 VSS 0.16fF
C588 vbg.t51 VSS 0.16fF
C589 vbg.n5 VSS 1.17fF $ **FLOATING
C590 vbg.t36 VSS 0.16fF
C591 vbg.t37 VSS 0.16fF
C592 vbg.n6 VSS 1.17fF $ **FLOATING
C593 vbg.t54 VSS 0.16fF
C594 vbg.t39 VSS 0.16fF
C595 vbg.n7 VSS 1.17fF $ **FLOATING
C596 vbg.t49 VSS 0.16fF
C597 vbg.t14 VSS 0.16fF
C598 vbg.n8 VSS 1.17fF $ **FLOATING
C599 vbg.t30 VSS 0.16fF
C600 vbg.t18 VSS 0.16fF
C601 vbg.n9 VSS 1.17fF $ **FLOATING
C602 vbg.t33 VSS 0.16fF
C603 vbg.t34 VSS 0.16fF
C604 vbg.n10 VSS 1.17fF $ **FLOATING
C605 vbg.t8 VSS 0.16fF
C606 vbg.t20 VSS 0.16fF
C607 vbg.n11 VSS 1.17fF $ **FLOATING
C608 vbg.t10 VSS 0.16fF
C609 vbg.t24 VSS 0.16fF
C610 vbg.n12 VSS 1.17fF $ **FLOATING
C611 vbg.t25 VSS 0.16fF
C612 vbg.t2 VSS 0.16fF
C613 vbg.n13 VSS 1.17fF $ **FLOATING
C614 vbg.t46 VSS 0.16fF
C615 vbg.t47 VSS 0.16fF
C616 vbg.n14 VSS 1.17fF $ **FLOATING
C617 vbg.t48 VSS 0.16fF
C618 vbg.t26 VSS 0.16fF
C619 vbg.n15 VSS 1.17fF $ **FLOATING
C620 vbg.t27 VSS 0.16fF
C621 vbg.t38 VSS 0.16fF
C622 vbg.n16 VSS 1.17fF $ **FLOATING
C623 vbg.t15 VSS 0.16fF
C624 vbg.t16 VSS 0.16fF
C625 vbg.n17 VSS 1.17fF $ **FLOATING
C626 vbg.t31 VSS 0.16fF
C627 vbg.t21 VSS 0.16fF
C628 vbg.n18 VSS 1.17fF $ **FLOATING
C629 vbg.t35 VSS 0.16fF
C630 vbg.t0 VSS 0.16fF
C631 vbg.n19 VSS 1.17fF $ **FLOATING
C632 vbg.t9 VSS 0.16fF
C633 vbg.t56 VSS 0.16fF
C634 vbg.n20 VSS 1.17fF $ **FLOATING
C635 vbg.t11 VSS 0.16fF
C636 vbg.t12 VSS 0.16fF
C637 vbg.n21 VSS 1.17fF $ **FLOATING
C638 vbg.t58 VSS 0.16fF
C639 vbg.t3 VSS 0.16fF
C640 vbg.n22 VSS 1.17fF $ **FLOATING
C641 vbg.t53 VSS 0.16fF
C642 vbg.t5 VSS 0.16fF
C643 vbg.n23 VSS 1.17fF $ **FLOATING
C644 vbg.t13 VSS 0.16fF
C645 vbg.t28 VSS 0.16fF
C646 vbg.n24 VSS 1.17fF $ **FLOATING
C647 vbg.t29 VSS 0.16fF
C648 vbg.t4 VSS 0.16fF
C649 vbg.n25 VSS 1.17fF $ **FLOATING
C650 vbg.t32 VSS 0.16fF
C651 vbg.t6 VSS 0.16fF
C652 vbg.n26 VSS 1.17fF $ **FLOATING
C653 vbg.t7 VSS 0.16fF
C654 vbg.t19 VSS 0.16fF
C655 vbg.n27 VSS 1.17fF $ **FLOATING
C656 vbg.t59 VSS 0.16fF
C657 vbg.t23 VSS 0.16fF
C658 vbg.n28 VSS 1.17fF $ **FLOATING
C659 vbg.t1 VSS 1.69fF
C660 vbg.n29 VSS 0.57fF $ **FLOATING
C661 vbg.n30 VSS 0.48fF $ **FLOATING
C662 vbg.n31 VSS 0.48fF $ **FLOATING
C663 vbg.n32 VSS 0.48fF $ **FLOATING
C664 vbg.n33 VSS 0.48fF $ **FLOATING
C665 vbg.n34 VSS 0.48fF $ **FLOATING
C666 vbg.n35 VSS 0.48fF $ **FLOATING
C667 vbg.n36 VSS 0.48fF $ **FLOATING
C668 vbg.n37 VSS 0.48fF $ **FLOATING
C669 vbg.n38 VSS 0.48fF $ **FLOATING
C670 vbg.n39 VSS 0.48fF $ **FLOATING
C671 vbg.n40 VSS 0.48fF $ **FLOATING
C672 vbg.n41 VSS 0.00fF $ **FLOATING
C673 vbg.n42 VSS 0.01fF $ **FLOATING
C674 vbg.t40 VSS 0.16fF
C675 vbg.n43 VSS 0.01fF $ **FLOATING
C676 vbg.n44 VSS 0.01fF $ **FLOATING
C677 vbg.n45 VSS 0.00fF $ **FLOATING
C678 vbg.n46 VSS 0.01fF $ **FLOATING
C679 vbg.n47 VSS 0.00fF $ **FLOATING
C680 vbg.n48 VSS 0.01fF $ **FLOATING
C681 vbg.n49 VSS 0.00fF $ **FLOATING
C682 vbg.n50 VSS 0.01fF $ **FLOATING
C683 vbg.n51 VSS 0.00fF $ **FLOATING
C684 vbg.n52 VSS 0.01fF $ **FLOATING
C685 vbg.n53 VSS 0.00fF $ **FLOATING
C686 vbg.n54 VSS 0.01fF $ **FLOATING
C687 vbg.n55 VSS 0.01fF $ **FLOATING
C688 vbg.t41 VSS 0.16fF
C689 vbg.n56 VSS 0.31fF $ **FLOATING
C690 vbg.n57 VSS 0.00fF $ **FLOATING
C691 vbg.n58 VSS 0.77fF $ **FLOATING
C692 vbg.n59 VSS 0.01fF $ **FLOATING
C693 vbg.n60 VSS 0.00fF $ **FLOATING
C694 vbg.n61 VSS 0.01fF $ **FLOATING
C695 vbg.n62 VSS 0.01fF $ **FLOATING
C696 vbg.n63 VSS 0.01fF $ **FLOATING
C697 vbg.n64 VSS 0.00fF $ **FLOATING
C698 vbg.n65 VSS 0.00fF $ **FLOATING
C699 vbg.n66 VSS 0.01fF $ **FLOATING
C700 vbg.n67 VSS 0.01fF $ **FLOATING
C701 vbg.n68 VSS 0.01fF $ **FLOATING
C702 vbg.n69 VSS 0.00fF $ **FLOATING
C703 vbg.n70 VSS 0.00fF $ **FLOATING
C704 vbg.n71 VSS 0.01fF $ **FLOATING
C705 vbg.n72 VSS 0.01fF $ **FLOATING
C706 vbg.n73 VSS 0.01fF $ **FLOATING
C707 vbg.n74 VSS 0.00fF $ **FLOATING
C708 vbg.n75 VSS 0.00fF $ **FLOATING
C709 vbg.n76 VSS 0.01fF $ **FLOATING
C710 vbg.n77 VSS 0.01fF $ **FLOATING
C711 vbg.n78 VSS 0.01fF $ **FLOATING
C712 vbg.n79 VSS 0.00fF $ **FLOATING
C713 vbg.n80 VSS 0.00fF $ **FLOATING
C714 vbg.n81 VSS 0.01fF $ **FLOATING
C715 vbg.n82 VSS 0.01fF $ **FLOATING
C716 vbg.n83 VSS 0.00fF $ **FLOATING
C717 vbg.n84 VSS 0.01fF $ **FLOATING
C718 vbg.n85 VSS 0.00fF $ **FLOATING
C719 vbg.n86 VSS 0.00fF $ **FLOATING
C720 vbg.n87 VSS 0.01fF $ **FLOATING
C721 vbg.n88 VSS 0.01fF $ **FLOATING
C722 vbg.n89 VSS 0.00fF $ **FLOATING
C723 vbg.n90 VSS 0.01fF $ **FLOATING
C724 vbg.n91 VSS 0.00fF $ **FLOATING
C725 vbg.n92 VSS 0.00fF $ **FLOATING
C726 vbg.n93 VSS 0.01fF $ **FLOATING
C727 vbg.n94 VSS 0.01fF $ **FLOATING
C728 vbg.n95 VSS 0.01fF $ **FLOATING
C729 vbg.n96 VSS 0.00fF $ **FLOATING
C730 vbg.n97 VSS 0.01fF $ **FLOATING
C731 vbg.n98 VSS 0.00fF $ **FLOATING
C732 vbg.n99 VSS 0.00fF $ **FLOATING
C733 vbg.n100 VSS 0.01fF $ **FLOATING
C734 vbg.n101 VSS 0.01fF $ **FLOATING
C735 vbg.n102 VSS 0.01fF $ **FLOATING
C736 vbg.n103 VSS 0.01fF $ **FLOATING
C737 vbg.n104 VSS 0.01fF $ **FLOATING
C738 vbg.n105 VSS 0.00fF $ **FLOATING
C739 vbg.n106 VSS 0.00fF $ **FLOATING
C740 vbg.n107 VSS 0.01fF $ **FLOATING
C741 vbg.n108 VSS 0.00fF $ **FLOATING
C742 vbg.n109 VSS 0.01fF $ **FLOATING
C743 vbg.n110 VSS 0.01fF $ **FLOATING
C744 vbg.n111 VSS 0.01fF $ **FLOATING
C745 vbg.n112 VSS 0.00fF $ **FLOATING
C746 vbg.n113 VSS 0.00fF $ **FLOATING
C747 vbg.n114 VSS 0.01fF $ **FLOATING
C748 vbg.n115 VSS 0.00fF $ **FLOATING
C749 vbg.n116 VSS 0.01fF $ **FLOATING
C750 vbg.n117 VSS 0.01fF $ **FLOATING
C751 vbg.n118 VSS 0.01fF $ **FLOATING
C752 vbg.n119 VSS 0.00fF $ **FLOATING
C753 vbg.n120 VSS 0.00fF $ **FLOATING
C754 vbg.n121 VSS 0.01fF $ **FLOATING
C755 vbg.n122 VSS 0.00fF $ **FLOATING
C756 vbg.n123 VSS 0.01fF $ **FLOATING
C757 vbg.n124 VSS 0.01fF $ **FLOATING
C758 vbg.n125 VSS 0.01fF $ **FLOATING
C759 vbg.n126 VSS 0.00fF $ **FLOATING
C760 vbg.n127 VSS 0.00fF $ **FLOATING
C761 vbg.n128 VSS 0.01fF $ **FLOATING
C762 vbg.n129 VSS 0.00fF $ **FLOATING
C763 vbg.n130 VSS 0.01fF $ **FLOATING
C764 vbg.n131 VSS 0.01fF $ **FLOATING
C765 vbg.n132 VSS 0.01fF $ **FLOATING
C766 vbg.n133 VSS 0.00fF $ **FLOATING
C767 vbg.n134 VSS 0.00fF $ **FLOATING
C768 vbg.n135 VSS 0.01fF $ **FLOATING
C769 vbg.n136 VSS 0.00fF $ **FLOATING
C770 vbg.n137 VSS 0.01fF $ **FLOATING
C771 vbg.n138 VSS 0.01fF $ **FLOATING
C772 vbg.n139 VSS 0.01fF $ **FLOATING
C773 vbg.n140 VSS 0.00fF $ **FLOATING
C774 vbg.n141 VSS 0.00fF $ **FLOATING
C775 vbg.n142 VSS 0.01fF $ **FLOATING
C776 vbg.n143 VSS 0.00fF $ **FLOATING
C777 vbg.n144 VSS 0.01fF $ **FLOATING
C778 vbg.n145 VSS 0.01fF $ **FLOATING
C779 vbg.n146 VSS 0.01fF $ **FLOATING
C780 vbg.n147 VSS 0.00fF $ **FLOATING
C781 vbg.n148 VSS 0.00fF $ **FLOATING
C782 vbg.n149 VSS 0.01fF $ **FLOATING
C783 vbg.n150 VSS 0.00fF $ **FLOATING
C784 vbg.n151 VSS 0.01fF $ **FLOATING
C785 vbg.n152 VSS 0.01fF $ **FLOATING
C786 vbg.n153 VSS 0.01fF $ **FLOATING
C787 vbg.n154 VSS 0.00fF $ **FLOATING
C788 vbg.n155 VSS 0.04fF $ **FLOATING
C789 vbg.n156 VSS 0.03fF $ **FLOATING
C790 vbg.n157 VSS 0.48fF $ **FLOATING
C791 vbg.n158 VSS 0.48fF $ **FLOATING
C792 vbg.n159 VSS 0.48fF $ **FLOATING
C793 vbg.n160 VSS 0.48fF $ **FLOATING
C794 vbg.n161 VSS 0.48fF $ **FLOATING
C795 vbg.n162 VSS 0.48fF $ **FLOATING
C796 vbg.n163 VSS 0.48fF $ **FLOATING
C797 vbg.n164 VSS 0.48fF $ **FLOATING
C798 vbg.n165 VSS 0.48fF $ **FLOATING
C799 vbg.n166 VSS 0.48fF $ **FLOATING
C800 vbg.n167 VSS 0.48fF $ **FLOATING
C801 vbg.n168 VSS 0.48fF $ **FLOATING
C802 vbg.n169 VSS 0.43fF $ **FLOATING
C803 vbg.n170 VSS 2.38fF $ **FLOATING
C804 vbg.n171 VSS 0.31fF $ **FLOATING
C805 vbg.n172 VSS 0.48fF $ **FLOATING
C806 vbg.n173 VSS 0.48fF $ **FLOATING
C807 vbg.n174 VSS 0.48fF $ **FLOATING
C808 vbg.n175 VSS 0.37fF $ **FLOATING
C809 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t16 VSS 0.08fF
C810 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t10 VSS 0.08fF
C811 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n0 VSS 0.58fF $ **FLOATING
C812 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t18 VSS 0.08fF
C813 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t20 VSS 0.08fF
C814 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n1 VSS 0.58fF $ **FLOATING
C815 sky130_asc_pfet_01v8_lvt_6_1/GATE VSS 0.04fF $ **FLOATING
C816 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t13 VSS 1.87fF
C817 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n2 VSS 0.34fF $ **FLOATING
C818 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n3 VSS 0.08fF $ **FLOATING
C819 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t15 VSS 1.87fF
C820 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n4 VSS 0.42fF $ **FLOATING
C821 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n5 VSS 0.07fF $ **FLOATING
C822 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n6 VSS 0.10fF $ **FLOATING
C823 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n7 VSS 0.07fF $ **FLOATING
C824 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n8 VSS 0.10fF $ **FLOATING
C825 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t9 VSS 1.87fF
C826 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n9 VSS 0.42fF $ **FLOATING
C827 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n10 VSS 0.07fF $ **FLOATING
C828 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n11 VSS 0.10fF $ **FLOATING
C829 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t17 VSS 1.87fF
C830 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n12 VSS 0.42fF $ **FLOATING
C831 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n13 VSS 0.07fF $ **FLOATING
C832 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n14 VSS 0.10fF $ **FLOATING
C833 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t19 VSS 1.87fF
C834 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n15 VSS 0.42fF $ **FLOATING
C835 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n16 VSS 0.07fF $ **FLOATING
C836 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n17 VSS 0.10fF $ **FLOATING
C837 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t11 VSS 1.87fF
C838 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n18 VSS 0.50fF $ **FLOATING
C839 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n19 VSS 0.09fF $ **FLOATING
C840 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n20 VSS 0.00fF $ **FLOATING
C841 sky130_asc_pfet_01v8_lvt_6_0/GATE VSS 0.04fF $ **FLOATING
C842 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n21 VSS 0.03fF $ **FLOATING
C843 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n22 VSS 0.00fF $ **FLOATING
C844 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t22 VSS 1.87fF
C845 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n23 VSS -0.01fF $ **FLOATING
C846 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n24 VSS 0.34fF $ **FLOATING
C847 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n25 VSS 0.00fF $ **FLOATING
C848 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t21 VSS 1.87fF
C849 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n26 VSS 0.42fF $ **FLOATING
C850 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n27 VSS 0.07fF $ **FLOATING
C851 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t23 VSS 2.01fF
C852 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n28 VSS 0.57fF $ **FLOATING
C853 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t24 VSS 1.87fF
C854 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n29 VSS 0.45fF $ **FLOATING
C855 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n30 VSS 0.07fF $ **FLOATING
C856 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n31 VSS 0.15fF $ **FLOATING
C857 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t25 VSS 1.87fF
C858 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n32 VSS 0.42fF $ **FLOATING
C859 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n33 VSS 0.07fF $ **FLOATING
C860 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n34 VSS 0.10fF $ **FLOATING
C861 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t26 VSS 1.87fF
C862 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n35 VSS 0.42fF $ **FLOATING
C863 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n36 VSS 0.07fF $ **FLOATING
C864 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n37 VSS 0.10fF $ **FLOATING
C865 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n38 VSS 0.10fF $ **FLOATING
C866 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n39 VSS 0.05fF $ **FLOATING
C867 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n40 VSS 0.01fF $ **FLOATING
C868 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n41 VSS 0.25fF $ **FLOATING
C869 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t2 VSS 0.05fF
C870 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t0 VSS 0.05fF
C871 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n42 VSS 0.35fF $ **FLOATING
C872 sky130_asc_nfet_01v8_lvt_9_2/DRAIN VSS 0.07fF $ **FLOATING
C873 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n43 VSS 0.08fF $ **FLOATING
C874 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t1 VSS 0.05fF
C875 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t4 VSS 0.05fF
C876 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n44 VSS 0.35fF $ **FLOATING
C877 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t5 VSS 0.05fF
C878 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t6 VSS 0.05fF
C879 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n45 VSS 0.35fF $ **FLOATING
C880 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t7 VSS 0.05fF
C881 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t8 VSS 0.05fF
C882 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n46 VSS 0.35fF $ **FLOATING
C883 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t3 VSS 0.55fF
C884 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n47 VSS 0.27fF $ **FLOATING
C885 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n48 VSS 0.24fF $ **FLOATING
C886 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n49 VSS 0.22fF $ **FLOATING
C887 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n50 VSS 0.11fF $ **FLOATING
C888 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n51 VSS 1.08fF $ **FLOATING
C889 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n52 VSS 1.00fF $ **FLOATING
C890 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t12 VSS 0.16fF
C891 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n53 VSS 0.68fF $ **FLOATING
C892 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n54 VSS 0.27fF $ **FLOATING
C893 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n55 VSS 0.24fF $ **FLOATING
C894 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.t14 VSS 0.67fF
C895 sky130_asc_pfet_01v8_lvt_6_1/DRAIN.n56 VSS 0.18fF $ **FLOATING
C896 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t8 VSS 1.05fF
C897 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t6 VSS 0.11fF
C898 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t7 VSS 0.11fF
C899 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n0 VSS 0.85fF $ **FLOATING
C900 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t18 VSS 1.03fF
C901 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n1 VSS 1.69fF $ **FLOATING
C902 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t15 VSS 1.05fF
C903 sky130_asc_nfet_01v8_lvt_9_2/SOURCE VSS 0.30fF $ **FLOATING
C904 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t17 VSS 0.11fF
C905 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t16 VSS 0.11fF
C906 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n2 VSS 0.85fF $ **FLOATING
C907 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t9 VSS 0.11fF
C908 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t11 VSS 0.11fF
C909 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n3 VSS 0.85fF $ **FLOATING
C910 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t12 VSS 0.11fF
C911 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t13 VSS 0.11fF
C912 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n4 VSS 0.85fF $ **FLOATING
C913 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t14 VSS 0.11fF
C914 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t10 VSS 0.11fF
C915 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n5 VSS 1.21fF $ **FLOATING
C916 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n6 VSS 0.80fF $ **FLOATING
C917 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n7 VSS 0.57fF $ **FLOATING
C918 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n8 VSS 0.39fF $ **FLOATING
C919 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n9 VSS 0.71fF $ **FLOATING
C920 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n10 VSS 2.43fF $ **FLOATING
C921 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t1 VSS 0.11fF
C922 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t2 VSS 0.11fF
C923 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n11 VSS 0.85fF $ **FLOATING
C924 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t3 VSS 0.11fF
C925 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t4 VSS 0.11fF
C926 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n12 VSS 0.85fF $ **FLOATING
C927 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t5 VSS 0.11fF
C928 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.t0 VSS 0.11fF
C929 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n13 VSS 1.21fF $ **FLOATING
C930 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n14 VSS 0.80fF $ **FLOATING
C931 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n15 VSS 0.57fF $ **FLOATING
C932 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n16 VSS 0.28fF $ **FLOATING
C933 sky130_asc_nfet_01v8_lvt_1_1/DRAIN.n17 VSS 0.32fF $ **FLOATING
C934 sky130_asc_nfet_01v8_lvt_9_1/SOURCE VSS 0.37fF $ **FLOATING
C935 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t48 VSS 1.11fF
C936 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t20 VSS 0.13fF
C937 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t32 VSS 0.13fF
C938 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n0 VSS 0.95fF $ **FLOATING
C939 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t0 VSS 0.42fF
C940 sky130_asc_res_xhigh_po_2p85_1_18/Rin VSS 0.70fF $ **FLOATING
C941 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n1 VSS 3.70fF $ **FLOATING
C942 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t61 VSS 0.42fF
C943 sky130_asc_res_xhigh_po_2p85_1_20/Rin VSS 0.70fF $ **FLOATING
C944 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n2 VSS 4.01fF $ **FLOATING
C945 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n3 VSS 0.64fF $ **FLOATING
C946 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t58 VSS 0.13fF
C947 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t59 VSS 0.13fF
C948 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n4 VSS 0.65fF $ **FLOATING
C949 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n5 VSS 0.58fF $ **FLOATING
C950 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t54 VSS 0.13fF
C951 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t55 VSS 0.13fF
C952 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n6 VSS 0.95fF $ **FLOATING
C953 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t56 VSS 0.13fF
C954 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t57 VSS 0.13fF
C955 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n7 VSS 0.95fF $ **FLOATING
C956 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t43 VSS 0.13fF
C957 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t44 VSS 0.13fF
C958 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n8 VSS 0.95fF $ **FLOATING
C959 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t26 VSS 0.13fF
C960 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t46 VSS 0.13fF
C961 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n9 VSS 0.95fF $ **FLOATING
C962 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t53 VSS 0.13fF
C963 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t29 VSS 0.13fF
C964 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n10 VSS 0.95fF $ **FLOATING
C965 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t40 VSS 0.13fF
C966 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t19 VSS 0.13fF
C967 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n11 VSS 0.95fF $ **FLOATING
C968 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t41 VSS 0.13fF
C969 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t22 VSS 0.13fF
C970 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n12 VSS 0.95fF $ **FLOATING
C971 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t23 VSS 0.13fF
C972 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t34 VSS 0.13fF
C973 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n13 VSS 0.95fF $ **FLOATING
C974 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t2 VSS 0.13fF
C975 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t36 VSS 0.13fF
C976 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n14 VSS 0.95fF $ **FLOATING
C977 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t42 VSS 0.13fF
C978 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t50 VSS 0.13fF
C979 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n15 VSS 0.95fF $ **FLOATING
C980 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t51 VSS 0.13fF
C981 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t35 VSS 0.13fF
C982 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n16 VSS 0.95fF $ **FLOATING
C983 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t52 VSS 0.13fF
C984 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t38 VSS 0.13fF
C985 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n17 VSS 0.95fF $ **FLOATING
C986 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t45 VSS 0.13fF
C987 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t16 VSS 0.13fF
C988 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n18 VSS 0.95fF $ **FLOATING
C989 sky130_asc_nfet_01v8_lvt_9_2/GATE VSS 0.06fF $ **FLOATING
C990 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t68 VSS 2.07fF
C991 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n19 VSS 0.32fF $ **FLOATING
C992 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t70 VSS 2.04fF
C993 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n20 VSS 0.58fF $ **FLOATING
C994 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t69 VSS 2.04fF
C995 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n21 VSS 0.59fF $ **FLOATING
C996 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t66 VSS 2.04fF
C997 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n22 VSS 0.58fF $ **FLOATING
C998 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t62 VSS 2.04fF
C999 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n23 VSS 0.52fF $ **FLOATING
C1000 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t67 VSS 2.20fF
C1001 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n24 VSS 0.67fF $ **FLOATING
C1002 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n25 VSS 0.11fF $ **FLOATING
C1003 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n26 VSS 0.23fF $ **FLOATING
C1004 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t63 VSS 2.04fF
C1005 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n27 VSS 0.46fF $ **FLOATING
C1006 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n28 VSS 0.11fF $ **FLOATING
C1007 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n29 VSS 0.16fF $ **FLOATING
C1008 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t64 VSS 2.04fF
C1009 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n30 VSS 0.46fF $ **FLOATING
C1010 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n31 VSS 0.11fF $ **FLOATING
C1011 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n32 VSS 0.16fF $ **FLOATING
C1012 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t65 VSS 2.04fF
C1013 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n33 VSS 0.46fF $ **FLOATING
C1014 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n34 VSS 0.11fF $ **FLOATING
C1015 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n35 VSS 0.16fF $ **FLOATING
C1016 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n36 VSS 0.16fF $ **FLOATING
C1017 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n37 VSS 0.16fF $ **FLOATING
C1018 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n38 VSS 0.16fF $ **FLOATING
C1019 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n39 VSS 0.11fF $ **FLOATING
C1020 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n40 VSS 1.15fF $ **FLOATING
C1021 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t27 VSS 0.13fF
C1022 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t47 VSS 0.13fF
C1023 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n41 VSS 0.95fF $ **FLOATING
C1024 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t30 VSS 0.13fF
C1025 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t31 VSS 0.13fF
C1026 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n42 VSS 0.95fF $ **FLOATING
C1027 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t8 VSS 0.13fF
C1028 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t9 VSS 0.13fF
C1029 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n43 VSS 0.95fF $ **FLOATING
C1030 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t12 VSS 0.13fF
C1031 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t13 VSS 0.13fF
C1032 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n44 VSS 0.95fF $ **FLOATING
C1033 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t24 VSS 0.13fF
C1034 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t3 VSS 0.13fF
C1035 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n45 VSS 0.95fF $ **FLOATING
C1036 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t4 VSS 0.13fF
C1037 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t5 VSS 0.13fF
C1038 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n46 VSS 0.95fF $ **FLOATING
C1039 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t6 VSS 0.13fF
C1040 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t15 VSS 0.13fF
C1041 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n47 VSS 0.95fF $ **FLOATING
C1042 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t25 VSS 0.13fF
C1043 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t37 VSS 0.13fF
C1044 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n48 VSS 0.95fF $ **FLOATING
C1045 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t28 VSS 0.13fF
C1046 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t39 VSS 0.13fF
C1047 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n49 VSS 0.95fF $ **FLOATING
C1048 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t7 VSS 0.13fF
C1049 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t17 VSS 0.13fF
C1050 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n50 VSS 0.95fF $ **FLOATING
C1051 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t18 VSS 0.13fF
C1052 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t21 VSS 0.13fF
C1053 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n51 VSS 0.95fF $ **FLOATING
C1054 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t33 VSS 0.13fF
C1055 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t1 VSS 0.13fF
C1056 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n52 VSS 0.95fF $ **FLOATING
C1057 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t10 VSS 0.13fF
C1058 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t11 VSS 0.13fF
C1059 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n53 VSS 0.95fF $ **FLOATING
C1060 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t14 VSS 1.37fF
C1061 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n54 VSS 0.46fF $ **FLOATING
C1062 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n55 VSS 0.39fF $ **FLOATING
C1063 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n56 VSS 0.39fF $ **FLOATING
C1064 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n57 VSS 0.39fF $ **FLOATING
C1065 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n58 VSS 0.39fF $ **FLOATING
C1066 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n59 VSS 0.39fF $ **FLOATING
C1067 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n60 VSS 0.39fF $ **FLOATING
C1068 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n61 VSS 0.39fF $ **FLOATING
C1069 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n62 VSS 0.39fF $ **FLOATING
C1070 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n63 VSS 0.39fF $ **FLOATING
C1071 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n64 VSS 0.39fF $ **FLOATING
C1072 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n65 VSS 0.39fF $ **FLOATING
C1073 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n66 VSS 0.37fF $ **FLOATING
C1074 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n67 VSS 1.27fF $ **FLOATING
C1075 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n68 VSS 0.23fF $ **FLOATING
C1076 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n69 VSS 0.39fF $ **FLOATING
C1077 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n70 VSS 0.39fF $ **FLOATING
C1078 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n71 VSS 0.39fF $ **FLOATING
C1079 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n72 VSS 0.39fF $ **FLOATING
C1080 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n73 VSS 0.39fF $ **FLOATING
C1081 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n74 VSS 0.39fF $ **FLOATING
C1082 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n75 VSS 0.39fF $ **FLOATING
C1083 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n76 VSS 0.39fF $ **FLOATING
C1084 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n77 VSS 0.39fF $ **FLOATING
C1085 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n78 VSS 0.39fF $ **FLOATING
C1086 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n79 VSS 0.39fF $ **FLOATING
C1087 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n80 VSS 0.39fF $ **FLOATING
C1088 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t60 VSS 0.13fF
C1089 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.t49 VSS 0.13fF
C1090 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n81 VSS 0.95fF $ **FLOATING
C1091 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n82 VSS 0.39fF $ **FLOATING
C1092 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n83 VSS 0.39fF $ **FLOATING
C1093 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n84 VSS 0.39fF $ **FLOATING
C1094 sky130_asc_pfet_01v8_lvt_60_1/DRAIN.n85 VSS 0.30fF $ **FLOATING
C1095 sky130_asc_res_xhigh_po_2p85_2_1/VPWR VSS 1.48fF $ **FLOATING
C1096 VDD.n0 VSS 108.44fF $ **FLOATING
C1097 sky130_asc_res_xhigh_po_2p85_1_3/VPWR VSS 0.92fF $ **FLOATING
C1098 sky130_asc_res_xhigh_po_2p85_1_4/VPWR VSS 0.92fF $ **FLOATING
C1099 sky130_asc_nfet_01v8_lvt_9_0/VPWR VSS 1.07fF $ **FLOATING
C1100 sky130_asc_pfet_01v8_lvt_12_0/VPWR VSS 0.03fF $ **FLOATING
C1101 VDD.n1 VSS 0.11fF $ **FLOATING
C1102 VDD.n2 VSS 0.08fF $ **FLOATING
C1103 VDD.n3 VSS 0.45fF $ **FLOATING
C1104 sky130_asc_res_xhigh_po_2p85_1_7/VPWR VSS 0.82fF $ **FLOATING
C1105 sky130_asc_pfet_01v8_lvt_60_2/VPWR VSS 0.03fF $ **FLOATING
C1106 VDD.n4 VSS 0.11fF $ **FLOATING
C1107 VDD.n5 VSS 0.08fF $ **FLOATING
C1108 VDD.n6 VSS 0.25fF $ **FLOATING
C1109 sky130_asc_cap_mim_m3_1_2/VPWR VSS 0.81fF $ **FLOATING
C1110 VDD.n8 VSS 0.03fF $ **FLOATING
C1111 VDD.n9 VSS 0.03fF $ **FLOATING
C1112 VDD.n10 VSS 0.03fF $ **FLOATING
C1113 VDD.n11 VSS 0.03fF $ **FLOATING
C1114 VDD.t119 VSS 0.04fF
C1115 VDD.t206 VSS 0.04fF
C1116 VDD.n13 VSS 0.29fF $ **FLOATING
C1117 VDD.t255 VSS 0.04fF
C1118 VDD.t306 VSS 0.04fF
C1119 VDD.n14 VSS 0.29fF $ **FLOATING
C1120 VDD.t243 VSS 0.04fF
C1121 VDD.t29 VSS 0.04fF
C1122 VDD.n15 VSS 0.29fF $ **FLOATING
C1123 VDD.t329 VSS 0.04fF
C1124 VDD.t148 VSS 0.04fF
C1125 VDD.n16 VSS 0.29fF $ **FLOATING
C1126 VDD.t320 VSS 0.04fF
C1127 VDD.t285 VSS 0.04fF
C1128 VDD.n17 VSS 0.29fF $ **FLOATING
C1129 VDD.t53 VSS 0.04fF
C1130 VDD.t277 VSS 0.04fF
C1131 VDD.n18 VSS 0.29fF $ **FLOATING
C1132 VDD.t177 VSS 0.04fF
C1133 VDD.t181 VSS 0.04fF
C1134 VDD.n19 VSS 0.29fF $ **FLOATING
C1135 VDD.t139 VSS 0.04fF
C1136 VDD.t160 VSS 0.04fF
C1137 VDD.n20 VSS 0.29fF $ **FLOATING
C1138 VDD.t210 VSS 0.04fF
C1139 VDD.t271 VSS 0.04fF
C1140 VDD.n21 VSS 0.29fF $ **FLOATING
C1141 VDD.t150 VSS 0.04fF
C1142 VDD.t218 VSS 0.04fF
C1143 VDD.n22 VSS 0.29fF $ **FLOATING
C1144 VDD.t299 VSS 0.04fF
C1145 VDD.t197 VSS 0.04fF
C1146 VDD.n23 VSS 0.29fF $ **FLOATING
C1147 VDD.t363 VSS 0.04fF
C1148 VDD.t295 VSS 0.04fF
C1149 VDD.n24 VSS 0.29fF $ **FLOATING
C1150 VDD.t27 VSS 0.04fF
C1151 VDD.t287 VSS 0.04fF
C1152 VDD.n25 VSS 0.29fF $ **FLOATING
C1153 VDD.t322 VSS 0.04fF
C1154 VDD.t355 VSS 0.04fF
C1155 VDD.n26 VSS 0.29fF $ **FLOATING
C1156 VDD.t311 VSS 0.04fF
C1157 VDD.t389 VSS 0.04fF
C1158 VDD.n27 VSS 0.29fF $ **FLOATING
C1159 VDD.t373 VSS 0.04fF
C1160 VDD.t375 VSS 0.04fF
C1161 VDD.n28 VSS 0.29fF $ **FLOATING
C1162 VDD.t316 VSS 0.04fF
C1163 VDD.t339 VSS 0.04fF
C1164 VDD.n29 VSS 0.29fF $ **FLOATING
C1165 VDD.t308 VSS 0.04fF
C1166 VDD.t129 VSS 0.04fF
C1167 VDD.n30 VSS 0.29fF $ **FLOATING
C1168 VDD.t257 VSS 0.04fF
C1169 VDD.t261 VSS 0.04fF
C1170 VDD.n31 VSS 0.29fF $ **FLOATING
C1171 VDD.t245 VSS 0.04fF
C1172 VDD.t337 VSS 0.04fF
C1173 VDD.n32 VSS 0.29fF $ **FLOATING
C1174 VDD.t291 VSS 0.04fF
C1175 VDD.t331 VSS 0.04fF
C1176 VDD.n33 VSS 0.29fF $ **FLOATING
C1177 VDD.t359 VSS 0.04fF
C1178 VDD.t393 VSS 0.04fF
C1179 VDD.n34 VSS 0.29fF $ **FLOATING
C1180 VDD.t353 VSS 0.04fF
C1181 VDD.t281 VSS 0.04fF
C1182 VDD.n35 VSS 0.29fF $ **FLOATING
C1183 VDD.t415 VSS 0.04fF
C1184 VDD.t345 VSS 0.04fF
C1185 VDD.n36 VSS 0.29fF $ **FLOATING
C1186 VDD.t409 VSS 0.04fF
C1187 VDD.t411 VSS 0.04fF
C1188 VDD.n37 VSS 0.29fF $ **FLOATING
C1189 VDD.t371 VSS 0.04fF
C1190 VDD.t407 VSS 0.04fF
C1191 VDD.n38 VSS 0.29fF $ **FLOATING
C1192 VDD.t429 VSS 0.04fF
C1193 VDD.t433 VSS 0.04fF
C1194 VDD.n39 VSS 0.29fF $ **FLOATING
C1195 VDD.t301 VSS 0.04fF
C1196 VDD.t425 VSS 0.04fF
C1197 VDD.n40 VSS 0.29fF $ **FLOATING
C1198 VDD.t367 VSS 0.04fF
C1199 VDD.t251 VSS 0.04fF
C1200 VDD.n41 VSS 0.29fF $ **FLOATING
C1201 sky130_asc_pfet_01v8_lvt_60_1/SOURCE VSS 0.02fF $ **FLOATING
C1202 VDD.n42 VSS 0.06fF $ **FLOATING
C1203 VDD.n43 VSS 0.08fF $ **FLOATING
C1204 VDD.n44 VSS 0.08fF $ **FLOATING
C1205 VDD.n45 VSS 0.08fF $ **FLOATING
C1206 VDD.n46 VSS 0.08fF $ **FLOATING
C1207 VDD.n47 VSS 0.08fF $ **FLOATING
C1208 VDD.n48 VSS 0.08fF $ **FLOATING
C1209 VDD.n49 VSS 0.08fF $ **FLOATING
C1210 VDD.n50 VSS 0.08fF $ **FLOATING
C1211 VDD.n51 VSS 0.08fF $ **FLOATING
C1212 VDD.n52 VSS 0.08fF $ **FLOATING
C1213 VDD.n53 VSS 0.08fF $ **FLOATING
C1214 VDD.n54 VSS 0.08fF $ **FLOATING
C1215 VDD.n55 VSS 0.08fF $ **FLOATING
C1216 VDD.n56 VSS 0.08fF $ **FLOATING
C1217 VDD.n57 VSS 0.08fF $ **FLOATING
C1218 VDD.n58 VSS 0.08fF $ **FLOATING
C1219 VDD.n59 VSS 0.08fF $ **FLOATING
C1220 VDD.n60 VSS 0.08fF $ **FLOATING
C1221 VDD.n61 VSS 0.08fF $ **FLOATING
C1222 VDD.n62 VSS 0.08fF $ **FLOATING
C1223 VDD.n63 VSS 0.08fF $ **FLOATING
C1224 VDD.n64 VSS 0.08fF $ **FLOATING
C1225 VDD.n65 VSS 0.08fF $ **FLOATING
C1226 VDD.n66 VSS 0.08fF $ **FLOATING
C1227 VDD.n67 VSS 0.08fF $ **FLOATING
C1228 VDD.n68 VSS 0.08fF $ **FLOATING
C1229 VDD.n69 VSS 0.08fF $ **FLOATING
C1230 VDD.n70 VSS 0.09fF $ **FLOATING
C1231 VDD.t212 VSS 0.04fF
C1232 VDD.t222 VSS 0.04fF
C1233 VDD.n71 VSS 0.20fF $ **FLOATING
C1234 VDD.n72 VSS 0.14fF $ **FLOATING
C1235 VDD.n73 VSS 0.00fF $ **FLOATING
C1236 VDD.t58 VSS 2.41fF
C1237 VDD.t15 VSS 2.19fF
C1238 VDD.t10 VSS 2.19fF
C1239 VDD.t334 VSS 2.19fF
C1240 VDD.t98 VSS 1.61fF
C1241 sky130_asc_cap_mim_m3_1_2/Cin VSS 0.03fF $ **FLOATING
C1242 VDD.t325 VSS 1.92fF
C1243 VDD.t22 VSS 2.19fF
C1244 VDD.t142 VSS 2.19fF
C1245 VDD.t56 VSS 2.19fF
C1246 VDD.t63 VSS 1.56fF
C1247 VDD.n74 VSS 1.24fF $ **FLOATING
C1248 VDD.n75 VSS 0.04fF $ **FLOATING
C1249 VDD.n76 VSS 0.63fF $ **FLOATING
C1250 VDD.n77 VSS 0.05fF $ **FLOATING
C1251 VDD.n78 VSS 0.00fF $ **FLOATING
C1252 VDD.n79 VSS 0.04fF $ **FLOATING
C1253 VDD.n80 VSS 0.81fF $ **FLOATING
C1254 sky130_asc_pfet_01v8_lvt_60_1/VPWR VSS 0.03fF $ **FLOATING
C1255 VDD.n81 VSS 0.11fF $ **FLOATING
C1256 VDD.n82 VSS 0.08fF $ **FLOATING
C1257 VDD.n83 VSS 0.79fF $ **FLOATING
C1258 VDD.n84 VSS 0.09fF $ **FLOATING
C1259 VDD.n85 VSS 0.05fF $ **FLOATING
C1260 VDD.n86 VSS 0.06fF $ **FLOATING
C1261 VDD.t118 VSS 1.58fF
C1262 VDD.t205 VSS 1.05fF
C1263 VDD.t221 VSS 2.01fF
C1264 VDD.t211 VSS 1.32fF
C1265 VDD.n87 VSS 0.79fF $ **FLOATING
C1266 VDD.n88 VSS 0.05fF $ **FLOATING
C1267 VDD.n89 VSS 0.04fF $ **FLOATING
C1268 VDD.n90 VSS 0.10fF $ **FLOATING
C1269 VDD.n91 VSS 0.04fF $ **FLOATING
C1270 VDD.n92 VSS 0.10fF $ **FLOATING
C1271 VDD.n93 VSS 0.05fF $ **FLOATING
C1272 VDD.n94 VSS 0.10fF $ **FLOATING
C1273 VDD.t254 VSS 1.17fF
C1274 VDD.t305 VSS 1.19fF
C1275 VDD.n95 VSS 0.79fF $ **FLOATING
C1276 VDD.n96 VSS 0.06fF $ **FLOATING
C1277 VDD.n97 VSS 0.04fF $ **FLOATING
C1278 VDD.n98 VSS 0.10fF $ **FLOATING
C1279 VDD.n99 VSS 0.04fF $ **FLOATING
C1280 VDD.n100 VSS 0.10fF $ **FLOATING
C1281 VDD.n101 VSS 0.05fF $ **FLOATING
C1282 VDD.n102 VSS 0.10fF $ **FLOATING
C1283 VDD.n103 VSS 0.04fF $ **FLOATING
C1284 VDD.n104 VSS 0.10fF $ **FLOATING
C1285 VDD.t147 VSS 1.30fF
C1286 VDD.t28 VSS 1.58fF
C1287 VDD.t242 VSS 1.07fF
C1288 VDD.n105 VSS 0.79fF $ **FLOATING
C1289 VDD.n106 VSS 0.06fF $ **FLOATING
C1290 VDD.n107 VSS 0.03fF $ **FLOATING
C1291 VDD.n108 VSS 0.10fF $ **FLOATING
C1292 VDD.n109 VSS 0.05fF $ **FLOATING
C1293 VDD.n110 VSS 0.10fF $ **FLOATING
C1294 VDD.n111 VSS 0.05fF $ **FLOATING
C1295 VDD.n112 VSS 0.10fF $ **FLOATING
C1296 VDD.t319 VSS 1.43fF
C1297 VDD.t328 VSS 1.58fF
C1298 VDD.t284 VSS 0.94fF
C1299 VDD.n113 VSS 0.79fF $ **FLOATING
C1300 VDD.n114 VSS 0.05fF $ **FLOATING
C1301 VDD.n115 VSS 0.04fF $ **FLOATING
C1302 VDD.n116 VSS 0.10fF $ **FLOATING
C1303 VDD.n117 VSS 0.05fF $ **FLOATING
C1304 VDD.n118 VSS 0.10fF $ **FLOATING
C1305 VDD.n119 VSS 0.05fF $ **FLOATING
C1306 VDD.n120 VSS 0.10fF $ **FLOATING
C1307 VDD.t180 VSS 1.56fF
C1308 VDD.t276 VSS 1.58fF
C1309 VDD.t52 VSS 0.81fF
C1310 VDD.n121 VSS 0.79fF $ **FLOATING
C1311 VDD.n122 VSS 0.05fF $ **FLOATING
C1312 VDD.n123 VSS 0.04fF $ **FLOATING
C1313 VDD.n124 VSS 0.10fF $ **FLOATING
C1314 VDD.n125 VSS 0.04fF $ **FLOATING
C1315 VDD.n126 VSS 0.10fF $ **FLOATING
C1316 VDD.n127 VSS 0.05fF $ **FLOATING
C1317 VDD.n128 VSS 0.10fF $ **FLOATING
C1318 VDD.t138 VSS 1.58fF
C1319 VDD.t159 VSS 0.89fF
C1320 VDD.t176 VSS 1.47fF
C1321 VDD.n129 VSS 0.79fF $ **FLOATING
C1322 VDD.n130 VSS 0.06fF $ **FLOATING
C1323 VDD.n131 VSS 0.04fF $ **FLOATING
C1324 VDD.n132 VSS 0.10fF $ **FLOATING
C1325 VDD.n133 VSS 0.04fF $ **FLOATING
C1326 VDD.n134 VSS 0.10fF $ **FLOATING
C1327 VDD.n135 VSS 0.05fF $ **FLOATING
C1328 VDD.n136 VSS 0.10fF $ **FLOATING
C1329 VDD.n137 VSS 0.04fF $ **FLOATING
C1330 VDD.n138 VSS 0.10fF $ **FLOATING
C1331 VDD.t217 VSS 1.58fF
C1332 VDD.t209 VSS 1.02fF
C1333 VDD.t270 VSS 1.35fF
C1334 VDD.n139 VSS 0.79fF $ **FLOATING
C1335 VDD.n140 VSS 0.06fF $ **FLOATING
C1336 VDD.n141 VSS 0.03fF $ **FLOATING
C1337 VDD.n142 VSS 0.10fF $ **FLOATING
C1338 VDD.n143 VSS 0.05fF $ **FLOATING
C1339 VDD.n144 VSS 0.10fF $ **FLOATING
C1340 VDD.n145 VSS 0.05fF $ **FLOATING
C1341 VDD.n146 VSS 0.10fF $ **FLOATING
C1342 VDD.t196 VSS 1.15fF
C1343 VDD.t149 VSS 1.22fF
C1344 VDD.n147 VSS 0.79fF $ **FLOATING
C1345 VDD.n148 VSS 0.05fF $ **FLOATING
C1346 VDD.n149 VSS 0.04fF $ **FLOATING
C1347 VDD.n150 VSS 0.10fF $ **FLOATING
C1348 VDD.n151 VSS 0.05fF $ **FLOATING
C1349 VDD.n152 VSS 0.10fF $ **FLOATING
C1350 VDD.n153 VSS 0.05fF $ **FLOATING
C1351 VDD.n154 VSS 0.10fF $ **FLOATING
C1352 VDD.t362 VSS 1.28fF
C1353 VDD.t298 VSS 1.58fF
C1354 VDD.t294 VSS 1.09fF
C1355 VDD.n155 VSS 0.79fF $ **FLOATING
C1356 VDD.n156 VSS 0.05fF $ **FLOATING
C1357 VDD.n157 VSS 0.04fF $ **FLOATING
C1358 VDD.n158 VSS 0.10fF $ **FLOATING
C1359 VDD.n159 VSS 0.04fF $ **FLOATING
C1360 VDD.n160 VSS 0.10fF $ **FLOATING
C1361 VDD.n161 VSS 0.05fF $ **FLOATING
C1362 VDD.n162 VSS 0.10fF $ **FLOATING
C1363 VDD.t354 VSS 1.40fF
C1364 VDD.t286 VSS 1.58fF
C1365 VDD.t26 VSS 0.96fF
C1366 VDD.n163 VSS 0.79fF $ **FLOATING
C1367 VDD.n164 VSS 0.06fF $ **FLOATING
C1368 VDD.n165 VSS 0.04fF $ **FLOATING
C1369 VDD.n166 VSS 0.10fF $ **FLOATING
C1370 VDD.n167 VSS 0.04fF $ **FLOATING
C1371 VDD.n168 VSS 0.10fF $ **FLOATING
C1372 VDD.n169 VSS 0.05fF $ **FLOATING
C1373 VDD.n170 VSS 0.10fF $ **FLOATING
C1374 VDD.n171 VSS 0.04fF $ **FLOATING
C1375 VDD.n172 VSS 0.10fF $ **FLOATING
C1376 VDD.t310 VSS 1.53fF
C1377 VDD.t321 VSS 1.58fF
C1378 VDD.t388 VSS 0.84fF
C1379 VDD.n173 VSS 0.79fF $ **FLOATING
C1380 VDD.n174 VSS 0.06fF $ **FLOATING
C1381 VDD.n175 VSS 0.03fF $ **FLOATING
C1382 VDD.n176 VSS 0.10fF $ **FLOATING
C1383 VDD.n177 VSS 0.05fF $ **FLOATING
C1384 VDD.n178 VSS 0.10fF $ **FLOATING
C1385 VDD.n179 VSS 0.05fF $ **FLOATING
C1386 VDD.n180 VSS 0.10fF $ **FLOATING
C1387 VDD.t338 VSS 1.58fF
C1388 VDD.t372 VSS 0.87fF
C1389 VDD.t374 VSS 1.50fF
C1390 VDD.n181 VSS 0.79fF $ **FLOATING
C1391 VDD.n182 VSS 0.05fF $ **FLOATING
C1392 VDD.n183 VSS 0.04fF $ **FLOATING
C1393 VDD.n184 VSS 0.10fF $ **FLOATING
C1394 VDD.n185 VSS 0.05fF $ **FLOATING
C1395 VDD.n186 VSS 0.10fF $ **FLOATING
C1396 VDD.n187 VSS 0.05fF $ **FLOATING
C1397 VDD.n188 VSS 0.10fF $ **FLOATING
C1398 VDD.t307 VSS 1.58fF
C1399 VDD.t128 VSS 1.00fF
C1400 VDD.t315 VSS 1.37fF
C1401 VDD.n189 VSS 0.79fF $ **FLOATING
C1402 VDD.n190 VSS 0.05fF $ **FLOATING
C1403 VDD.n191 VSS 0.04fF $ **FLOATING
C1404 VDD.n192 VSS 0.10fF $ **FLOATING
C1405 VDD.n193 VSS 0.04fF $ **FLOATING
C1406 VDD.n194 VSS 0.10fF $ **FLOATING
C1407 VDD.n195 VSS 0.05fF $ **FLOATING
C1408 VDD.n196 VSS 0.10fF $ **FLOATING
C1409 VDD.t256 VSS 1.13fF
C1410 VDD.t260 VSS 1.24fF
C1411 VDD.n197 VSS 0.79fF $ **FLOATING
C1412 VDD.n198 VSS 0.06fF $ **FLOATING
C1413 VDD.n199 VSS 0.04fF $ **FLOATING
C1414 VDD.n200 VSS 0.10fF $ **FLOATING
C1415 VDD.n201 VSS 0.04fF $ **FLOATING
C1416 VDD.n202 VSS 0.10fF $ **FLOATING
C1417 VDD.n203 VSS 0.05fF $ **FLOATING
C1418 VDD.n204 VSS 0.10fF $ **FLOATING
C1419 VDD.n205 VSS 0.04fF $ **FLOATING
C1420 VDD.n206 VSS 0.10fF $ **FLOATING
C1421 VDD.t330 VSS 1.25fF
C1422 VDD.t336 VSS 1.58fF
C1423 VDD.t244 VSS 1.11fF
C1424 VDD.n207 VSS 0.79fF $ **FLOATING
C1425 VDD.n208 VSS 0.06fF $ **FLOATING
C1426 VDD.n209 VSS 0.03fF $ **FLOATING
C1427 VDD.n210 VSS 0.10fF $ **FLOATING
C1428 VDD.n211 VSS 0.05fF $ **FLOATING
C1429 VDD.n212 VSS 0.10fF $ **FLOATING
C1430 VDD.n213 VSS 0.05fF $ **FLOATING
C1431 VDD.n214 VSS 0.10fF $ **FLOATING
C1432 VDD.t358 VSS 1.38fF
C1433 VDD.t290 VSS 1.58fF
C1434 VDD.t392 VSS 0.99fF
C1435 VDD.n215 VSS 0.79fF $ **FLOATING
C1436 VDD.n216 VSS 0.05fF $ **FLOATING
C1437 VDD.n217 VSS 0.04fF $ **FLOATING
C1438 VDD.n218 VSS 0.10fF $ **FLOATING
C1439 VDD.n219 VSS 0.05fF $ **FLOATING
C1440 VDD.n220 VSS 0.10fF $ **FLOATING
C1441 VDD.n221 VSS 0.05fF $ **FLOATING
C1442 VDD.n222 VSS 0.10fF $ **FLOATING
C1443 VDD.t344 VSS 1.51fF
C1444 VDD.t280 VSS 1.58fF
C1445 VDD.t352 VSS 0.86fF
C1446 VDD.n223 VSS 0.79fF $ **FLOATING
C1447 VDD.n224 VSS 0.05fF $ **FLOATING
C1448 VDD.n225 VSS 0.04fF $ **FLOATING
C1449 VDD.n226 VSS 0.10fF $ **FLOATING
C1450 VDD.n227 VSS 0.04fF $ **FLOATING
C1451 VDD.n228 VSS 0.10fF $ **FLOATING
C1452 VDD.n229 VSS 0.05fF $ **FLOATING
C1453 VDD.n230 VSS 0.10fF $ **FLOATING
C1454 VDD.t408 VSS 1.58fF
C1455 VDD.t410 VSS 0.85fF
C1456 VDD.t414 VSS 1.52fF
C1457 VDD.n231 VSS 0.79fF $ **FLOATING
C1458 VDD.n232 VSS 0.06fF $ **FLOATING
C1459 VDD.n233 VSS 0.04fF $ **FLOATING
C1460 VDD.n234 VSS 0.10fF $ **FLOATING
C1461 VDD.n235 VSS 0.04fF $ **FLOATING
C1462 VDD.n236 VSS 0.10fF $ **FLOATING
C1463 VDD.n237 VSS 0.05fF $ **FLOATING
C1464 VDD.n238 VSS 0.10fF $ **FLOATING
C1465 VDD.n239 VSS 0.04fF $ **FLOATING
C1466 VDD.n240 VSS 0.10fF $ **FLOATING
C1467 VDD.t432 VSS 1.58fF
C1468 VDD.t370 VSS 0.97fF
C1469 VDD.t406 VSS 1.39fF
C1470 VDD.n241 VSS 0.79fF $ **FLOATING
C1471 VDD.n242 VSS 0.06fF $ **FLOATING
C1472 VDD.n243 VSS 0.03fF $ **FLOATING
C1473 VDD.n244 VSS 0.10fF $ **FLOATING
C1474 VDD.n245 VSS 0.05fF $ **FLOATING
C1475 VDD.n246 VSS 0.10fF $ **FLOATING
C1476 VDD.n247 VSS 0.05fF $ **FLOATING
C1477 VDD.n248 VSS 0.11fF $ **FLOATING
C1478 VDD.t366 VSS 1.80fF
C1479 VDD.t250 VSS 1.58fF
C1480 VDD.t300 VSS 1.58fF
C1481 VDD.t424 VSS 1.10fF
C1482 VDD.t428 VSS 1.27fF
C1483 VDD.n249 VSS 0.79fF $ **FLOATING
C1484 VDD.n250 VSS 0.07fF $ **FLOATING
C1485 VDD.n251 VSS 0.68fF $ **FLOATING
C1486 VDD.n252 VSS 0.53fF $ **FLOATING
C1487 VDD.n253 VSS 0.05fF $ **FLOATING
C1488 VDD.n254 VSS 0.00fF $ **FLOATING
C1489 VDD.n255 VSS 0.05fF $ **FLOATING
C1490 VDD.n256 VSS 0.01fF $ **FLOATING
C1491 VDD.n257 VSS 0.06fF $ **FLOATING
C1492 VDD.n258 VSS 0.00fF $ **FLOATING
C1493 VDD.n259 VSS 0.05fF $ **FLOATING
C1494 VDD.n260 VSS 0.01fF $ **FLOATING
C1495 VDD.n261 VSS 0.06fF $ **FLOATING
C1496 VDD.n262 VSS 0.00fF $ **FLOATING
C1497 VDD.n263 VSS 0.05fF $ **FLOATING
C1498 VDD.n264 VSS 0.01fF $ **FLOATING
C1499 VDD.n265 VSS 0.06fF $ **FLOATING
C1500 VDD.n266 VSS 0.00fF $ **FLOATING
C1501 VDD.n267 VSS 0.05fF $ **FLOATING
C1502 VDD.n268 VSS 0.01fF $ **FLOATING
C1503 VDD.n269 VSS 0.05fF $ **FLOATING
C1504 VDD.n270 VSS 0.01fF $ **FLOATING
C1505 VDD.n271 VSS 0.03fF $ **FLOATING
C1506 VDD.n272 VSS 0.01fF $ **FLOATING
C1507 VDD.n273 VSS 0.03fF $ **FLOATING
C1508 VDD.n274 VSS 0.00fF $ **FLOATING
C1509 VDD.n275 VSS 0.34fF $ **FLOATING
C1510 VDD.n276 VSS 0.03fF $ **FLOATING
C1511 VDD.n277 VSS 0.03fF $ **FLOATING
C1512 VDD.t445 VSS 0.04fF
C1513 VDD.t493 VSS 0.04fF
C1514 VDD.n279 VSS 0.20fF $ **FLOATING
C1515 VDD.t487 VSS 0.04fF
C1516 VDD.t3 VSS 0.04fF
C1517 VDD.n280 VSS 0.29fF $ **FLOATING
C1518 sky130_asc_pfet_01v8_lvt_6_1/SOURCE VSS 0.02fF $ **FLOATING
C1519 VDD.n281 VSS 0.06fF $ **FLOATING
C1520 VDD.t5 VSS 0.04fF
C1521 VDD.t1 VSS 0.04fF
C1522 VDD.n282 VSS 0.37fF $ **FLOATING
C1523 VDD.n283 VSS 0.09fF $ **FLOATING
C1524 VDD.n284 VSS 0.07fF $ **FLOATING
C1525 VDD.t122 VSS 1.80fF
C1526 VDD.t274 VSS 1.58fF
C1527 VDD.t168 VSS 1.58fF
C1528 VDD.t172 VSS 1.10fF
C1529 VDD.t227 VSS 1.27fF
C1530 VDD.n285 VSS 0.79fF $ **FLOATING
C1531 VDD.n286 VSS 0.07fF $ **FLOATING
C1532 VDD.t47 VSS 0.04fF
C1533 VDD.t115 VSS 0.04fF
C1534 VDD.n287 VSS 0.29fF $ **FLOATING
C1535 VDD.t241 VSS 0.04fF
C1536 VDD.t201 VSS 0.04fF
C1537 VDD.n288 VSS 0.29fF $ **FLOATING
C1538 VDD.t395 VSS 0.04fF
C1539 VDD.t189 VSS 0.04fF
C1540 VDD.n289 VSS 0.29fF $ **FLOATING
C1541 VDD.t65 VSS 0.04fF
C1542 VDD.t69 VSS 0.04fF
C1543 VDD.n290 VSS 0.29fF $ **FLOATING
C1544 VDD.t39 VSS 0.04fF
C1545 VDD.t55 VSS 0.04fF
C1546 VDD.n291 VSS 0.29fF $ **FLOATING
C1547 VDD.t175 VSS 0.04fF
C1548 VDD.t179 VSS 0.04fF
C1549 VDD.n292 VSS 0.29fF $ **FLOATING
C1550 VDD.t82 VSS 0.04fF
C1551 VDD.t95 VSS 0.04fF
C1552 VDD.n293 VSS 0.29fF $ **FLOATING
C1553 VDD.t208 VSS 0.04fF
C1554 VDD.t76 VSS 0.04fF
C1555 VDD.n294 VSS 0.29fF $ **FLOATING
C1556 VDD.t133 VSS 0.04fF
C1557 VDD.t216 VSS 0.04fF
C1558 VDD.n295 VSS 0.29fF $ **FLOATING
C1559 VDD.t111 VSS 0.04fF
C1560 VDD.t191 VSS 0.04fF
C1561 VDD.n296 VSS 0.29fF $ **FLOATING
C1562 VDD.t249 VSS 0.04fF
C1563 VDD.t297 VSS 0.04fF
C1564 VDD.n297 VSS 0.29fF $ **FLOATING
C1565 VDD.t45 VSS 0.04fF
C1566 VDD.t361 VSS 0.04fF
C1567 VDD.n298 VSS 0.29fF $ **FLOATING
C1568 VDD.t318 VSS 0.04fF
C1569 VDD.t233 VSS 0.04fF
C1570 VDD.n299 VSS 0.29fF $ **FLOATING
C1571 VDD.t239 VSS 0.04fF
C1572 VDD.t283 VSS 0.04fF
C1573 VDD.n300 VSS 0.29fF $ **FLOATING
C1574 VDD.t228 VSS 0.04fF
C1575 VDD.t31 VSS 0.04fF
C1576 VDD.n301 VSS 0.29fF $ **FLOATING
C1577 VDD.t169 VSS 0.04fF
C1578 VDD.t173 VSS 0.04fF
C1579 VDD.n302 VSS 0.29fF $ **FLOATING
C1580 VDD.t123 VSS 0.04fF
C1581 VDD.t275 VSS 0.04fF
C1582 VDD.n303 VSS 0.29fF $ **FLOATING
C1583 sky130_asc_pfet_01v8_lvt_60_2/SOURCE VSS 0.02fF $ **FLOATING
C1584 VDD.n304 VSS 0.06fF $ **FLOATING
C1585 VDD.n305 VSS 0.08fF $ **FLOATING
C1586 VDD.n306 VSS 0.08fF $ **FLOATING
C1587 VDD.n307 VSS 0.08fF $ **FLOATING
C1588 VDD.n308 VSS 0.08fF $ **FLOATING
C1589 VDD.n309 VSS 0.08fF $ **FLOATING
C1590 VDD.n310 VSS 0.08fF $ **FLOATING
C1591 VDD.n311 VSS 0.08fF $ **FLOATING
C1592 VDD.n312 VSS 0.08fF $ **FLOATING
C1593 VDD.n313 VSS 0.08fF $ **FLOATING
C1594 VDD.n314 VSS 0.08fF $ **FLOATING
C1595 VDD.n315 VSS 0.08fF $ **FLOATING
C1596 VDD.n316 VSS 0.08fF $ **FLOATING
C1597 VDD.n317 VSS 0.08fF $ **FLOATING
C1598 VDD.n318 VSS 0.08fF $ **FLOATING
C1599 VDD.n319 VSS 0.08fF $ **FLOATING
C1600 VDD.n320 VSS 0.08fF $ **FLOATING
C1601 VDD.t164 VSS 0.04fF
C1602 VDD.t226 VSS 0.04fF
C1603 VDD.n321 VSS 0.29fF $ **FLOATING
C1604 VDD.t439 VSS 0.04fF
C1605 VDD.t90 VSS 0.04fF
C1606 VDD.n322 VSS 0.29fF $ **FLOATING
C1607 VDD.t377 VSS 0.04fF
C1608 VDD.t102 VSS 0.04fF
C1609 VDD.n323 VSS 0.29fF $ **FLOATING
C1610 VDD.t104 VSS 0.04fF
C1611 VDD.t397 VSS 0.04fF
C1612 VDD.n324 VSS 0.29fF $ **FLOATING
C1613 VDD.t419 VSS 0.04fF
C1614 VDD.t351 VSS 0.04fF
C1615 VDD.n325 VSS 0.29fF $ **FLOATING
C1616 VDD.t43 VSS 0.04fF
C1617 VDD.t365 VSS 0.04fF
C1618 VDD.n326 VSS 0.29fF $ **FLOATING
C1619 VDD.t399 VSS 0.04fF
C1620 VDD.t401 VSS 0.04fF
C1621 VDD.n327 VSS 0.29fF $ **FLOATING
C1622 VDD.t333 VSS 0.04fF
C1623 VDD.t71 VSS 0.04fF
C1624 VDD.n328 VSS 0.29fF $ **FLOATING
C1625 VDD.t403 VSS 0.04fF
C1626 VDD.t405 VSS 0.04fF
C1627 VDD.n329 VSS 0.29fF $ **FLOATING
C1628 VDD.t427 VSS 0.04fF
C1629 VDD.t49 VSS 0.04fF
C1630 VDD.n330 VSS 0.29fF $ **FLOATING
C1631 VDD.t7 VSS 0.04fF
C1632 VDD.t379 VSS 0.04fF
C1633 VDD.n331 VSS 0.29fF $ **FLOATING
C1634 VDD.t381 VSS 0.04fF
C1635 VDD.t314 VSS 0.04fF
C1636 VDD.n332 VSS 0.37fF $ **FLOATING
C1637 VDD.n333 VSS 0.09fF $ **FLOATING
C1638 VDD.n334 VSS 0.08fF $ **FLOATING
C1639 VDD.n335 VSS 0.08fF $ **FLOATING
C1640 VDD.n336 VSS 0.08fF $ **FLOATING
C1641 VDD.n337 VSS 0.08fF $ **FLOATING
C1642 VDD.n338 VSS 0.08fF $ **FLOATING
C1643 VDD.n339 VSS 0.08fF $ **FLOATING
C1644 VDD.n340 VSS 0.08fF $ **FLOATING
C1645 VDD.n341 VSS 0.08fF $ **FLOATING
C1646 VDD.n342 VSS 0.08fF $ **FLOATING
C1647 VDD.n343 VSS 0.08fF $ **FLOATING
C1648 VDD.n344 VSS 0.08fF $ **FLOATING
C1649 VDD.t121 VSS 0.04fF
C1650 VDD.t204 VSS 0.04fF
C1651 VDD.n345 VSS 0.20fF $ **FLOATING
C1652 VDD.n346 VSS 0.06fF $ **FLOATING
C1653 VDD.n347 VSS 0.05fF $ **FLOATING
C1654 VDD.n348 VSS 0.10fF $ **FLOATING
C1655 VDD.t6 VSS 1.58fF
C1656 VDD.t378 VSS 1.05fF
C1657 VDD.t313 VSS 2.01fF
C1658 VDD.t380 VSS 1.32fF
C1659 VDD.n349 VSS 0.79fF $ **FLOATING
C1660 VDD.n350 VSS 0.05fF $ **FLOATING
C1661 VDD.n351 VSS 0.04fF $ **FLOATING
C1662 VDD.n352 VSS 0.10fF $ **FLOATING
C1663 VDD.n353 VSS 0.04fF $ **FLOATING
C1664 VDD.n354 VSS 0.10fF $ **FLOATING
C1665 VDD.n355 VSS 0.05fF $ **FLOATING
C1666 VDD.n356 VSS 0.10fF $ **FLOATING
C1667 VDD.t426 VSS 1.17fF
C1668 VDD.t48 VSS 1.19fF
C1669 VDD.n357 VSS 0.79fF $ **FLOATING
C1670 VDD.n358 VSS 0.06fF $ **FLOATING
C1671 VDD.n359 VSS 0.04fF $ **FLOATING
C1672 VDD.n360 VSS 0.10fF $ **FLOATING
C1673 VDD.n361 VSS 0.04fF $ **FLOATING
C1674 VDD.n362 VSS 0.10fF $ **FLOATING
C1675 VDD.n363 VSS 0.05fF $ **FLOATING
C1676 VDD.n364 VSS 0.10fF $ **FLOATING
C1677 VDD.n365 VSS 0.04fF $ **FLOATING
C1678 VDD.n366 VSS 0.10fF $ **FLOATING
C1679 VDD.t70 VSS 1.30fF
C1680 VDD.t404 VSS 1.58fF
C1681 VDD.t402 VSS 1.07fF
C1682 VDD.n367 VSS 0.79fF $ **FLOATING
C1683 VDD.n368 VSS 0.06fF $ **FLOATING
C1684 VDD.n369 VSS 0.03fF $ **FLOATING
C1685 VDD.n370 VSS 0.10fF $ **FLOATING
C1686 VDD.n371 VSS 0.05fF $ **FLOATING
C1687 VDD.n372 VSS 0.10fF $ **FLOATING
C1688 VDD.n373 VSS 0.05fF $ **FLOATING
C1689 VDD.n374 VSS 0.10fF $ **FLOATING
C1690 VDD.t398 VSS 1.43fF
C1691 VDD.t332 VSS 1.58fF
C1692 VDD.t400 VSS 0.94fF
C1693 VDD.n375 VSS 0.79fF $ **FLOATING
C1694 VDD.n376 VSS 0.05fF $ **FLOATING
C1695 VDD.n377 VSS 0.04fF $ **FLOATING
C1696 VDD.n378 VSS 0.10fF $ **FLOATING
C1697 VDD.n379 VSS 0.05fF $ **FLOATING
C1698 VDD.n380 VSS 0.10fF $ **FLOATING
C1699 VDD.n381 VSS 0.05fF $ **FLOATING
C1700 VDD.n382 VSS 0.10fF $ **FLOATING
C1701 VDD.t350 VSS 1.56fF
C1702 VDD.t364 VSS 1.58fF
C1703 VDD.t42 VSS 0.81fF
C1704 VDD.n383 VSS 0.79fF $ **FLOATING
C1705 VDD.n384 VSS 0.05fF $ **FLOATING
C1706 VDD.n385 VSS 0.04fF $ **FLOATING
C1707 VDD.n386 VSS 0.10fF $ **FLOATING
C1708 VDD.n387 VSS 0.04fF $ **FLOATING
C1709 VDD.n388 VSS 0.10fF $ **FLOATING
C1710 VDD.n389 VSS 0.05fF $ **FLOATING
C1711 VDD.n390 VSS 0.10fF $ **FLOATING
C1712 VDD.t103 VSS 1.58fF
C1713 VDD.t396 VSS 0.89fF
C1714 VDD.t418 VSS 1.47fF
C1715 VDD.n391 VSS 0.79fF $ **FLOATING
C1716 VDD.n392 VSS 0.06fF $ **FLOATING
C1717 VDD.n393 VSS 0.04fF $ **FLOATING
C1718 VDD.n394 VSS 0.10fF $ **FLOATING
C1719 VDD.n395 VSS 0.04fF $ **FLOATING
C1720 VDD.n396 VSS 0.10fF $ **FLOATING
C1721 VDD.n397 VSS 0.05fF $ **FLOATING
C1722 VDD.n398 VSS 0.10fF $ **FLOATING
C1723 VDD.n399 VSS 0.04fF $ **FLOATING
C1724 VDD.n400 VSS 0.10fF $ **FLOATING
C1725 VDD.t89 VSS 1.58fF
C1726 VDD.t376 VSS 1.02fF
C1727 VDD.t101 VSS 1.35fF
C1728 VDD.n401 VSS 0.79fF $ **FLOATING
C1729 VDD.n402 VSS 0.06fF $ **FLOATING
C1730 VDD.n403 VSS 0.03fF $ **FLOATING
C1731 VDD.n404 VSS 0.10fF $ **FLOATING
C1732 VDD.n405 VSS 0.05fF $ **FLOATING
C1733 VDD.n406 VSS 0.10fF $ **FLOATING
C1734 VDD.n407 VSS 0.05fF $ **FLOATING
C1735 VDD.n408 VSS 0.10fF $ **FLOATING
C1736 VDD.t225 VSS 1.15fF
C1737 VDD.t438 VSS 1.22fF
C1738 VDD.n409 VSS 0.79fF $ **FLOATING
C1739 VDD.n410 VSS 0.05fF $ **FLOATING
C1740 VDD.n411 VSS 0.04fF $ **FLOATING
C1741 VDD.n412 VSS 0.10fF $ **FLOATING
C1742 VDD.n413 VSS 0.05fF $ **FLOATING
C1743 VDD.n414 VSS 0.10fF $ **FLOATING
C1744 VDD.n415 VSS 0.05fF $ **FLOATING
C1745 VDD.n416 VSS 0.10fF $ **FLOATING
C1746 VDD.t120 VSS 1.28fF
C1747 VDD.t163 VSS 1.58fF
C1748 VDD.t203 VSS 1.09fF
C1749 VDD.n417 VSS 0.79fF $ **FLOATING
C1750 VDD.n418 VSS 0.05fF $ **FLOATING
C1751 VDD.n419 VSS 0.04fF $ **FLOATING
C1752 VDD.n420 VSS 0.06fF $ **FLOATING
C1753 VDD.n421 VSS 0.09fF $ **FLOATING
C1754 VDD.n422 VSS 0.04fF $ **FLOATING
C1755 VDD.n423 VSS 0.09fF $ **FLOATING
C1756 VDD.n424 VSS 0.05fF $ **FLOATING
C1757 VDD.n425 VSS 0.10fF $ **FLOATING
C1758 VDD.t200 VSS 1.40fF
C1759 VDD.t114 VSS 1.58fF
C1760 VDD.t46 VSS 0.96fF
C1761 VDD.n426 VSS 0.79fF $ **FLOATING
C1762 VDD.n427 VSS 0.06fF $ **FLOATING
C1763 VDD.n428 VSS 0.04fF $ **FLOATING
C1764 VDD.n429 VSS 0.10fF $ **FLOATING
C1765 VDD.n430 VSS 0.04fF $ **FLOATING
C1766 VDD.n431 VSS 0.10fF $ **FLOATING
C1767 VDD.n432 VSS 0.05fF $ **FLOATING
C1768 VDD.n433 VSS 0.10fF $ **FLOATING
C1769 VDD.n434 VSS 0.04fF $ **FLOATING
C1770 VDD.n435 VSS 0.10fF $ **FLOATING
C1771 VDD.t394 VSS 1.53fF
C1772 VDD.t240 VSS 1.58fF
C1773 VDD.t188 VSS 0.84fF
C1774 VDD.n436 VSS 0.79fF $ **FLOATING
C1775 VDD.n437 VSS 0.06fF $ **FLOATING
C1776 VDD.n438 VSS 0.03fF $ **FLOATING
C1777 VDD.n439 VSS 0.10fF $ **FLOATING
C1778 VDD.n440 VSS 0.05fF $ **FLOATING
C1779 VDD.n441 VSS 0.10fF $ **FLOATING
C1780 VDD.n442 VSS 0.05fF $ **FLOATING
C1781 VDD.n443 VSS 0.10fF $ **FLOATING
C1782 VDD.t54 VSS 1.58fF
C1783 VDD.t64 VSS 0.87fF
C1784 VDD.t68 VSS 1.50fF
C1785 VDD.n444 VSS 0.79fF $ **FLOATING
C1786 VDD.n445 VSS 0.05fF $ **FLOATING
C1787 VDD.n446 VSS 0.04fF $ **FLOATING
C1788 VDD.n447 VSS 0.10fF $ **FLOATING
C1789 VDD.n448 VSS 0.05fF $ **FLOATING
C1790 VDD.n449 VSS 0.10fF $ **FLOATING
C1791 VDD.n450 VSS 0.05fF $ **FLOATING
C1792 VDD.n451 VSS 0.10fF $ **FLOATING
C1793 VDD.t174 VSS 1.58fF
C1794 VDD.t178 VSS 1.00fF
C1795 VDD.t38 VSS 1.37fF
C1796 VDD.n452 VSS 0.79fF $ **FLOATING
C1797 VDD.n453 VSS 0.05fF $ **FLOATING
C1798 VDD.n454 VSS 0.04fF $ **FLOATING
C1799 VDD.n455 VSS 0.10fF $ **FLOATING
C1800 VDD.n456 VSS 0.04fF $ **FLOATING
C1801 VDD.n457 VSS 0.10fF $ **FLOATING
C1802 VDD.n458 VSS 0.05fF $ **FLOATING
C1803 VDD.n459 VSS 0.10fF $ **FLOATING
C1804 VDD.t81 VSS 1.13fF
C1805 VDD.t94 VSS 1.24fF
C1806 VDD.n460 VSS 0.79fF $ **FLOATING
C1807 VDD.n461 VSS 0.06fF $ **FLOATING
C1808 VDD.n462 VSS 0.04fF $ **FLOATING
C1809 VDD.n463 VSS 0.10fF $ **FLOATING
C1810 VDD.n464 VSS 0.04fF $ **FLOATING
C1811 VDD.n465 VSS 0.10fF $ **FLOATING
C1812 VDD.n466 VSS 0.05fF $ **FLOATING
C1813 VDD.n467 VSS 0.10fF $ **FLOATING
C1814 VDD.n468 VSS 0.04fF $ **FLOATING
C1815 VDD.n469 VSS 0.10fF $ **FLOATING
C1816 VDD.t215 VSS 1.25fF
C1817 VDD.t75 VSS 1.58fF
C1818 VDD.t207 VSS 1.11fF
C1819 VDD.n470 VSS 0.79fF $ **FLOATING
C1820 VDD.n471 VSS 0.06fF $ **FLOATING
C1821 VDD.n472 VSS 0.03fF $ **FLOATING
C1822 VDD.n473 VSS 0.10fF $ **FLOATING
C1823 VDD.n474 VSS 0.05fF $ **FLOATING
C1824 VDD.n475 VSS 0.10fF $ **FLOATING
C1825 VDD.n476 VSS 0.05fF $ **FLOATING
C1826 VDD.n477 VSS 0.10fF $ **FLOATING
C1827 VDD.t110 VSS 1.38fF
C1828 VDD.t132 VSS 1.58fF
C1829 VDD.t190 VSS 0.99fF
C1830 VDD.n478 VSS 0.79fF $ **FLOATING
C1831 VDD.n479 VSS 0.05fF $ **FLOATING
C1832 VDD.n480 VSS 0.04fF $ **FLOATING
C1833 VDD.n481 VSS 0.10fF $ **FLOATING
C1834 VDD.n482 VSS 0.05fF $ **FLOATING
C1835 VDD.n483 VSS 0.10fF $ **FLOATING
C1836 VDD.n484 VSS 0.05fF $ **FLOATING
C1837 VDD.n485 VSS 0.10fF $ **FLOATING
C1838 VDD.t360 VSS 1.51fF
C1839 VDD.t296 VSS 1.58fF
C1840 VDD.t248 VSS 0.86fF
C1841 VDD.n486 VSS 0.79fF $ **FLOATING
C1842 VDD.n487 VSS 0.05fF $ **FLOATING
C1843 VDD.n488 VSS 0.04fF $ **FLOATING
C1844 VDD.n489 VSS 0.10fF $ **FLOATING
C1845 VDD.n490 VSS 0.04fF $ **FLOATING
C1846 VDD.n491 VSS 0.10fF $ **FLOATING
C1847 VDD.n492 VSS 0.05fF $ **FLOATING
C1848 VDD.n493 VSS 0.10fF $ **FLOATING
C1849 VDD.t317 VSS 1.58fF
C1850 VDD.t232 VSS 0.85fF
C1851 VDD.t44 VSS 1.52fF
C1852 VDD.n494 VSS 0.79fF $ **FLOATING
C1853 VDD.n495 VSS 0.06fF $ **FLOATING
C1854 VDD.n496 VSS 0.04fF $ **FLOATING
C1855 VDD.n497 VSS 0.10fF $ **FLOATING
C1856 VDD.n498 VSS 0.04fF $ **FLOATING
C1857 VDD.n499 VSS 0.10fF $ **FLOATING
C1858 VDD.n500 VSS 0.05fF $ **FLOATING
C1859 VDD.n501 VSS 0.10fF $ **FLOATING
C1860 VDD.n502 VSS 0.04fF $ **FLOATING
C1861 VDD.n503 VSS 0.10fF $ **FLOATING
C1862 VDD.t30 VSS 1.58fF
C1863 VDD.t238 VSS 0.97fF
C1864 VDD.t282 VSS 1.39fF
C1865 VDD.n504 VSS 0.79fF $ **FLOATING
C1866 VDD.n505 VSS 0.06fF $ **FLOATING
C1867 VDD.n506 VSS 0.03fF $ **FLOATING
C1868 VDD.n507 VSS 0.10fF $ **FLOATING
C1869 VDD.n508 VSS 0.05fF $ **FLOATING
C1870 VDD.n509 VSS 0.10fF $ **FLOATING
C1871 VDD.n510 VSS 0.05fF $ **FLOATING
C1872 VDD.n511 VSS 0.11fF $ **FLOATING
C1873 VDD.n512 VSS 0.49fF $ **FLOATING
C1874 sky130_asc_pfet_01v8_lvt_6_1/VPWR VSS 0.03fF $ **FLOATING
C1875 VDD.n513 VSS 0.11fF $ **FLOATING
C1876 VDD.n514 VSS 0.08fF $ **FLOATING
C1877 VDD.n515 VSS 0.43fF $ **FLOATING
C1878 VDD.n516 VSS 0.05fF $ **FLOATING
C1879 VDD.n517 VSS 0.10fF $ **FLOATING
C1880 VDD.t486 VSS 1.80fF
C1881 VDD.t2 VSS 1.58fF
C1882 VDD.t444 VSS 1.58fF
C1883 VDD.t492 VSS 1.05fF
C1884 VDD.t0 VSS 2.01fF
C1885 VDD.t4 VSS 1.32fF
C1886 VDD.n518 VSS 0.79fF $ **FLOATING
C1887 VDD.n519 VSS 0.05fF $ **FLOATING
C1888 VDD.n520 VSS 0.04fF $ **FLOATING
C1889 VDD.n521 VSS 0.09fF $ **FLOATING
C1890 VDD.n522 VSS 0.10fF $ **FLOATING
C1891 VDD.n523 VSS 0.38fF $ **FLOATING
C1892 sky130_asc_res_xhigh_po_2p85_1_20/VPWR VSS 0.82fF $ **FLOATING
C1893 sky130_asc_res_xhigh_po_2p85_1_18/VPWR VSS 1.13fF $ **FLOATING
C1894 VDD.n524 VSS 0.56fF $ **FLOATING
C1895 VDD.n525 VSS 0.05fF $ **FLOATING
C1896 VDD.n526 VSS 0.00fF $ **FLOATING
C1897 VDD.n527 VSS 0.05fF $ **FLOATING
C1898 VDD.n528 VSS 0.01fF $ **FLOATING
C1899 VDD.n529 VSS 0.06fF $ **FLOATING
C1900 VDD.n530 VSS 0.00fF $ **FLOATING
C1901 VDD.n531 VSS 0.05fF $ **FLOATING
C1902 VDD.n532 VSS 0.01fF $ **FLOATING
C1903 VDD.n533 VSS 0.06fF $ **FLOATING
C1904 VDD.n534 VSS 0.00fF $ **FLOATING
C1905 VDD.n535 VSS 0.05fF $ **FLOATING
C1906 VDD.n536 VSS 0.01fF $ **FLOATING
C1907 VDD.n537 VSS 0.06fF $ **FLOATING
C1908 VDD.n538 VSS 0.00fF $ **FLOATING
C1909 VDD.n539 VSS 0.05fF $ **FLOATING
C1910 VDD.n540 VSS 0.01fF $ **FLOATING
C1911 VDD.n541 VSS 0.05fF $ **FLOATING
C1912 VDD.n542 VSS 0.01fF $ **FLOATING
C1913 VDD.n543 VSS 0.03fF $ **FLOATING
C1914 VDD.n544 VSS 0.01fF $ **FLOATING
C1915 VDD.n545 VSS 0.03fF $ **FLOATING
C1916 VDD.n546 VSS 0.00fF $ **FLOATING
C1917 VDD.n547 VSS 0.34fF $ **FLOATING
C1918 VDD.n548 VSS 0.03fF $ **FLOATING
C1919 VDD.n549 VSS 0.03fF $ **FLOATING
C1920 VDD.n551 VSS 0.06fF $ **FLOATING
C1921 VDD.n552 VSS 0.10fF $ **FLOATING
C1922 VDD.n553 VSS 0.06fF $ **FLOATING
C1923 VDD.n554 VSS 0.10fF $ **FLOATING
C1924 VDD.n555 VSS 0.05fF $ **FLOATING
C1925 VDD.n556 VSS 0.07fF $ **FLOATING
C1926 sky130_asc_pfet_01v8_lvt_12_1/VPWR VSS 0.03fF $ **FLOATING
C1927 VDD.t134 VSS 1.80fF
C1928 VDD.t430 VSS 1.58fF
C1929 VDD.t434 VSS 1.58fF
C1930 VDD.t79 VSS 1.30fF
C1931 VDD.n557 VSS 0.79fF $ **FLOATING
C1932 VDD.t34 VSS 1.07fF
C1933 VDD.t96 VSS 1.58fF
C1934 VDD.t386 VSS 1.17fF
C1935 VDD.n558 VSS 0.79fF $ **FLOATING
C1936 VDD.t412 VSS 1.19fF
C1937 VDD.t346 VSS 1.58fF
C1938 VDD.t422 VSS 1.05fF
C1939 VDD.n559 VSS 0.79fF $ **FLOATING
C1940 VDD.t59 VSS 1.32fF
C1941 VDD.t416 VSS 2.01fF
C1942 VDD.n560 VSS 0.11fF $ **FLOATING
C1943 VDD.t347 VSS 0.04fF
C1944 VDD.t423 VSS 0.04fF
C1945 VDD.n561 VSS 0.29fF $ **FLOATING
C1946 VDD.t387 VSS 0.04fF
C1947 VDD.t413 VSS 0.04fF
C1948 VDD.n562 VSS 0.29fF $ **FLOATING
C1949 VDD.t35 VSS 0.04fF
C1950 VDD.t97 VSS 0.04fF
C1951 VDD.n563 VSS 0.29fF $ **FLOATING
C1952 VDD.t435 VSS 0.04fF
C1953 VDD.t80 VSS 0.04fF
C1954 VDD.n564 VSS 0.29fF $ **FLOATING
C1955 VDD.t135 VSS 0.04fF
C1956 VDD.t431 VSS 0.04fF
C1957 VDD.n565 VSS 0.29fF $ **FLOATING
C1958 sky130_asc_pfet_01v8_lvt_12_1/SOURCE VSS 0.02fF $ **FLOATING
C1959 VDD.n566 VSS 0.06fF $ **FLOATING
C1960 VDD.n567 VSS 0.08fF $ **FLOATING
C1961 VDD.n568 VSS 0.08fF $ **FLOATING
C1962 VDD.n569 VSS 0.08fF $ **FLOATING
C1963 VDD.n570 VSS 0.09fF $ **FLOATING
C1964 VDD.t60 VSS 0.04fF
C1965 VDD.t417 VSS 0.04fF
C1966 VDD.n571 VSS 0.19fF $ **FLOATING
C1967 VDD.n572 VSS 0.15fF $ **FLOATING
C1968 VDD.n573 VSS 0.09fF $ **FLOATING
C1969 VDD.n574 VSS 0.53fF $ **FLOATING
C1970 VDD.n575 VSS 0.08fF $ **FLOATING
C1971 VDD.n576 VSS 0.05fF $ **FLOATING
C1972 VDD.n577 VSS 0.04fF $ **FLOATING
C1973 VDD.n578 VSS 0.10fF $ **FLOATING
C1974 VDD.n579 VSS 0.10fF $ **FLOATING
C1975 VDD.n580 VSS 0.04fF $ **FLOATING
C1976 VDD.n581 VSS 0.05fF $ **FLOATING
C1977 VDD.n582 VSS 0.04fF $ **FLOATING
C1978 VDD.n583 VSS 0.10fF $ **FLOATING
C1979 VDD.n584 VSS 0.10fF $ **FLOATING
C1980 VDD.n585 VSS 0.04fF $ **FLOATING
C1981 VDD.n586 VSS 0.05fF $ **FLOATING
C1982 VDD.n587 VSS 0.04fF $ **FLOATING
C1983 VDD.n588 VSS 0.11fF $ **FLOATING
C1984 VDD.n589 VSS 0.44fF $ **FLOATING
C1985 sky130_asc_cap_mim_m3_1_9/VPWR VSS 1.78fF $ **FLOATING
C1986 sky130_asc_nfet_01v8_lvt_9_1/VPWR VSS 2.37fF $ **FLOATING
C1987 sky130_asc_pnp_05v5_W3p40L3p40_8_2/VPWR VSS 3.03fF $ **FLOATING
C1988 sky130_asc_res_xhigh_po_2p85_1_0/VPWR VSS 2.78fF $ **FLOATING
C1989 VDD.n590 VSS 0.60fF $ **FLOATING
C1990 VDD.n591 VSS 0.05fF $ **FLOATING
C1991 VDD.n592 VSS 0.00fF $ **FLOATING
C1992 VDD.n593 VSS 0.05fF $ **FLOATING
C1993 VDD.n594 VSS 0.01fF $ **FLOATING
C1994 VDD.n595 VSS 0.06fF $ **FLOATING
C1995 VDD.n596 VSS 0.00fF $ **FLOATING
C1996 VDD.n597 VSS 0.05fF $ **FLOATING
C1997 VDD.n598 VSS 0.01fF $ **FLOATING
C1998 VDD.n599 VSS 0.06fF $ **FLOATING
C1999 VDD.n600 VSS 0.00fF $ **FLOATING
C2000 VDD.n601 VSS 0.05fF $ **FLOATING
C2001 VDD.n602 VSS 0.01fF $ **FLOATING
C2002 VDD.n603 VSS 0.06fF $ **FLOATING
C2003 VDD.n604 VSS 0.00fF $ **FLOATING
C2004 VDD.n605 VSS 0.05fF $ **FLOATING
C2005 VDD.n606 VSS 0.01fF $ **FLOATING
C2006 VDD.n607 VSS 0.05fF $ **FLOATING
C2007 VDD.n608 VSS 0.01fF $ **FLOATING
C2008 VDD.n609 VSS 0.03fF $ **FLOATING
C2009 VDD.n610 VSS 0.01fF $ **FLOATING
C2010 VDD.n611 VSS 0.03fF $ **FLOATING
C2011 VDD.n612 VSS 0.00fF $ **FLOATING
C2012 VDD.n613 VSS 0.34fF $ **FLOATING
C2013 VDD.n614 VSS 0.03fF $ **FLOATING
C2014 VDD.n615 VSS 0.03fF $ **FLOATING
C2015 VDD.t459 VSS 1.80fF
C2016 VDD.t477 VSS 1.58fF
C2017 VDD.t480 VSS 1.58fF
C2018 VDD.t447 VSS 1.30fF
C2019 VDD.t456 VSS 1.58fF
C2020 VDD.t450 VSS 1.07fF
C2021 VDD.n617 VSS 0.79fF $ **FLOATING
C2022 VDD.n618 VSS 0.06fF $ **FLOATING
C2023 VDD.t463 VSS 0.04fF
C2024 VDD.t466 VSS 0.04fF
C2025 VDD.n619 VSS 0.29fF $ **FLOATING
C2026 VDD.t469 VSS 0.04fF
C2027 VDD.t454 VSS 0.04fF
C2028 VDD.n620 VSS 0.29fF $ **FLOATING
C2029 VDD.t451 VSS 0.04fF
C2030 VDD.t457 VSS 0.04fF
C2031 VDD.n621 VSS 0.29fF $ **FLOATING
C2032 VDD.t481 VSS 0.04fF
C2033 VDD.t448 VSS 0.04fF
C2034 VDD.n622 VSS 0.29fF $ **FLOATING
C2035 VDD.t460 VSS 0.04fF
C2036 VDD.t478 VSS 0.04fF
C2037 VDD.n623 VSS 0.29fF $ **FLOATING
C2038 sky130_asc_pfet_01v8_lvt_12_0/SOURCE VSS 0.02fF $ **FLOATING
C2039 VDD.n624 VSS 0.06fF $ **FLOATING
C2040 VDD.n625 VSS 0.08fF $ **FLOATING
C2041 VDD.n626 VSS 0.08fF $ **FLOATING
C2042 VDD.n627 VSS 0.08fF $ **FLOATING
C2043 VDD.n628 VSS 0.08fF $ **FLOATING
C2044 VDD.t472 VSS 0.04fF
C2045 VDD.t475 VSS 0.04fF
C2046 VDD.n629 VSS 0.32fF $ **FLOATING
C2047 VDD.n630 VSS 0.06fF $ **FLOATING
C2048 sky130_asc_pfet_01v8_lvt_12_0/GATE VSS 0.02fF $ **FLOATING
C2049 VDD.t458 VSS 0.95fF
C2050 VDD.n631 VSS 0.26fF $ **FLOATING
C2051 VDD.n632 VSS 0.04fF $ **FLOATING
C2052 VDD.n633 VSS 0.04fF $ **FLOATING
C2053 VDD.n634 VSS 0.05fF $ **FLOATING
C2054 VDD.t476 VSS 0.95fF
C2055 VDD.n635 VSS 0.22fF $ **FLOATING
C2056 VDD.n636 VSS 0.04fF $ **FLOATING
C2057 VDD.n637 VSS 0.05fF $ **FLOATING
C2058 VDD.t479 VSS 0.95fF
C2059 VDD.n638 VSS 0.22fF $ **FLOATING
C2060 VDD.n639 VSS 0.04fF $ **FLOATING
C2061 VDD.n640 VSS 0.05fF $ **FLOATING
C2062 VDD.t446 VSS 0.95fF
C2063 VDD.n641 VSS 0.22fF $ **FLOATING
C2064 VDD.n642 VSS 0.04fF $ **FLOATING
C2065 VDD.n643 VSS 0.05fF $ **FLOATING
C2066 VDD.t449 VSS 0.95fF
C2067 VDD.n644 VSS 0.22fF $ **FLOATING
C2068 VDD.n645 VSS 0.04fF $ **FLOATING
C2069 VDD.n646 VSS 0.05fF $ **FLOATING
C2070 VDD.t455 VSS 0.95fF
C2071 VDD.n647 VSS 0.25fF $ **FLOATING
C2072 VDD.n648 VSS 0.05fF $ **FLOATING
C2073 VDD.t467 VSS 0.95fF
C2074 VDD.n649 VSS 0.26fF $ **FLOATING
C2075 VDD.n650 VSS 0.05fF $ **FLOATING
C2076 VDD.t452 VSS 0.95fF
C2077 VDD.n651 VSS 0.22fF $ **FLOATING
C2078 VDD.n652 VSS 0.04fF $ **FLOATING
C2079 VDD.n653 VSS 0.05fF $ **FLOATING
C2080 VDD.n654 VSS 0.04fF $ **FLOATING
C2081 VDD.n655 VSS 0.05fF $ **FLOATING
C2082 VDD.t461 VSS 0.95fF
C2083 VDD.n656 VSS 0.22fF $ **FLOATING
C2084 VDD.n657 VSS 0.04fF $ **FLOATING
C2085 VDD.n658 VSS 0.05fF $ **FLOATING
C2086 VDD.t464 VSS 0.95fF
C2087 VDD.n659 VSS 0.22fF $ **FLOATING
C2088 VDD.n660 VSS 0.04fF $ **FLOATING
C2089 VDD.n661 VSS 0.05fF $ **FLOATING
C2090 VDD.t470 VSS 0.95fF
C2091 VDD.n662 VSS 0.23fF $ **FLOATING
C2092 VDD.t473 VSS 1.03fF
C2093 VDD.n663 VSS 0.25fF $ **FLOATING
C2094 VDD.n664 VSS 0.11fF $ **FLOATING
C2095 VDD.n665 VSS 0.07fF $ **FLOATING
C2096 VDD.n666 VSS 0.05fF $ **FLOATING
C2097 VDD.n667 VSS 0.06fF $ **FLOATING
C2098 VDD.n668 VSS 0.05fF $ **FLOATING
C2099 VDD.t462 VSS 1.58fF
C2100 VDD.t465 VSS 1.05fF
C2101 VDD.t474 VSS 2.01fF
C2102 VDD.t471 VSS 1.32fF
C2103 VDD.n669 VSS 0.79fF $ **FLOATING
C2104 VDD.n670 VSS 0.05fF $ **FLOATING
C2105 VDD.n671 VSS 0.04fF $ **FLOATING
C2106 VDD.n672 VSS 0.09fF $ **FLOATING
C2107 VDD.n673 VSS 0.04fF $ **FLOATING
C2108 VDD.n674 VSS 0.10fF $ **FLOATING
C2109 VDD.n675 VSS 0.05fF $ **FLOATING
C2110 VDD.n676 VSS 0.10fF $ **FLOATING
C2111 VDD.t468 VSS 1.17fF
C2112 VDD.t453 VSS 1.19fF
C2113 VDD.n677 VSS 0.79fF $ **FLOATING
C2114 VDD.n678 VSS 0.06fF $ **FLOATING
C2115 VDD.n679 VSS 0.04fF $ **FLOATING
C2116 VDD.n680 VSS 0.10fF $ **FLOATING
C2117 VDD.n681 VSS 0.04fF $ **FLOATING
C2118 VDD.n682 VSS 0.10fF $ **FLOATING
C2119 VDD.n683 VSS 0.05fF $ **FLOATING
C2120 VDD.n684 VSS 0.10fF $ **FLOATING
C2121 VDD.n685 VSS 0.04fF $ **FLOATING
C2122 VDD.n686 VSS 0.11fF $ **FLOATING
C2123 VDD.n687 VSS 0.44fF $ **FLOATING
C2124 sky130_asc_cap_mim_m3_1_5/VPWR VSS 1.76fF $ **FLOATING
C2125 sky130_asc_pnp_05v5_W3p40L3p40_1_0/VPWR VSS 1.72fF $ **FLOATING
C2126 sky130_asc_nfet_01v8_lvt_9_2/VPWR VSS 1.30fF $ **FLOATING
C2127 sky130_asc_pnp_05v5_W3p40L3p40_8_1/VPWR VSS 3.03fF $ **FLOATING
C2128 sky130_asc_res_xhigh_po_2p85_1_8/VPWR VSS 2.78fF $ **FLOATING
C2129 VDD.n688 VSS 0.60fF $ **FLOATING
C2130 VDD.n689 VSS 0.05fF $ **FLOATING
C2131 VDD.n690 VSS 0.00fF $ **FLOATING
C2132 VDD.n691 VSS 0.05fF $ **FLOATING
C2133 VDD.n692 VSS 0.01fF $ **FLOATING
C2134 VDD.n693 VSS 0.06fF $ **FLOATING
C2135 VDD.n694 VSS 0.00fF $ **FLOATING
C2136 VDD.n695 VSS 0.05fF $ **FLOATING
C2137 VDD.n696 VSS 0.01fF $ **FLOATING
C2138 VDD.n697 VSS 0.06fF $ **FLOATING
C2139 VDD.n698 VSS 0.00fF $ **FLOATING
C2140 VDD.n699 VSS 0.05fF $ **FLOATING
C2141 VDD.n700 VSS 0.01fF $ **FLOATING
C2142 VDD.n701 VSS 0.06fF $ **FLOATING
C2143 VDD.n702 VSS 0.00fF $ **FLOATING
C2144 VDD.n703 VSS 0.05fF $ **FLOATING
C2145 VDD.n704 VSS 0.01fF $ **FLOATING
C2146 VDD.n705 VSS 0.05fF $ **FLOATING
C2147 VDD.n706 VSS 0.01fF $ **FLOATING
C2148 VDD.n707 VSS 0.03fF $ **FLOATING
C2149 VDD.n708 VSS 0.01fF $ **FLOATING
C2150 VDD.n709 VSS 0.03fF $ **FLOATING
C2151 VDD.n710 VSS 0.00fF $ **FLOATING
C2152 VDD.n711 VSS 0.34fF $ **FLOATING
C2153 VDD.n712 VSS 0.03fF $ **FLOATING
C2154 VDD.n713 VSS 0.03fF $ **FLOATING
C2155 VDD.n715 VSS 0.05fF $ **FLOATING
C2156 VDD.t491 VSS 0.04fF
C2157 VDD.t489 VSS 0.04fF
C2158 VDD.n716 VSS 0.29fF $ **FLOATING
C2159 sky130_asc_pfet_01v8_lvt_6_0/SOURCE VSS 0.02fF $ **FLOATING
C2160 VDD.n717 VSS 0.03fF $ **FLOATING
C2161 VDD.t485 VSS 0.04fF
C2162 VDD.t483 VSS 0.04fF
C2163 VDD.n718 VSS 0.29fF $ **FLOATING
C2164 VDD.t443 VSS 0.04fF
C2165 VDD.t441 VSS 0.04fF
C2166 VDD.n719 VSS 0.37fF $ **FLOATING
C2167 VDD.n720 VSS 0.09fF $ **FLOATING
C2168 VDD.n721 VSS 0.04fF $ **FLOATING
C2169 VDD.n722 VSS 0.10fF $ **FLOATING
C2170 VDD.t490 VSS 1.80fF
C2171 VDD.t488 VSS 1.58fF
C2172 VDD.t484 VSS 1.58fF
C2173 VDD.t482 VSS 1.05fF
C2174 VDD.n723 VSS 0.79fF $ **FLOATING
C2175 VDD.n724 VSS 0.05fF $ **FLOATING
C2176 sky130_asc_res_xhigh_po_2p85_1_5/VPWR VSS 1.33fF $ **FLOATING
C2177 sky130_asc_res_xhigh_po_2p85_1_6/VPWR VSS 0.99fF $ **FLOATING
C2178 sky130_asc_cap_mim_m3_1_7/VPWR VSS 1.99fF $ **FLOATING
C2179 sky130_asc_pfet_01v8_lvt_6_0/VPWR VSS 0.03fF $ **FLOATING
C2180 VDD.t442 VSS 1.32fF
C2181 VDD.t440 VSS 2.01fF
C2182 VDD.n725 VSS 0.11fF $ **FLOATING
C2183 VDD.n726 VSS 0.08fF $ **FLOATING
C2184 VDD.n727 VSS 1.46fF $ **FLOATING
C2185 VDD.n728 VSS 0.10fF $ **FLOATING
C2186 VDD.n729 VSS 0.10fF $ **FLOATING
C2187 VDD.n730 VSS 0.04fF $ **FLOATING
C2188 VDD.n731 VSS 0.05fF $ **FLOATING
C2189 VDD.n732 VSS 0.04fF $ **FLOATING
C2190 VDD.n733 VSS 0.05fF $ **FLOATING
C2191 VDD.n734 VSS 0.10fF $ **FLOATING
C2192 VDD.n735 VSS 0.05fF $ **FLOATING
C2193 VDD.n736 VSS 0.06fF $ **FLOATING
C2194 VDD.n737 VSS 0.32fF $ **FLOATING
C2195 sky130_asc_pnp_05v5_W3p40L3p40_8_0/VPWR VSS 2.29fF $ **FLOATING
C2196 sky130_asc_res_xhigh_po_2p85_1_17/VPWR VSS 2.82fF $ **FLOATING
C2197 VDD.n738 VSS 0.65fF $ **FLOATING
C2198 VDD.n739 VSS 0.05fF $ **FLOATING
C2199 VDD.n740 VSS 0.00fF $ **FLOATING
C2200 VDD.n741 VSS 0.05fF $ **FLOATING
C2201 VDD.n742 VSS 0.01fF $ **FLOATING
C2202 VDD.n743 VSS 0.06fF $ **FLOATING
C2203 VDD.n744 VSS 0.00fF $ **FLOATING
C2204 VDD.n745 VSS 0.05fF $ **FLOATING
C2205 VDD.n746 VSS 0.01fF $ **FLOATING
C2206 VDD.n747 VSS 0.06fF $ **FLOATING
C2207 VDD.n748 VSS 0.00fF $ **FLOATING
C2208 VDD.n749 VSS 0.05fF $ **FLOATING
C2209 VDD.n750 VSS 0.01fF $ **FLOATING
C2210 VDD.n751 VSS 0.06fF $ **FLOATING
C2211 VDD.n752 VSS 0.00fF $ **FLOATING
C2212 VDD.n753 VSS 0.05fF $ **FLOATING
C2213 VDD.n754 VSS 0.01fF $ **FLOATING
C2214 VDD.n755 VSS 0.05fF $ **FLOATING
C2215 VDD.n756 VSS 0.01fF $ **FLOATING
C2216 VDD.n757 VSS 0.03fF $ **FLOATING
C2217 VDD.n758 VSS 0.01fF $ **FLOATING
C2218 VDD.n759 VSS 0.03fF $ **FLOATING
C2219 VDD.n760 VSS 0.00fF $ **FLOATING
C2220 VDD.n761 VSS 0.34fF $ **FLOATING
C2221 VDD.n762 VSS 0.03fF $ **FLOATING
C2222 VDD.n763 VSS 0.03fF $ **FLOATING
C2223 sky130_asc_res_xhigh_po_2p85_1_2/VPWR VSS 1.00fF $ **FLOATING
C2224 sky130_asc_res_xhigh_po_2p85_1_9/VPWR VSS 0.99fF $ **FLOATING
C2225 sky130_asc_cap_mim_m3_1_6/VPWR VSS 1.88fF $ **FLOATING
C2226 sky130_asc_res_xhigh_po_2p85_1_22/VPWR VSS 2.18fF $ **FLOATING
C2227 sky130_asc_pnp_05v5_W3p40L3p40_8_3/VPWR VSS 2.74fF $ **FLOATING
C2228 sky130_asc_res_xhigh_po_2p85_1_16/VPWR VSS 2.82fF $ **FLOATING
C2229 VDD.n765 VSS 0.65fF $ **FLOATING
C2230 VDD.n766 VSS 0.05fF $ **FLOATING
C2231 VDD.n767 VSS 0.00fF $ **FLOATING
C2232 VDD.n768 VSS 0.05fF $ **FLOATING
C2233 VDD.n769 VSS 0.01fF $ **FLOATING
C2234 VDD.n770 VSS 0.06fF $ **FLOATING
C2235 VDD.n771 VSS 0.00fF $ **FLOATING
C2236 VDD.n772 VSS 0.05fF $ **FLOATING
C2237 VDD.n773 VSS 0.01fF $ **FLOATING
C2238 VDD.n774 VSS 0.06fF $ **FLOATING
C2239 VDD.n775 VSS 0.00fF $ **FLOATING
C2240 VDD.n776 VSS 0.05fF $ **FLOATING
C2241 VDD.n777 VSS 0.01fF $ **FLOATING
C2242 VDD.n778 VSS 0.06fF $ **FLOATING
C2243 VDD.n779 VSS 0.00fF $ **FLOATING
C2244 VDD.n780 VSS 0.05fF $ **FLOATING
C2245 VDD.n781 VSS 0.01fF $ **FLOATING
C2246 VDD.n782 VSS 0.05fF $ **FLOATING
C2247 VDD.n783 VSS 0.01fF $ **FLOATING
C2248 VDD.n784 VSS 0.03fF $ **FLOATING
C2249 VDD.n785 VSS 0.01fF $ **FLOATING
C2250 VDD.n786 VSS 0.03fF $ **FLOATING
C2251 VDD.n787 VSS 0.00fF $ **FLOATING
C2252 VDD.n788 VSS 0.34fF $ **FLOATING
C2253 VDD.n789 VSS 0.03fF $ **FLOATING
C2254 VDD.n790 VSS 0.03fF $ **FLOATING
C2255 sky130_asc_res_xhigh_po_2p85_1_24/VPWR VSS 1.00fF $ **FLOATING
C2256 sky130_asc_res_xhigh_po_2p85_1_21/VPWR VSS 0.99fF $ **FLOATING
C2257 sky130_asc_cap_mim_m3_1_8/VPWR VSS 1.88fF $ **FLOATING
C2258 sky130_asc_res_xhigh_po_2p85_2_0/VPWR VSS 1.99fF $ **FLOATING
C2259 sky130_asc_res_xhigh_po_2p85_1_29/VPWR VSS 1.10fF $ **FLOATING
C2260 sky130_asc_res_xhigh_po_2p85_1_30/VPWR VSS 1.00fF $ **FLOATING
C2261 sky130_asc_res_xhigh_po_2p85_1_10/VPWR VSS 1.00fF $ **FLOATING
C2262 sky130_asc_res_xhigh_po_2p85_1_14/VPWR VSS 1.00fF $ **FLOATING
C2263 sky130_asc_res_xhigh_po_2p85_1_12/VPWR VSS 1.45fF $ **FLOATING
C2264 VDD.n792 VSS 0.81fF $ **FLOATING
C2265 VDD.n793 VSS 0.05fF $ **FLOATING
C2266 VDD.n794 VSS 0.00fF $ **FLOATING
C2267 VDD.n795 VSS 0.05fF $ **FLOATING
C2268 VDD.n796 VSS 0.01fF $ **FLOATING
C2269 VDD.n797 VSS 0.06fF $ **FLOATING
C2270 VDD.n798 VSS 0.00fF $ **FLOATING
C2271 VDD.n799 VSS 0.05fF $ **FLOATING
C2272 VDD.n800 VSS 0.01fF $ **FLOATING
C2273 VDD.n801 VSS 0.06fF $ **FLOATING
C2274 VDD.n802 VSS 0.00fF $ **FLOATING
C2275 VDD.n803 VSS 0.05fF $ **FLOATING
C2276 VDD.n804 VSS 0.01fF $ **FLOATING
C2277 VDD.n805 VSS 0.06fF $ **FLOATING
C2278 VDD.n806 VSS 0.00fF $ **FLOATING
C2279 VDD.n807 VSS 0.05fF $ **FLOATING
C2280 VDD.n808 VSS 0.01fF $ **FLOATING
C2281 VDD.n809 VSS 0.05fF $ **FLOATING
C2282 VDD.n810 VSS 0.01fF $ **FLOATING
C2283 VDD.n811 VSS 0.03fF $ **FLOATING
C2284 VDD.n812 VSS 0.01fF $ **FLOATING
C2285 VDD.n813 VSS 0.03fF $ **FLOATING
C2286 VDD.n814 VSS 0.00fF $ **FLOATING
C2287 VDD.n815 VSS 0.34fF $ **FLOATING
C2288 sky130_asc_res_xhigh_po_2p85_1_27/VPWR VSS 1.10fF $ **FLOATING
C2289 sky130_asc_res_xhigh_po_2p85_1_25/VPWR VSS 1.00fF $ **FLOATING
C2290 sky130_asc_res_xhigh_po_2p85_1_23/VPWR VSS 1.00fF $ **FLOATING
C2291 sky130_asc_res_xhigh_po_2p85_1_26/VPWR VSS 1.00fF $ **FLOATING
C2292 sky130_asc_res_xhigh_po_2p85_1_28/VPWR VSS 1.00fF $ **FLOATING
C2293 sky130_asc_res_xhigh_po_2p85_1_13/VPWR VSS 1.17fF $ **FLOATING
C2294 sky130_asc_res_xhigh_po_2p85_1_11/VPWR VSS 1.09fF $ **FLOATING
C2295 sky130_asc_res_xhigh_po_2p85_1_15/VPWR VSS 1.47fF $ **FLOATING
C2296 VDD.n816 VSS 104.86fF $ **FLOATING
C2297 VDD.n817 VSS 6.43fF $ **FLOATING
C2298 VDD.n818 VSS 0.09fF $ **FLOATING
C2299 VDD.n819 VSS 6.54fF $ **FLOATING
C2300 VDD.n820 VSS 6.43fF $ **FLOATING
C2301 VDD.n821 VSS 0.09fF $ **FLOATING
C2302 VDD.n822 VSS 6.54fF $ **FLOATING
C2303 VDD.n823 VSS 6.43fF $ **FLOATING
C2304 VDD.n824 VSS 0.09fF $ **FLOATING
C2305 VDD.n825 VSS 6.54fF $ **FLOATING
C2306 VDD.n826 VSS 6.43fF $ **FLOATING
C2307 VDD.n827 VSS 0.09fF $ **FLOATING
C2308 VDD.n828 VSS 6.54fF $ **FLOATING
C2309 VDD.n829 VSS 6.43fF $ **FLOATING
C2310 VDD.n830 VSS 0.09fF $ **FLOATING
C2311 VDD.n831 VSS 6.54fF $ **FLOATING
C2312 VDD.n832 VSS 6.43fF $ **FLOATING
C2313 VDD.n833 VSS 0.09fF $ **FLOATING
C2314 VDD.n834 VSS 6.54fF $ **FLOATING
C2315 VDD.n835 VSS 6.43fF $ **FLOATING
C2316 VDD.n836 VSS 0.09fF $ **FLOATING
C2317 VDD.n837 VSS 6.54fF $ **FLOATING
C2318 VDD.n838 VSS 6.43fF $ **FLOATING
C2319 VDD.n839 VSS 0.09fF $ **FLOATING
C2320 VDD.n840 VSS 0.34fF $ **FLOATING
C2321 VDD.n841 VSS 0.00fF $ **FLOATING
C2322 VDD.n842 VSS 0.03fF $ **FLOATING
C2323 VDD.n843 VSS 0.01fF $ **FLOATING
C2324 VDD.n844 VSS 0.03fF $ **FLOATING
C2325 VDD.n845 VSS 0.01fF $ **FLOATING
C2326 VDD.n846 VSS 0.05fF $ **FLOATING
C2327 VDD.n847 VSS 0.01fF $ **FLOATING
C2328 VDD.n848 VSS 0.05fF $ **FLOATING
C2329 VDD.n849 VSS 0.00fF $ **FLOATING
C2330 VDD.n850 VSS 0.06fF $ **FLOATING
C2331 VDD.n851 VSS 0.01fF $ **FLOATING
C2332 VDD.n852 VSS 0.05fF $ **FLOATING
C2333 VDD.n853 VSS 0.00fF $ **FLOATING
C2334 VDD.n854 VSS 0.06fF $ **FLOATING
C2335 VDD.n855 VSS 0.01fF $ **FLOATING
C2336 VDD.n856 VSS 0.05fF $ **FLOATING
C2337 VDD.n857 VSS 0.00fF $ **FLOATING
C2338 VDD.n858 VSS 0.06fF $ **FLOATING
C2339 VDD.n859 VSS 0.01fF $ **FLOATING
C2340 VDD.n860 VSS 0.05fF $ **FLOATING
C2341 VDD.n861 VSS 0.00fF $ **FLOATING
C2342 VDD.n862 VSS 0.05fF $ **FLOATING
C2343 VDD.n863 VSS 0.60fF $ **FLOATING
C2344 sky130_asc_res_xhigh_po_2p85_1_19/VPWR VSS 2.50fF $ **FLOATING
C2345 sky130_asc_pnp_05v5_W3p40L3p40_7_0/VPWR VSS 2.05fF $ **FLOATING
C2346 sky130_asc_nfet_01v8_lvt_1_1/VPWR VSS 0.33fF $ **FLOATING
C2347 VDD.n864 VSS 0.00fF $ **FLOATING
C2348 VDD.n865 VSS 0.00fF $ **FLOATING
C2349 sky130_asc_cap_mim_m3_1_0/Cin VSS 0.03fF $ **FLOATING
C2350 VDD.t348 VSS 1.92fF
C2351 VDD.t13 VSS 2.19fF
C2352 VDD.t57 VSS 2.19fF
C2353 VDD.t349 VSS 2.19fF
C2354 VDD.t14 VSS 2.19fF
C2355 VDD.t107 VSS 2.19fF
C2356 VDD.t312 VSS 2.19fF
C2357 VDD.t343 VSS 2.19fF
C2358 VDD.t229 VSS 2.19fF
C2359 VDD.t36 VSS 2.32fF
C2360 VDD.n866 VSS 0.10fF $ **FLOATING
C2361 VDD.n867 VSS 0.01fF $ **FLOATING
C2362 VDD.n868 VSS -0.01fF $ **FLOATING
C2363 VDD.n869 VSS 0.01fF $ **FLOATING
C2364 VDD.n870 VSS 1.40fF $ **FLOATING
C2365 sky130_asc_cap_mim_m3_1_0/VPWR VSS 2.04fF $ **FLOATING
C2366 VDD.n871 VSS 0.00fF $ **FLOATING
C2367 VDD.n872 VSS 0.00fF $ **FLOATING
C2368 VDD.t17 VSS 2.41fF
C2369 VDD.t144 VSS 2.19fF
C2370 VDD.t304 VSS 2.19fF
C2371 VDD.t87 VSS 2.19fF
C2372 VDD.t265 VSS 1.61fF
C2373 sky130_asc_cap_mim_m3_1_3/Cin VSS 0.03fF $ **FLOATING
C2374 VDD.t20 VSS 1.92fF
C2375 VDD.t141 VSS 2.19fF
C2376 VDD.t264 VSS 2.19fF
C2377 VDD.t12 VSS 2.19fF
C2378 VDD.t9 VSS 1.56fF
C2379 VDD.n873 VSS 1.15fF $ **FLOATING
C2380 VDD.n874 VSS 0.08fF $ **FLOATING
C2381 VDD.n875 VSS 0.01fF $ **FLOATING
C2382 VDD.n876 VSS -0.01fF $ **FLOATING
C2383 VDD.n877 VSS 0.01fF $ **FLOATING
C2384 VDD.n878 VSS 1.40fF $ **FLOATING
C2385 sky130_asc_cap_mim_m3_1_3/VPWR VSS 0.71fF $ **FLOATING
C2386 VDD.n879 VSS 0.00fF $ **FLOATING
C2387 VDD.n880 VSS 0.00fF $ **FLOATING
C2388 sky130_asc_cap_mim_m3_1_1/Cin VSS 0.03fF $ **FLOATING
C2389 VDD.t37 VSS 1.92fF
C2390 VDD.t91 VSS 2.19fF
C2391 VDD.t309 VSS 2.19fF
C2392 VDD.t124 VSS 2.19fF
C2393 VDD.t202 VSS 2.19fF
C2394 VDD.t72 VSS 2.19fF
C2395 VDD.t88 VSS 2.19fF
C2396 VDD.t23 VSS 2.19fF
C2397 VDD.t143 VSS 2.19fF
C2398 VDD.t340 VSS 2.32fF
C2399 VDD.n881 VSS 0.10fF $ **FLOATING
C2400 VDD.n882 VSS 0.01fF $ **FLOATING
C2401 VDD.n883 VSS -0.01fF $ **FLOATING
C2402 VDD.n884 VSS 0.01fF $ **FLOATING
C2403 VDD.n885 VSS 1.39fF $ **FLOATING
C2404 sky130_asc_cap_mim_m3_1_1/VPWR VSS 1.51fF $ **FLOATING
C2405 sky130_asc_nfet_01v8_lvt_1_0/VPWR VSS 0.34fF $ **FLOATING
C2406 VDD.n887 VSS 0.05fF $ **FLOATING
C2407 VDD.n888 VSS 0.01fF $ **FLOATING
C2408 VDD.n889 VSS 0.06fF $ **FLOATING
C2409 VDD.n890 VSS 0.00fF $ **FLOATING
C2410 VDD.n892 VSS 0.13fF $ **FLOATING
C2411 VDD.n893 VSS 6.54fF $ **FLOATING
C2412 VDD.n894 VSS 6.37fF $ **FLOATING
C2413 VDD.n895 VSS 0.00fF $ **FLOATING
C2414 VDD.n897 VSS 0.03fF $ **FLOATING
C2415 VDD.n898 VSS 0.01fF $ **FLOATING
C2416 VDD.n899 VSS 0.03fF $ **FLOATING
C2417 VDD.n900 VSS 0.01fF $ **FLOATING
C2418 VDD.n901 VSS 0.06fF $ **FLOATING
C2419 VDD.n902 VSS 0.01fF $ **FLOATING
C2420 VDD.n903 VSS 0.05fF $ **FLOATING
C2421 VDD.n904 VSS 0.00fF $ **FLOATING
C2422 VDD.n906 VSS 0.06fF $ **FLOATING
C2423 VDD.n907 VSS 0.01fF $ **FLOATING
C2424 VDD.n908 VSS 0.05fF $ **FLOATING
C2425 VDD.n909 VSS 0.00fF $ **FLOATING
C2426 VDD.n910 VSS 0.06fF $ **FLOATING
C2427 VDD.n911 VSS 0.00fF $ **FLOATING
C2428 VDD.n912 VSS 0.03fF $ **FLOATING
C2429 VDD.n913 VSS 0.03fF $ **FLOATING
C2430 VDD.n914 VSS 0.01fF $ **FLOATING
C2431 VDD.n915 VSS 0.05fF $ **FLOATING
C2432 VDD.n916 VSS 0.01fF $ **FLOATING
C2433 VDD.n917 VSS 0.05fF $ **FLOATING
C2434 VDD.n918 VSS 0.06fF $ **FLOATING
C2435 VDD.n919 VSS 0.00fF $ **FLOATING
C2436 VDD.n920 VSS 0.01fF $ **FLOATING
C2437 VDD.n921 VSS 0.05fF $ **FLOATING
C2438 VDD.n922 VSS 0.06fF $ **FLOATING
C2439 VDD.n923 VSS 0.00fF $ **FLOATING
C2440 VDD.n924 VSS 0.01fF $ **FLOATING
C2441 VDD.n925 VSS 0.05fF $ **FLOATING
C2442 VDD.t266 VSS 1.80fF
C2443 VDD.t268 VSS 1.58fF
C2444 VDD.t136 VSS 1.58fF
C2445 VDD.t278 VSS 1.10fF
C2446 VDD.t151 VSS 1.27fF
C2447 VDD.n927 VSS 0.79fF $ **FLOATING
C2448 VDD.n928 VSS 0.07fF $ **FLOATING
C2449 VDD.t263 VSS 0.04fF
C2450 VDD.t131 VSS 0.04fF
C2451 VDD.n929 VSS 0.29fF $ **FLOATING
C2452 VDD.t247 VSS 0.04fF
C2453 VDD.t259 VSS 0.04fF
C2454 VDD.n930 VSS 0.29fF $ **FLOATING
C2455 VDD.t193 VSS 0.04fF
C2456 VDD.t195 VSS 0.04fF
C2457 VDD.n931 VSS 0.29fF $ **FLOATING
C2458 VDD.t289 VSS 0.04fF
C2459 VDD.t293 VSS 0.04fF
C2460 VDD.n932 VSS 0.29fF $ **FLOATING
C2461 VDD.t62 VSS 0.04fF
C2462 VDD.t25 VSS 0.04fF
C2463 VDD.n933 VSS 0.29fF $ **FLOATING
C2464 VDD.t185 VSS 0.04fF
C2465 VDD.t187 VSS 0.04fF
C2466 VDD.n934 VSS 0.29fF $ **FLOATING
C2467 VDD.t166 VSS 0.04fF
C2468 VDD.t100 VSS 0.04fF
C2469 VDD.n935 VSS 0.29fF $ **FLOATING
C2470 VDD.t224 VSS 0.04fF
C2471 VDD.t86 VSS 0.04fF
C2472 VDD.n936 VSS 0.29fF $ **FLOATING
C2473 VDD.t158 VSS 0.04fF
C2474 VDD.t220 VSS 0.04fF
C2475 VDD.n937 VSS 0.29fF $ **FLOATING
C2476 VDD.t117 VSS 0.04fF
C2477 VDD.t156 VSS 0.04fF
C2478 VDD.n938 VSS 0.29fF $ **FLOATING
C2479 VDD.t253 VSS 0.04fF
C2480 VDD.t303 VSS 0.04fF
C2481 VDD.n939 VSS 0.29fF $ **FLOATING
C2482 VDD.t237 VSS 0.04fF
C2483 VDD.t369 VSS 0.04fF
C2484 VDD.n940 VSS 0.29fF $ **FLOATING
C2485 VDD.t327 VSS 0.04fF
C2486 VDD.t235 VSS 0.04fF
C2487 VDD.n941 VSS 0.29fF $ **FLOATING
C2488 VDD.t391 VSS 0.04fF
C2489 VDD.t324 VSS 0.04fF
C2490 VDD.n942 VSS 0.29fF $ **FLOATING
C2491 VDD.t383 VSS 0.04fF
C2492 VDD.t273 VSS 0.04fF
C2493 VDD.n943 VSS 0.29fF $ **FLOATING
C2494 VDD.t152 VSS 0.04fF
C2495 VDD.t342 VSS 0.04fF
C2496 VDD.n944 VSS 0.29fF $ **FLOATING
C2497 VDD.t137 VSS 0.04fF
C2498 VDD.t279 VSS 0.04fF
C2499 VDD.n945 VSS 0.29fF $ **FLOATING
C2500 VDD.t267 VSS 0.04fF
C2501 VDD.t269 VSS 0.04fF
C2502 VDD.n946 VSS 0.29fF $ **FLOATING
C2503 sky130_asc_pfet_01v8_lvt_60_0/SOURCE VSS 0.02fF $ **FLOATING
C2504 VDD.n947 VSS 0.06fF $ **FLOATING
C2505 VDD.n948 VSS 0.08fF $ **FLOATING
C2506 VDD.n949 VSS 0.08fF $ **FLOATING
C2507 VDD.n950 VSS 0.08fF $ **FLOATING
C2508 VDD.n951 VSS 0.08fF $ **FLOATING
C2509 VDD.n952 VSS 0.08fF $ **FLOATING
C2510 VDD.n953 VSS 0.08fF $ **FLOATING
C2511 VDD.n954 VSS 0.08fF $ **FLOATING
C2512 VDD.n955 VSS 0.08fF $ **FLOATING
C2513 VDD.n956 VSS 0.08fF $ **FLOATING
C2514 VDD.n957 VSS 0.08fF $ **FLOATING
C2515 VDD.n958 VSS 0.08fF $ **FLOATING
C2516 VDD.n959 VSS 0.08fF $ **FLOATING
C2517 VDD.n960 VSS 0.08fF $ **FLOATING
C2518 VDD.n961 VSS 0.08fF $ **FLOATING
C2519 VDD.n962 VSS 0.08fF $ **FLOATING
C2520 VDD.n963 VSS 0.08fF $ **FLOATING
C2521 VDD.n964 VSS 0.08fF $ **FLOATING
C2522 VDD.t171 VSS 0.04fF
C2523 VDD.t231 VSS 0.04fF
C2524 VDD.n965 VSS 0.29fF $ **FLOATING
C2525 VDD.t33 VSS 0.04fF
C2526 VDD.t93 VSS 0.04fF
C2527 VDD.n966 VSS 0.29fF $ **FLOATING
C2528 VDD.t385 VSS 0.04fF
C2529 VDD.t106 VSS 0.04fF
C2530 VDD.n967 VSS 0.29fF $ **FLOATING
C2531 VDD.t109 VSS 0.04fF
C2532 VDD.t421 VSS 0.04fF
C2533 VDD.n968 VSS 0.29fF $ **FLOATING
C2534 VDD.t67 VSS 0.04fF
C2535 VDD.t357 VSS 0.04fF
C2536 VDD.n969 VSS 0.29fF $ **FLOATING
C2537 VDD.t74 VSS 0.04fF
C2538 VDD.t113 VSS 0.04fF
C2539 VDD.n970 VSS 0.29fF $ **FLOATING
C2540 VDD.t154 VSS 0.04fF
C2541 VDD.t199 VSS 0.04fF
C2542 VDD.n971 VSS 0.29fF $ **FLOATING
C2543 VDD.t51 VSS 0.04fF
C2544 VDD.t146 VSS 0.04fF
C2545 VDD.n972 VSS 0.29fF $ **FLOATING
C2546 VDD.t78 VSS 0.04fF
C2547 VDD.t84 VSS 0.04fF
C2548 VDD.n973 VSS 0.29fF $ **FLOATING
C2549 VDD.t162 VSS 0.04fF
C2550 VDD.t437 VSS 0.04fF
C2551 VDD.n974 VSS 0.29fF $ **FLOATING
C2552 VDD.t183 VSS 0.04fF
C2553 VDD.t41 VSS 0.04fF
C2554 VDD.n975 VSS 0.37fF $ **FLOATING
C2555 VDD.n976 VSS 0.09fF $ **FLOATING
C2556 VDD.n977 VSS 0.08fF $ **FLOATING
C2557 VDD.n978 VSS 0.08fF $ **FLOATING
C2558 VDD.n979 VSS 0.08fF $ **FLOATING
C2559 VDD.n980 VSS 0.08fF $ **FLOATING
C2560 VDD.n981 VSS 0.08fF $ **FLOATING
C2561 VDD.n982 VSS 0.08fF $ **FLOATING
C2562 VDD.n983 VSS 0.08fF $ **FLOATING
C2563 VDD.n984 VSS 0.08fF $ **FLOATING
C2564 VDD.n985 VSS 0.08fF $ **FLOATING
C2565 VDD.n986 VSS 0.08fF $ **FLOATING
C2566 VDD.t127 VSS 0.04fF
C2567 VDD.t214 VSS 0.04fF
C2568 VDD.n987 VSS 0.20fF $ **FLOATING
C2569 VDD.n988 VSS 0.06fF $ **FLOATING
C2570 sky130_asc_cap_mim_m3_1_4/VPWR VSS 1.19fF $ **FLOATING
C2571 VDD.t18 VSS 2.41fF
C2572 VDD.t8 VSS 1.61fF
C2573 sky130_asc_cap_mim_m3_1_4/Cin VSS 0.03fF $ **FLOATING
C2574 VDD.t19 VSS 1.92fF
C2575 VDD.t140 VSS 2.19fF
C2576 VDD.t335 VSS 2.19fF
C2577 VDD.t21 VSS 2.19fF
C2578 VDD.t16 VSS 2.19fF
C2579 VDD.t125 VSS 2.19fF
C2580 VDD.t167 VSS 2.19fF
C2581 VDD.t11 VSS 1.56fF
C2582 VDD.n989 VSS 1.24fF $ **FLOATING
C2583 VDD.n990 VSS 1.57fF $ **FLOATING
C2584 VDD.n991 VSS 0.11fF $ **FLOATING
C2585 VDD.n992 VSS 0.08fF $ **FLOATING
C2586 VDD.n993 VSS 0.45fF $ **FLOATING
C2587 VDD.n994 VSS 0.05fF $ **FLOATING
C2588 VDD.n995 VSS 0.10fF $ **FLOATING
C2589 VDD.t161 VSS 1.58fF
C2590 VDD.t436 VSS 1.05fF
C2591 VDD.t40 VSS 2.01fF
C2592 VDD.t182 VSS 1.32fF
C2593 VDD.n996 VSS 0.79fF $ **FLOATING
C2594 VDD.n997 VSS 0.05fF $ **FLOATING
C2595 VDD.n998 VSS 0.04fF $ **FLOATING
C2596 VDD.n999 VSS 0.10fF $ **FLOATING
C2597 VDD.n1000 VSS 0.04fF $ **FLOATING
C2598 VDD.n1001 VSS 0.10fF $ **FLOATING
C2599 VDD.n1002 VSS 0.05fF $ **FLOATING
C2600 VDD.n1003 VSS 0.10fF $ **FLOATING
C2601 VDD.t77 VSS 1.17fF
C2602 VDD.t83 VSS 1.19fF
C2603 VDD.n1004 VSS 0.79fF $ **FLOATING
C2604 VDD.n1005 VSS 0.06fF $ **FLOATING
C2605 VDD.n1006 VSS 0.04fF $ **FLOATING
C2606 VDD.n1007 VSS 0.10fF $ **FLOATING
C2607 VDD.n1008 VSS 0.04fF $ **FLOATING
C2608 VDD.n1009 VSS 0.10fF $ **FLOATING
C2609 VDD.n1010 VSS 0.05fF $ **FLOATING
C2610 VDD.n1011 VSS 0.10fF $ **FLOATING
C2611 VDD.n1012 VSS 0.04fF $ **FLOATING
C2612 VDD.n1013 VSS 0.10fF $ **FLOATING
C2613 VDD.t198 VSS 1.30fF
C2614 VDD.t145 VSS 1.58fF
C2615 VDD.t50 VSS 1.07fF
C2616 VDD.n1014 VSS 0.79fF $ **FLOATING
C2617 VDD.n1015 VSS 0.06fF $ **FLOATING
C2618 VDD.n1016 VSS 0.03fF $ **FLOATING
C2619 VDD.n1017 VSS 0.10fF $ **FLOATING
C2620 VDD.n1018 VSS 0.05fF $ **FLOATING
C2621 VDD.n1019 VSS 0.10fF $ **FLOATING
C2622 VDD.n1020 VSS 0.05fF $ **FLOATING
C2623 VDD.n1021 VSS 0.10fF $ **FLOATING
C2624 VDD.t73 VSS 1.43fF
C2625 VDD.t153 VSS 1.58fF
C2626 VDD.t112 VSS 0.94fF
C2627 VDD.n1022 VSS 0.79fF $ **FLOATING
C2628 VDD.n1023 VSS 0.05fF $ **FLOATING
C2629 VDD.n1024 VSS 0.04fF $ **FLOATING
C2630 VDD.n1025 VSS 0.10fF $ **FLOATING
C2631 VDD.n1026 VSS 0.05fF $ **FLOATING
C2632 VDD.n1027 VSS 0.10fF $ **FLOATING
C2633 VDD.n1028 VSS 0.05fF $ **FLOATING
C2634 VDD.n1029 VSS 0.10fF $ **FLOATING
C2635 VDD.t420 VSS 1.56fF
C2636 VDD.t356 VSS 1.58fF
C2637 VDD.t66 VSS 0.81fF
C2638 VDD.n1030 VSS 0.79fF $ **FLOATING
C2639 VDD.n1031 VSS 0.05fF $ **FLOATING
C2640 VDD.n1032 VSS 0.04fF $ **FLOATING
C2641 VDD.n1033 VSS 0.10fF $ **FLOATING
C2642 VDD.n1034 VSS 0.04fF $ **FLOATING
C2643 VDD.n1035 VSS 0.10fF $ **FLOATING
C2644 VDD.n1036 VSS 0.05fF $ **FLOATING
C2645 VDD.n1037 VSS 0.10fF $ **FLOATING
C2646 VDD.t384 VSS 1.58fF
C2647 VDD.t105 VSS 0.89fF
C2648 VDD.t108 VSS 1.47fF
C2649 VDD.n1038 VSS 0.79fF $ **FLOATING
C2650 VDD.n1039 VSS 0.06fF $ **FLOATING
C2651 VDD.n1040 VSS 0.04fF $ **FLOATING
C2652 VDD.n1041 VSS 0.10fF $ **FLOATING
C2653 VDD.n1042 VSS 0.04fF $ **FLOATING
C2654 VDD.n1043 VSS 0.10fF $ **FLOATING
C2655 VDD.n1044 VSS 0.05fF $ **FLOATING
C2656 VDD.n1045 VSS 0.10fF $ **FLOATING
C2657 VDD.n1046 VSS 0.04fF $ **FLOATING
C2658 VDD.n1047 VSS 0.10fF $ **FLOATING
C2659 VDD.t230 VSS 1.58fF
C2660 VDD.t32 VSS 1.02fF
C2661 VDD.t92 VSS 1.35fF
C2662 VDD.n1048 VSS 0.79fF $ **FLOATING
C2663 VDD.n1049 VSS 0.06fF $ **FLOATING
C2664 VDD.n1050 VSS 0.03fF $ **FLOATING
C2665 VDD.n1051 VSS 0.10fF $ **FLOATING
C2666 VDD.n1052 VSS 0.05fF $ **FLOATING
C2667 VDD.n1053 VSS 0.10fF $ **FLOATING
C2668 VDD.n1054 VSS 0.05fF $ **FLOATING
C2669 VDD.n1055 VSS 0.10fF $ **FLOATING
C2670 VDD.t213 VSS 1.15fF
C2671 VDD.t170 VSS 1.22fF
C2672 VDD.n1056 VSS 0.79fF $ **FLOATING
C2673 VDD.n1057 VSS 0.05fF $ **FLOATING
C2674 VDD.n1058 VSS 0.04fF $ **FLOATING
C2675 VDD.n1059 VSS 0.10fF $ **FLOATING
C2676 VDD.n1060 VSS 0.09fF $ **FLOATING
C2677 VDD.n1061 VSS 0.05fF $ **FLOATING
C2678 VDD.n1062 VSS 0.05fF $ **FLOATING
C2679 VDD.n1063 VSS 0.05fF $ **FLOATING
C2680 VDD.n1064 VSS 0.10fF $ **FLOATING
C2681 VDD.t262 VSS 1.28fF
C2682 VDD.t126 VSS 1.58fF
C2683 VDD.t130 VSS 1.09fF
C2684 VDD.n1065 VSS 0.79fF $ **FLOATING
C2685 VDD.n1066 VSS 0.05fF $ **FLOATING
C2686 VDD.n1067 VSS 0.04fF $ **FLOATING
C2687 VDD.n1068 VSS 0.10fF $ **FLOATING
C2688 VDD.n1069 VSS 0.04fF $ **FLOATING
C2689 VDD.n1070 VSS 0.10fF $ **FLOATING
C2690 VDD.n1071 VSS 0.05fF $ **FLOATING
C2691 VDD.n1072 VSS 0.10fF $ **FLOATING
C2692 VDD.t194 VSS 1.40fF
C2693 VDD.t258 VSS 1.58fF
C2694 VDD.t246 VSS 0.96fF
C2695 VDD.n1073 VSS 0.79fF $ **FLOATING
C2696 VDD.n1074 VSS 0.06fF $ **FLOATING
C2697 VDD.n1075 VSS 0.04fF $ **FLOATING
C2698 VDD.n1076 VSS 0.10fF $ **FLOATING
C2699 VDD.n1077 VSS 0.04fF $ **FLOATING
C2700 VDD.n1078 VSS 0.10fF $ **FLOATING
C2701 VDD.n1079 VSS 0.05fF $ **FLOATING
C2702 VDD.n1080 VSS 0.10fF $ **FLOATING
C2703 VDD.n1081 VSS 0.04fF $ **FLOATING
C2704 VDD.n1082 VSS 0.10fF $ **FLOATING
C2705 VDD.t288 VSS 1.53fF
C2706 VDD.t192 VSS 1.58fF
C2707 VDD.t292 VSS 0.84fF
C2708 VDD.n1083 VSS 0.79fF $ **FLOATING
C2709 VDD.n1084 VSS 0.06fF $ **FLOATING
C2710 VDD.n1085 VSS 0.03fF $ **FLOATING
C2711 VDD.n1086 VSS 0.10fF $ **FLOATING
C2712 VDD.n1087 VSS 0.05fF $ **FLOATING
C2713 VDD.n1088 VSS 0.10fF $ **FLOATING
C2714 VDD.n1089 VSS 0.05fF $ **FLOATING
C2715 VDD.n1090 VSS 0.10fF $ **FLOATING
C2716 VDD.t186 VSS 1.58fF
C2717 VDD.t61 VSS 0.87fF
C2718 VDD.t24 VSS 1.50fF
C2719 VDD.n1091 VSS 0.79fF $ **FLOATING
C2720 VDD.n1092 VSS 0.05fF $ **FLOATING
C2721 VDD.n1093 VSS 0.04fF $ **FLOATING
C2722 VDD.n1094 VSS 0.10fF $ **FLOATING
C2723 VDD.n1095 VSS 0.05fF $ **FLOATING
C2724 VDD.n1096 VSS 0.10fF $ **FLOATING
C2725 VDD.n1097 VSS 0.05fF $ **FLOATING
C2726 VDD.n1098 VSS 0.10fF $ **FLOATING
C2727 VDD.t165 VSS 1.58fF
C2728 VDD.t99 VSS 1.00fF
C2729 VDD.t184 VSS 1.37fF
C2730 VDD.n1099 VSS 0.79fF $ **FLOATING
C2731 VDD.n1100 VSS 0.05fF $ **FLOATING
C2732 VDD.n1101 VSS 0.04fF $ **FLOATING
C2733 VDD.n1102 VSS 0.10fF $ **FLOATING
C2734 VDD.n1103 VSS 0.04fF $ **FLOATING
C2735 VDD.n1104 VSS 0.10fF $ **FLOATING
C2736 VDD.n1105 VSS 0.05fF $ **FLOATING
C2737 VDD.n1106 VSS 0.10fF $ **FLOATING
C2738 VDD.t223 VSS 1.13fF
C2739 VDD.t85 VSS 1.24fF
C2740 VDD.n1107 VSS 0.79fF $ **FLOATING
C2741 VDD.n1108 VSS 0.06fF $ **FLOATING
C2742 VDD.n1109 VSS 0.04fF $ **FLOATING
C2743 VDD.n1110 VSS 0.10fF $ **FLOATING
C2744 VDD.n1111 VSS 0.04fF $ **FLOATING
C2745 VDD.n1112 VSS 0.10fF $ **FLOATING
C2746 VDD.n1113 VSS 0.05fF $ **FLOATING
C2747 VDD.n1114 VSS 0.10fF $ **FLOATING
C2748 VDD.n1115 VSS 0.04fF $ **FLOATING
C2749 VDD.n1116 VSS 0.10fF $ **FLOATING
C2750 VDD.t155 VSS 1.25fF
C2751 VDD.t219 VSS 1.58fF
C2752 VDD.t157 VSS 1.11fF
C2753 VDD.n1117 VSS 0.79fF $ **FLOATING
C2754 VDD.n1118 VSS 0.06fF $ **FLOATING
C2755 VDD.n1119 VSS 0.03fF $ **FLOATING
C2756 VDD.n1120 VSS 0.10fF $ **FLOATING
C2757 VDD.n1121 VSS 0.05fF $ **FLOATING
C2758 VDD.n1122 VSS 0.10fF $ **FLOATING
C2759 VDD.n1123 VSS 0.05fF $ **FLOATING
C2760 VDD.n1124 VSS 0.10fF $ **FLOATING
C2761 VDD.t252 VSS 1.38fF
C2762 VDD.t116 VSS 1.58fF
C2763 VDD.t302 VSS 0.99fF
C2764 VDD.n1125 VSS 0.79fF $ **FLOATING
C2765 VDD.n1126 VSS 0.05fF $ **FLOATING
C2766 VDD.n1127 VSS 0.04fF $ **FLOATING
C2767 VDD.n1128 VSS 0.10fF $ **FLOATING
C2768 VDD.n1129 VSS 0.05fF $ **FLOATING
C2769 VDD.n1130 VSS 0.10fF $ **FLOATING
C2770 VDD.n1131 VSS 0.05fF $ **FLOATING
C2771 VDD.n1132 VSS 0.10fF $ **FLOATING
C2772 VDD.t234 VSS 1.51fF
C2773 VDD.t368 VSS 1.58fF
C2774 VDD.t236 VSS 0.86fF
C2775 VDD.n1133 VSS 0.79fF $ **FLOATING
C2776 VDD.n1134 VSS 0.05fF $ **FLOATING
C2777 VDD.n1135 VSS 0.04fF $ **FLOATING
C2778 VDD.n1136 VSS 0.10fF $ **FLOATING
C2779 VDD.n1137 VSS 0.04fF $ **FLOATING
C2780 VDD.n1138 VSS 0.10fF $ **FLOATING
C2781 VDD.n1139 VSS 0.05fF $ **FLOATING
C2782 VDD.n1140 VSS 0.10fF $ **FLOATING
C2783 VDD.t390 VSS 1.58fF
C2784 VDD.t323 VSS 0.85fF
C2785 VDD.t326 VSS 1.52fF
C2786 VDD.n1141 VSS 0.79fF $ **FLOATING
C2787 VDD.n1142 VSS 0.06fF $ **FLOATING
C2788 VDD.n1143 VSS 0.04fF $ **FLOATING
C2789 VDD.n1144 VSS 0.10fF $ **FLOATING
C2790 VDD.n1145 VSS 0.04fF $ **FLOATING
C2791 VDD.n1146 VSS 0.10fF $ **FLOATING
C2792 VDD.n1147 VSS 0.05fF $ **FLOATING
C2793 VDD.n1148 VSS 0.10fF $ **FLOATING
C2794 VDD.n1149 VSS 0.04fF $ **FLOATING
C2795 VDD.n1150 VSS 0.10fF $ **FLOATING
C2796 VDD.t341 VSS 1.58fF
C2797 VDD.t382 VSS 0.97fF
C2798 VDD.t272 VSS 1.39fF
C2799 VDD.n1151 VSS 0.79fF $ **FLOATING
C2800 VDD.n1152 VSS 0.06fF $ **FLOATING
C2801 VDD.n1153 VSS 0.03fF $ **FLOATING
C2802 VDD.n1154 VSS 0.10fF $ **FLOATING
C2803 VDD.n1155 VSS 0.05fF $ **FLOATING
C2804 VDD.n1156 VSS 0.10fF $ **FLOATING
C2805 VDD.n1157 VSS 0.05fF $ **FLOATING
C2806 VDD.n1158 VSS 0.11fF $ **FLOATING
C2807 VDD.n1159 VSS 0.56fF $ **FLOATING
C2808 VDD.n1160 VSS 0.44fF $ **FLOATING
C2809 VDD.n1161 VSS 0.04fF $ **FLOATING
C2810 VDD.n1162 VSS 0.01fF $ **FLOATING
C2811 VDD.n1163 VSS 0.06fF $ **FLOATING
C2812 VDD.n1164 VSS 0.01fF $ **FLOATING
C2813 VDD.n1165 VSS 0.06fF $ **FLOATING
C2814 VDD.n1166 VSS 0.00fF $ **FLOATING
C2815 VDD.n1167 VSS 102.87fF $ **FLOATING
C2816 VDD.n1168 VSS 110.44fF $ **FLOATING
C2817 VDD.n1169 VSS 14.13fF $ **FLOATING
C2818 VDD.n1170 VSS 14.23fF $ **FLOATING
C2819 VDD.n1171 VSS 14.17fF $ **FLOATING
C2820 VDD.n1172 VSS 14.25fF $ **FLOATING
C2821 VDD.n1173 VSS 14.40fF $ **FLOATING
C2822 VDD.n1174 VSS 14.14fF $ **FLOATING
C2823 VDD.n1175 VSS 14.40fF $ **FLOATING
C2824 VDD.n1176 VSS 14.40fF $ **FLOATING
C2825 VDD.n1177 VSS 14.03fF $ **FLOATING
C2826 sky130_asc_res_xhigh_po_2p85_1_1/VPWR VSS 1.44fF $ **FLOATING
C2827 sky130_asc_pfet_01v8_lvt_60_0/GATE.n0 VSS 0.04fF $ **FLOATING
C2828 sky130_asc_pfet_01v8_lvt_60_0/GATE.t40 VSS 6.86fF
C2829 sky130_asc_pfet_01v8_lvt_60_0/GATE.n1 VSS 0.02fF $ **FLOATING
C2830 sky130_asc_pfet_01v8_lvt_60_0/GATE.n2 VSS 0.02fF $ **FLOATING
C2831 sky130_asc_pfet_01v8_lvt_60_0/GATE.t89 VSS 5.09fF
C2832 sky130_asc_cap_mim_m3_1_3/Cout VSS 4.46fF
C2833 sky130_asc_pfet_01v8_lvt_60_0/GATE.n3 VSS 0.01fF $ **FLOATING
C2834 sky130_asc_pfet_01v8_lvt_60_0/GATE.n4 VSS 0.40fF $ **FLOATING
C2835 sky130_asc_pfet_01v8_lvt_60_0/GATE.t75 VSS 4.46fF
C2836 sky130_asc_pfet_01v8_lvt_60_0/GATE.t157 VSS 5.03fF
C2837 sky130_asc_pfet_01v8_lvt_60_0/GATE.t27 VSS 5.10fF
C2838 sky130_asc_pfet_01v8_lvt_60_0/GATE.t93 VSS 5.10fF
C2839 sky130_asc_pfet_01v8_lvt_60_0/GATE.t33 VSS 4.39fF
C2840 sky130_asc_pfet_01v8_lvt_60_0/GATE.t43 VSS 5.10fF
C2841 sky130_asc_pfet_01v8_lvt_60_0/GATE.t34 VSS 5.10fF
C2842 sky130_asc_pfet_01v8_lvt_60_0/GATE.t97 VSS 4.39fF
C2843 sky130_asc_pfet_01v8_lvt_60_0/GATE.t73 VSS 5.10fF
C2844 sky130_asc_pfet_01v8_lvt_60_0/GATE.t55 VSS 5.11fF
C2845 sky130_asc_pfet_01v8_lvt_60_0/GATE.t106 VSS 4.30fF
C2846 sky130_asc_pfet_01v8_lvt_60_0/GATE.t46 VSS 3.85fF
C2847 sky130_asc_pfet_01v8_lvt_60_0/GATE.t26 VSS 5.11fF
C2848 sky130_asc_pfet_01v8_lvt_60_0/GATE.t50 VSS 5.10fF
C2849 sky130_asc_pfet_01v8_lvt_60_0/GATE.t109 VSS 5.10fF
C2850 sky130_asc_pfet_01v8_lvt_60_0/GATE.t54 VSS 4.39fF
C2851 sky130_asc_pfet_01v8_lvt_60_0/GATE.t155 VSS 4.14fF
C2852 sky130_asc_pfet_01v8_lvt_60_0/GATE.t81 VSS 5.11fF
C2853 sky130_asc_pfet_01v8_lvt_60_0/GATE.t44 VSS 5.10fF
C2854 sky130_asc_pfet_01v8_lvt_60_0/GATE.t162 VSS 5.10fF
C2855 sky130_asc_pfet_01v8_lvt_60_0/GATE.t38 VSS 4.39fF
C2856 sky130_asc_pfet_01v8_lvt_60_0/GATE.t130 VSS 2.08fF
C2857 sky130_asc_pfet_01v8_lvt_60_0/GATE.t36 VSS 2.08fF
C2858 sky130_asc_pfet_01v8_lvt_60_0/GATE.t72 VSS 2.08fF
C2859 sky130_asc_pfet_01v8_lvt_60_0/GATE.t51 VSS 2.08fF
C2860 sky130_asc_pfet_01v8_lvt_60_0/GATE.t21 VSS 0.52fF
C2861 sky130_asc_pfet_01v8_lvt_60_0/GATE.t20 VSS 0.06fF
C2862 sky130_asc_pfet_01v8_lvt_60_0/GATE.t19 VSS 0.06fF
C2863 sky130_asc_pfet_01v8_lvt_60_0/GATE.n5 VSS 0.44fF $ **FLOATING
C2864 sky130_asc_pfet_01v8_lvt_60_0/GATE.t18 VSS 0.06fF
C2865 sky130_asc_pfet_01v8_lvt_60_0/GATE.t7 VSS 0.06fF
C2866 sky130_asc_pfet_01v8_lvt_60_0/GATE.n6 VSS 0.44fF $ **FLOATING
C2867 sky130_asc_pfet_01v8_lvt_60_0/GATE.t11 VSS 0.04fF
C2868 sky130_asc_pfet_01v8_lvt_60_0/GATE.t15 VSS 0.04fF
C2869 sky130_asc_pfet_01v8_lvt_60_0/GATE.n7 VSS 0.27fF $ **FLOATING
C2870 sky130_asc_pfet_01v8_lvt_60_0/GATE.t10 VSS 0.04fF
C2871 sky130_asc_pfet_01v8_lvt_60_0/GATE.t13 VSS 0.04fF
C2872 sky130_asc_pfet_01v8_lvt_60_0/GATE.n8 VSS 0.27fF $ **FLOATING
C2873 sky130_asc_pfet_01v8_lvt_60_0/GATE.t9 VSS 0.04fF
C2874 sky130_asc_pfet_01v8_lvt_60_0/GATE.t14 VSS 0.04fF
C2875 sky130_asc_pfet_01v8_lvt_60_0/GATE.n9 VSS 0.27fF $ **FLOATING
C2876 sky130_asc_pfet_01v8_lvt_60_0/GATE.t17 VSS 0.04fF
C2877 sky130_asc_pfet_01v8_lvt_60_0/GATE.t12 VSS 0.04fF
C2878 sky130_asc_pfet_01v8_lvt_60_0/GATE.n10 VSS 0.27fF $ **FLOATING
C2879 sky130_asc_nfet_01v8_lvt_9_1/DRAIN VSS 0.05fF $ **FLOATING
C2880 sky130_asc_pfet_01v8_lvt_60_0/GATE.n11 VSS 0.14fF $ **FLOATING
C2881 sky130_asc_pfet_01v8_lvt_60_0/GATE.n12 VSS 0.18fF $ **FLOATING
C2882 sky130_asc_pfet_01v8_lvt_60_0/GATE.n13 VSS 0.18fF $ **FLOATING
C2883 sky130_asc_pfet_01v8_lvt_60_0/GATE.n14 VSS 0.14fF $ **FLOATING
C2884 sky130_asc_pfet_01v8_lvt_60_0/GATE.t16 VSS 0.37fF
C2885 sky130_asc_pfet_01v8_lvt_60_0/GATE.n15 VSS 0.12fF $ **FLOATING
C2886 sky130_asc_pfet_01v8_lvt_60_2/GATE VSS 0.03fF $ **FLOATING
C2887 sky130_asc_pfet_01v8_lvt_60_0/GATE.n16 VSS 0.09fF $ **FLOATING
C2888 sky130_asc_pfet_01v8_lvt_60_0/GATE.t207 VSS 1.44fF
C2889 sky130_asc_pfet_01v8_lvt_60_0/GATE.n17 VSS 0.37fF $ **FLOATING
C2890 sky130_asc_pfet_01v8_lvt_60_0/GATE.n18 VSS 0.05fF $ **FLOATING
C2891 sky130_asc_pfet_01v8_lvt_60_0/GATE.n19 VSS 0.08fF $ **FLOATING
C2892 sky130_asc_pfet_01v8_lvt_60_0/GATE.t127 VSS 1.44fF
C2893 sky130_asc_pfet_01v8_lvt_60_0/GATE.n20 VSS 0.33fF $ **FLOATING
C2894 sky130_asc_pfet_01v8_lvt_60_0/GATE.n21 VSS 0.05fF $ **FLOATING
C2895 sky130_asc_pfet_01v8_lvt_60_0/GATE.n22 VSS 0.08fF $ **FLOATING
C2896 sky130_asc_pfet_01v8_lvt_60_0/GATE.t194 VSS 1.44fF
C2897 sky130_asc_pfet_01v8_lvt_60_0/GATE.n23 VSS 0.33fF $ **FLOATING
C2898 sky130_asc_pfet_01v8_lvt_60_0/GATE.n24 VSS 0.05fF $ **FLOATING
C2899 sky130_asc_pfet_01v8_lvt_60_0/GATE.n25 VSS 0.08fF $ **FLOATING
C2900 sky130_asc_pfet_01v8_lvt_60_0/GATE.t193 VSS 1.44fF
C2901 sky130_asc_pfet_01v8_lvt_60_0/GATE.n26 VSS 0.38fF $ **FLOATING
C2902 sky130_asc_pfet_01v8_lvt_60_0/GATE.n27 VSS 0.08fF $ **FLOATING
C2903 sky130_asc_pfet_01v8_lvt_60_0/GATE.t156 VSS 1.44fF
C2904 sky130_asc_pfet_01v8_lvt_60_0/GATE.n28 VSS 0.39fF $ **FLOATING
C2905 sky130_asc_pfet_01v8_lvt_60_0/GATE.n29 VSS 0.08fF $ **FLOATING
C2906 sky130_asc_pfet_01v8_lvt_60_0/GATE.t243 VSS 1.44fF
C2907 sky130_asc_pfet_01v8_lvt_60_0/GATE.n30 VSS 0.33fF $ **FLOATING
C2908 sky130_asc_pfet_01v8_lvt_60_0/GATE.n31 VSS 0.05fF $ **FLOATING
C2909 sky130_asc_pfet_01v8_lvt_60_0/GATE.n32 VSS 0.08fF $ **FLOATING
C2910 sky130_asc_pfet_01v8_lvt_60_0/GATE.n33 VSS 0.05fF $ **FLOATING
C2911 sky130_asc_pfet_01v8_lvt_60_0/GATE.n34 VSS 0.08fF $ **FLOATING
C2912 sky130_asc_pfet_01v8_lvt_60_0/GATE.t147 VSS 1.44fF
C2913 sky130_asc_pfet_01v8_lvt_60_0/GATE.n35 VSS 0.33fF $ **FLOATING
C2914 sky130_asc_pfet_01v8_lvt_60_0/GATE.n36 VSS 0.05fF $ **FLOATING
C2915 sky130_asc_pfet_01v8_lvt_60_0/GATE.n37 VSS 0.08fF $ **FLOATING
C2916 sky130_asc_pfet_01v8_lvt_60_0/GATE.t122 VSS 1.44fF
C2917 sky130_asc_pfet_01v8_lvt_60_0/GATE.n38 VSS 0.33fF $ **FLOATING
C2918 sky130_asc_pfet_01v8_lvt_60_0/GATE.n39 VSS 0.05fF $ **FLOATING
C2919 sky130_asc_pfet_01v8_lvt_60_0/GATE.n40 VSS 0.08fF $ **FLOATING
C2920 sky130_asc_pfet_01v8_lvt_60_0/GATE.t103 VSS 1.44fF
C2921 sky130_asc_pfet_01v8_lvt_60_0/GATE.n41 VSS 0.33fF $ **FLOATING
C2922 sky130_asc_pfet_01v8_lvt_60_0/GATE.n42 VSS 0.05fF $ **FLOATING
C2923 sky130_asc_pfet_01v8_lvt_60_0/GATE.n43 VSS 0.08fF $ **FLOATING
C2924 sky130_asc_pfet_01v8_lvt_60_0/GATE.t153 VSS 1.44fF
C2925 sky130_asc_pfet_01v8_lvt_60_0/GATE.n44 VSS 0.33fF $ **FLOATING
C2926 sky130_asc_pfet_01v8_lvt_60_0/GATE.n45 VSS 0.05fF $ **FLOATING
C2927 sky130_asc_pfet_01v8_lvt_60_0/GATE.n46 VSS 0.08fF $ **FLOATING
C2928 sky130_asc_pfet_01v8_lvt_60_0/GATE.t151 VSS 1.44fF
C2929 sky130_asc_pfet_01v8_lvt_60_0/GATE.n47 VSS 0.38fF $ **FLOATING
C2930 sky130_asc_pfet_01v8_lvt_60_0/GATE.n48 VSS 0.08fF $ **FLOATING
C2931 sky130_asc_pfet_01v8_lvt_60_0/GATE.t80 VSS 1.44fF
C2932 sky130_asc_pfet_01v8_lvt_60_0/GATE.n49 VSS 0.39fF $ **FLOATING
C2933 sky130_asc_pfet_01v8_lvt_60_0/GATE.n50 VSS 0.08fF $ **FLOATING
C2934 sky130_asc_pfet_01v8_lvt_60_0/GATE.t141 VSS 1.44fF
C2935 sky130_asc_pfet_01v8_lvt_60_0/GATE.n51 VSS 0.33fF $ **FLOATING
C2936 sky130_asc_pfet_01v8_lvt_60_0/GATE.n52 VSS 0.05fF $ **FLOATING
C2937 sky130_asc_pfet_01v8_lvt_60_0/GATE.n53 VSS 0.08fF $ **FLOATING
C2938 sky130_asc_pfet_01v8_lvt_60_0/GATE.n54 VSS 0.05fF $ **FLOATING
C2939 sky130_asc_pfet_01v8_lvt_60_0/GATE.n55 VSS 0.08fF $ **FLOATING
C2940 sky130_asc_pfet_01v8_lvt_60_0/GATE.t115 VSS 1.44fF
C2941 sky130_asc_pfet_01v8_lvt_60_0/GATE.n56 VSS 0.33fF $ **FLOATING
C2942 sky130_asc_pfet_01v8_lvt_60_0/GATE.n57 VSS 0.05fF $ **FLOATING
C2943 sky130_asc_pfet_01v8_lvt_60_0/GATE.n58 VSS 0.08fF $ **FLOATING
C2944 sky130_asc_pfet_01v8_lvt_60_0/GATE.t213 VSS 1.44fF
C2945 sky130_asc_pfet_01v8_lvt_60_0/GATE.n59 VSS 0.33fF $ **FLOATING
C2946 sky130_asc_pfet_01v8_lvt_60_0/GATE.n60 VSS 0.05fF $ **FLOATING
C2947 sky130_asc_pfet_01v8_lvt_60_0/GATE.n61 VSS 0.08fF $ **FLOATING
C2948 sky130_asc_pfet_01v8_lvt_60_0/GATE.t177 VSS 1.44fF
C2949 sky130_asc_pfet_01v8_lvt_60_0/GATE.n62 VSS 0.33fF $ **FLOATING
C2950 sky130_asc_pfet_01v8_lvt_60_0/GATE.n63 VSS 0.05fF $ **FLOATING
C2951 sky130_asc_pfet_01v8_lvt_60_0/GATE.n64 VSS 0.08fF $ **FLOATING
C2952 sky130_asc_pfet_01v8_lvt_60_0/GATE.t203 VSS 1.44fF
C2953 sky130_asc_pfet_01v8_lvt_60_0/GATE.n65 VSS 0.33fF $ **FLOATING
C2954 sky130_asc_pfet_01v8_lvt_60_0/GATE.n66 VSS 0.05fF $ **FLOATING
C2955 sky130_asc_pfet_01v8_lvt_60_0/GATE.n67 VSS 0.08fF $ **FLOATING
C2956 sky130_asc_pfet_01v8_lvt_60_0/GATE.t167 VSS 1.44fF
C2957 sky130_asc_pfet_01v8_lvt_60_0/GATE.n68 VSS 0.38fF $ **FLOATING
C2958 sky130_asc_pfet_01v8_lvt_60_0/GATE.n69 VSS 0.08fF $ **FLOATING
C2959 sky130_asc_pfet_01v8_lvt_60_0/GATE.t164 VSS 1.44fF
C2960 sky130_asc_pfet_01v8_lvt_60_0/GATE.n70 VSS 0.39fF $ **FLOATING
C2961 sky130_asc_pfet_01v8_lvt_60_0/GATE.n71 VSS 0.08fF $ **FLOATING
C2962 sky130_asc_pfet_01v8_lvt_60_0/GATE.t228 VSS 1.44fF
C2963 sky130_asc_pfet_01v8_lvt_60_0/GATE.n72 VSS 0.38fF $ **FLOATING
C2964 sky130_asc_pfet_01v8_lvt_60_0/GATE.n73 VSS 0.08fF $ **FLOATING
C2965 sky130_asc_pfet_01v8_lvt_60_0/GATE.n74 VSS 0.05fF $ **FLOATING
C2966 sky130_asc_pfet_01v8_lvt_60_0/GATE.n75 VSS 0.08fF $ **FLOATING
C2967 sky130_asc_pfet_01v8_lvt_60_0/GATE.n76 VSS 0.08fF $ **FLOATING
C2968 sky130_asc_pfet_01v8_lvt_60_0/GATE.t240 VSS 1.44fF
C2969 sky130_asc_pfet_01v8_lvt_60_0/GATE.n77 VSS 0.38fF $ **FLOATING
C2970 sky130_asc_pfet_01v8_lvt_60_0/GATE.t238 VSS 1.44fF
C2971 sky130_asc_pfet_01v8_lvt_60_0/GATE.n78 VSS 0.39fF $ **FLOATING
C2972 sky130_asc_pfet_01v8_lvt_60_0/GATE.t235 VSS 1.44fF
C2973 sky130_asc_pfet_01v8_lvt_60_0/GATE.n79 VSS 0.38fF $ **FLOATING
C2974 sky130_asc_pfet_01v8_lvt_60_0/GATE.t137 VSS 1.44fF
C2975 sky130_asc_pfet_01v8_lvt_60_0/GATE.n80 VSS 0.39fF $ **FLOATING
C2976 sky130_asc_pfet_01v8_lvt_60_0/GATE.t211 VSS 1.44fF
C2977 sky130_asc_pfet_01v8_lvt_60_0/GATE.n81 VSS 0.38fF $ **FLOATING
C2978 sky130_asc_pfet_01v8_lvt_60_0/GATE.t222 VSS 1.44fF
C2979 sky130_asc_pfet_01v8_lvt_60_0/GATE.n82 VSS 0.39fF $ **FLOATING
C2980 sky130_asc_pfet_01v8_lvt_60_0/GATE.t69 VSS 1.44fF
C2981 sky130_asc_pfet_01v8_lvt_60_0/GATE.n83 VSS 0.38fF $ **FLOATING
C2982 sky130_asc_pfet_01v8_lvt_12_1/GATE VSS 0.03fF $ **FLOATING
C2983 sky130_asc_pfet_01v8_lvt_60_0/GATE.t202 VSS 1.44fF
C2984 sky130_asc_pfet_01v8_lvt_60_0/GATE.n84 VSS 0.39fF $ **FLOATING
C2985 sky130_asc_pfet_01v8_lvt_60_0/GATE.n85 VSS 0.06fF $ **FLOATING
C2986 sky130_asc_pfet_01v8_lvt_60_0/GATE.n86 VSS 0.05fF $ **FLOATING
C2987 sky130_asc_pfet_01v8_lvt_60_0/GATE.n87 VSS 0.08fF $ **FLOATING
C2988 sky130_asc_pfet_01v8_lvt_60_0/GATE.t30 VSS 1.44fF
C2989 sky130_asc_pfet_01v8_lvt_60_0/GATE.n88 VSS 0.33fF $ **FLOATING
C2990 sky130_asc_pfet_01v8_lvt_60_0/GATE.n89 VSS 0.05fF $ **FLOATING
C2991 sky130_asc_pfet_01v8_lvt_60_0/GATE.n90 VSS 0.08fF $ **FLOATING
C2992 sky130_asc_pfet_01v8_lvt_60_0/GATE.t28 VSS 1.44fF
C2993 sky130_asc_pfet_01v8_lvt_60_0/GATE.n91 VSS 0.33fF $ **FLOATING
C2994 sky130_asc_pfet_01v8_lvt_60_0/GATE.n92 VSS 0.05fF $ **FLOATING
C2995 sky130_asc_pfet_01v8_lvt_60_0/GATE.n93 VSS 0.08fF $ **FLOATING
C2996 sky130_asc_pfet_01v8_lvt_60_0/GATE.t226 VSS 1.44fF
C2997 sky130_asc_pfet_01v8_lvt_60_0/GATE.n94 VSS 0.33fF $ **FLOATING
C2998 sky130_asc_pfet_01v8_lvt_60_0/GATE.n95 VSS 0.05fF $ **FLOATING
C2999 sky130_asc_pfet_01v8_lvt_60_0/GATE.n96 VSS 0.08fF $ **FLOATING
C3000 sky130_asc_pfet_01v8_lvt_60_0/GATE.t241 VSS 1.44fF
C3001 sky130_asc_pfet_01v8_lvt_60_0/GATE.n97 VSS 0.33fF $ **FLOATING
C3002 sky130_asc_pfet_01v8_lvt_60_0/GATE.n98 VSS 0.05fF $ **FLOATING
C3003 sky130_asc_pfet_01v8_lvt_60_0/GATE.n99 VSS 0.07fF $ **FLOATING
C3004 sky130_asc_pfet_01v8_lvt_60_0/GATE.n100 VSS 0.04fF $ **FLOATING
C3005 sky130_asc_pfet_01v8_lvt_60_0/GATE.t64 VSS 1.44fF
C3006 sky130_asc_pfet_01v8_lvt_60_0/GATE.n101 VSS 0.39fF $ **FLOATING
C3007 sky130_asc_nfet_01v8_lvt_9_0/DRAIN VSS 0.05fF $ **FLOATING
C3008 sky130_asc_pfet_01v8_lvt_60_0/GATE.t8 VSS 0.04fF
C3009 sky130_asc_pfet_01v8_lvt_60_0/GATE.t23 VSS 0.04fF
C3010 sky130_asc_pfet_01v8_lvt_60_0/GATE.n102 VSS 0.27fF $ **FLOATING
C3011 sky130_asc_pfet_01v8_lvt_60_0/GATE.t1 VSS 0.04fF
C3012 sky130_asc_pfet_01v8_lvt_60_0/GATE.t3 VSS 0.04fF
C3013 sky130_asc_pfet_01v8_lvt_60_0/GATE.n103 VSS 0.27fF $ **FLOATING
C3014 sky130_asc_pfet_01v8_lvt_60_0/GATE.t4 VSS 0.04fF
C3015 sky130_asc_pfet_01v8_lvt_60_0/GATE.t2 VSS 0.04fF
C3016 sky130_asc_pfet_01v8_lvt_60_0/GATE.n104 VSS 0.27fF $ **FLOATING
C3017 sky130_asc_pfet_01v8_lvt_60_0/GATE.t5 VSS 0.42fF
C3018 sky130_asc_pfet_01v8_lvt_60_0/GATE.n105 VSS 0.21fF $ **FLOATING
C3019 sky130_asc_pfet_01v8_lvt_60_0/GATE.n106 VSS 0.18fF $ **FLOATING
C3020 sky130_asc_pfet_01v8_lvt_60_0/GATE.n107 VSS 0.18fF $ **FLOATING
C3021 sky130_asc_pfet_01v8_lvt_60_0/GATE.n108 VSS 0.13fF $ **FLOATING
C3022 sky130_asc_pfet_01v8_lvt_60_0/GATE.n109 VSS 0.00fF $ **FLOATING
C3023 sky130_asc_pfet_01v8_lvt_60_0/GATE.n110 VSS 0.01fF $ **FLOATING
C3024 sky130_asc_pfet_01v8_lvt_60_0/GATE.n111 VSS 0.00fF $ **FLOATING
C3025 sky130_asc_pfet_01v8_lvt_60_0/GATE.n112 VSS 0.00fF $ **FLOATING
C3026 sky130_asc_pfet_01v8_lvt_60_0/GATE.n113 VSS 0.00fF $ **FLOATING
C3027 sky130_asc_pfet_01v8_lvt_60_0/GATE.n114 VSS 0.00fF $ **FLOATING
C3028 sky130_asc_pfet_01v8_lvt_60_0/GATE.n115 VSS 0.00fF $ **FLOATING
C3029 sky130_asc_pfet_01v8_lvt_60_0/GATE.n116 VSS 0.00fF $ **FLOATING
C3030 sky130_asc_pfet_01v8_lvt_60_0/GATE.n117 VSS 0.00fF $ **FLOATING
C3031 sky130_asc_pfet_01v8_lvt_60_0/GATE.n118 VSS 0.00fF $ **FLOATING
C3032 sky130_asc_pfet_01v8_lvt_60_0/GATE.n119 VSS 0.00fF $ **FLOATING
C3033 sky130_asc_pfet_01v8_lvt_60_0/GATE.n120 VSS 0.00fF $ **FLOATING
C3034 sky130_asc_pfet_01v8_lvt_60_0/GATE.n121 VSS 0.00fF $ **FLOATING
C3035 sky130_asc_pfet_01v8_lvt_60_0/GATE.n122 VSS 0.00fF $ **FLOATING
C3036 sky130_asc_pfet_01v8_lvt_60_0/GATE.n123 VSS 0.00fF $ **FLOATING
C3037 sky130_asc_pfet_01v8_lvt_60_0/GATE.n124 VSS 0.00fF $ **FLOATING
C3038 sky130_asc_pfet_01v8_lvt_60_0/GATE.n125 VSS 0.00fF $ **FLOATING
C3039 sky130_asc_pfet_01v8_lvt_60_0/GATE.n126 VSS 0.00fF $ **FLOATING
C3040 sky130_asc_pfet_01v8_lvt_60_0/GATE.n127 VSS 0.00fF $ **FLOATING
C3041 sky130_asc_pfet_01v8_lvt_60_0/GATE.n128 VSS 0.01fF $ **FLOATING
C3042 sky130_asc_pfet_01v8_lvt_60_0/GATE.n129 VSS 0.00fF $ **FLOATING
C3043 sky130_asc_pfet_01v8_lvt_60_0/GATE.n130 VSS 0.00fF $ **FLOATING
C3044 sky130_asc_pfet_01v8_lvt_60_0/GATE.n131 VSS 0.00fF $ **FLOATING
C3045 sky130_asc_pfet_01v8_lvt_60_0/GATE.n132 VSS 0.00fF $ **FLOATING
C3046 sky130_asc_pfet_01v8_lvt_60_0/GATE.n133 VSS 0.00fF $ **FLOATING
C3047 sky130_asc_pfet_01v8_lvt_60_0/GATE.n134 VSS 0.00fF $ **FLOATING
C3048 sky130_asc_pfet_01v8_lvt_60_0/GATE.n135 VSS 0.00fF $ **FLOATING
C3049 sky130_asc_pfet_01v8_lvt_60_0/GATE.n136 VSS 0.00fF $ **FLOATING
C3050 sky130_asc_pfet_01v8_lvt_60_0/GATE.n137 VSS 0.00fF $ **FLOATING
C3051 sky130_asc_pfet_01v8_lvt_60_0/GATE.n138 VSS 0.00fF $ **FLOATING
C3052 sky130_asc_pfet_01v8_lvt_60_0/GATE.n139 VSS 0.00fF $ **FLOATING
C3053 sky130_asc_pfet_01v8_lvt_60_0/GATE.n140 VSS 0.00fF $ **FLOATING
C3054 sky130_asc_pfet_01v8_lvt_60_0/GATE.n141 VSS 0.00fF $ **FLOATING
C3055 sky130_asc_pfet_01v8_lvt_60_0/GATE.n142 VSS 0.00fF $ **FLOATING
C3056 sky130_asc_pfet_01v8_lvt_60_0/GATE.n143 VSS 0.00fF $ **FLOATING
C3057 sky130_asc_pfet_01v8_lvt_60_0/GATE.t0 VSS 0.04fF
C3058 sky130_asc_pfet_01v8_lvt_60_0/GATE.t22 VSS 0.04fF
C3059 sky130_asc_pfet_01v8_lvt_60_0/GATE.n144 VSS 0.07fF $ **FLOATING
C3060 sky130_asc_pfet_01v8_lvt_60_0/GATE.n145 VSS 0.01fF $ **FLOATING
C3061 sky130_asc_pfet_01v8_lvt_60_0/GATE.t45 VSS 1.44fF
C3062 sky130_asc_pfet_01v8_lvt_60_0/GATE.n146 VSS 0.38fF $ **FLOATING
C3063 sky130_asc_pfet_01v8_lvt_60_0/GATE.n147 VSS 0.30fF $ **FLOATING
C3064 sky130_asc_pfet_01v8_lvt_60_0/GATE.n148 VSS 0.05fF $ **FLOATING
C3065 sky130_asc_pfet_01v8_lvt_60_0/GATE.n149 VSS 0.08fF $ **FLOATING
C3066 sky130_asc_pfet_01v8_lvt_60_0/GATE.t234 VSS 1.44fF
C3067 sky130_asc_pfet_01v8_lvt_60_0/GATE.n150 VSS 0.33fF $ **FLOATING
C3068 sky130_asc_pfet_01v8_lvt_60_0/GATE.n151 VSS 0.05fF $ **FLOATING
C3069 sky130_asc_pfet_01v8_lvt_60_0/GATE.n152 VSS 0.08fF $ **FLOATING
C3070 sky130_asc_pfet_01v8_lvt_60_0/GATE.t37 VSS 1.44fF
C3071 sky130_asc_pfet_01v8_lvt_60_0/GATE.n153 VSS 0.33fF $ **FLOATING
C3072 sky130_asc_pfet_01v8_lvt_60_0/GATE.n154 VSS 0.05fF $ **FLOATING
C3073 sky130_asc_pfet_01v8_lvt_60_0/GATE.n155 VSS 0.08fF $ **FLOATING
C3074 sky130_asc_pfet_01v8_lvt_60_0/GATE.t87 VSS 1.44fF
C3075 sky130_asc_pfet_01v8_lvt_60_0/GATE.n156 VSS 0.33fF $ **FLOATING
C3076 sky130_asc_pfet_01v8_lvt_60_0/GATE.n157 VSS 0.05fF $ **FLOATING
C3077 sky130_asc_pfet_01v8_lvt_60_0/GATE.n158 VSS 0.08fF $ **FLOATING
C3078 sky130_asc_pfet_01v8_lvt_60_0/GATE.t47 VSS 1.44fF
C3079 sky130_asc_pfet_01v8_lvt_60_0/GATE.n159 VSS 0.33fF $ **FLOATING
C3080 sky130_asc_pfet_01v8_lvt_60_0/GATE.n160 VSS 0.05fF $ **FLOATING
C3081 sky130_asc_pfet_01v8_lvt_60_0/GATE.n161 VSS 0.08fF $ **FLOATING
C3082 sky130_asc_pfet_01v8_lvt_60_0/GATE.n162 VSS 0.08fF $ **FLOATING
C3083 sky130_asc_pfet_01v8_lvt_60_0/GATE.n163 VSS 0.04fF $ **FLOATING
C3084 sky130_asc_pfet_01v8_lvt_60_0/GATE.n164 VSS 0.00fF $ **FLOATING
C3085 sky130_asc_pfet_01v8_lvt_60_0/GATE.t219 VSS 1.44fF
C3086 sky130_asc_pfet_01v8_lvt_60_0/GATE.n165 VSS 0.12fF $ **FLOATING
C3087 sky130_asc_pfet_01v8_lvt_60_0/GATE.n166 VSS 0.26fF $ **FLOATING
C3088 sky130_asc_pfet_01v8_lvt_60_0/GATE.n167 VSS 0.00fF $ **FLOATING
C3089 sky130_asc_pfet_01v8_lvt_60_0/GATE.n168 VSS 0.18fF $ **FLOATING
C3090 sky130_asc_pfet_01v8_lvt_60_0/GATE.t231 VSS 1.44fF
C3091 sky130_asc_pfet_01v8_lvt_60_0/GATE.n169 VSS 0.38fF $ **FLOATING
C3092 sky130_asc_pfet_01v8_lvt_60_0/GATE.t78 VSS 1.44fF
C3093 sky130_asc_pfet_01v8_lvt_60_0/GATE.n170 VSS 0.38fF $ **FLOATING
C3094 sky130_asc_pfet_01v8_lvt_60_0/GATE.t56 VSS 1.44fF
C3095 sky130_asc_pfet_01v8_lvt_60_0/GATE.n171 VSS 0.38fF $ **FLOATING
C3096 sky130_asc_pfet_01v8_lvt_60_0/GATE.t32 VSS 1.44fF
C3097 sky130_asc_pfet_01v8_lvt_60_0/GATE.n172 VSS 0.39fF $ **FLOATING
C3098 sky130_asc_pfet_01v8_lvt_60_0/GATE.t107 VSS 1.55fF
C3099 sky130_asc_pfet_01v8_lvt_60_0/GATE.n173 VSS 0.44fF $ **FLOATING
C3100 sky130_asc_pfet_01v8_lvt_60_0/GATE.t67 VSS 1.44fF
C3101 sky130_asc_pfet_01v8_lvt_60_0/GATE.n174 VSS 0.34fF $ **FLOATING
C3102 sky130_asc_pfet_01v8_lvt_60_0/GATE.n175 VSS 0.05fF $ **FLOATING
C3103 sky130_asc_pfet_01v8_lvt_60_0/GATE.n176 VSS 0.11fF $ **FLOATING
C3104 sky130_asc_pfet_01v8_lvt_60_0/GATE.t68 VSS 1.44fF
C3105 sky130_asc_pfet_01v8_lvt_60_0/GATE.n177 VSS 0.33fF $ **FLOATING
C3106 sky130_asc_pfet_01v8_lvt_60_0/GATE.n178 VSS 0.05fF $ **FLOATING
C3107 sky130_asc_pfet_01v8_lvt_60_0/GATE.n179 VSS 0.08fF $ **FLOATING
C3108 sky130_asc_pfet_01v8_lvt_60_0/GATE.t244 VSS 1.44fF
C3109 sky130_asc_pfet_01v8_lvt_60_0/GATE.n180 VSS 0.33fF $ **FLOATING
C3110 sky130_asc_pfet_01v8_lvt_60_0/GATE.n181 VSS 0.05fF $ **FLOATING
C3111 sky130_asc_pfet_01v8_lvt_60_0/GATE.n182 VSS 0.08fF $ **FLOATING
C3112 sky130_asc_pfet_01v8_lvt_60_0/GATE.t95 VSS 1.44fF
C3113 sky130_asc_pfet_01v8_lvt_60_0/GATE.n183 VSS 0.33fF $ **FLOATING
C3114 sky130_asc_pfet_01v8_lvt_60_0/GATE.n184 VSS 0.05fF $ **FLOATING
C3115 sky130_asc_pfet_01v8_lvt_60_0/GATE.n185 VSS 0.08fF $ **FLOATING
C3116 sky130_asc_pfet_01v8_lvt_60_0/GATE.n186 VSS 0.08fF $ **FLOATING
C3117 sky130_asc_pfet_01v8_lvt_60_0/GATE.n187 VSS 0.08fF $ **FLOATING
C3118 sky130_asc_pfet_01v8_lvt_60_0/GATE.t57 VSS 1.44fF
C3119 sky130_asc_pfet_01v8_lvt_60_0/GATE.n188 VSS 0.33fF $ **FLOATING
C3120 sky130_asc_pfet_01v8_lvt_60_0/GATE.n189 VSS 0.05fF $ **FLOATING
C3121 sky130_asc_pfet_01v8_lvt_60_0/GATE.n190 VSS 0.08fF $ **FLOATING
C3122 sky130_asc_pfet_01v8_lvt_60_0/GATE.n191 VSS 0.05fF $ **FLOATING
C3123 sky130_asc_pfet_01v8_lvt_60_0/GATE.n192 VSS 0.08fF $ **FLOATING
C3124 sky130_asc_pfet_01v8_lvt_60_0/GATE.t230 VSS 1.44fF
C3125 sky130_asc_pfet_01v8_lvt_60_0/GATE.n193 VSS 0.33fF $ **FLOATING
C3126 sky130_asc_pfet_01v8_lvt_60_0/GATE.n194 VSS 0.05fF $ **FLOATING
C3127 sky130_asc_pfet_01v8_lvt_60_0/GATE.n195 VSS 0.08fF $ **FLOATING
C3128 sky130_asc_pfet_01v8_lvt_60_0/GATE.t96 VSS 1.44fF
C3129 sky130_asc_pfet_01v8_lvt_60_0/GATE.n196 VSS 0.33fF $ **FLOATING
C3130 sky130_asc_pfet_01v8_lvt_60_0/GATE.n197 VSS 0.05fF $ **FLOATING
C3131 sky130_asc_pfet_01v8_lvt_60_0/GATE.n198 VSS 0.08fF $ **FLOATING
C3132 sky130_asc_pfet_01v8_lvt_60_0/GATE.t58 VSS 1.44fF
C3133 sky130_asc_pfet_01v8_lvt_60_0/GATE.n199 VSS 0.33fF $ **FLOATING
C3134 sky130_asc_pfet_01v8_lvt_60_0/GATE.n200 VSS 0.05fF $ **FLOATING
C3135 sky130_asc_pfet_01v8_lvt_60_0/GATE.n201 VSS 0.08fF $ **FLOATING
C3136 sky130_asc_pfet_01v8_lvt_60_0/GATE.t59 VSS 1.44fF
C3137 sky130_asc_pfet_01v8_lvt_60_0/GATE.n202 VSS 0.33fF $ **FLOATING
C3138 sky130_asc_pfet_01v8_lvt_60_0/GATE.n203 VSS 0.05fF $ **FLOATING
C3139 sky130_asc_pfet_01v8_lvt_60_0/GATE.n204 VSS 0.08fF $ **FLOATING
C3140 sky130_asc_pfet_01v8_lvt_60_0/GATE.n205 VSS 0.08fF $ **FLOATING
C3141 sky130_asc_pfet_01v8_lvt_60_0/GATE.n206 VSS 0.07fF $ **FLOATING
C3142 sky130_asc_pfet_01v8_lvt_60_0/GATE.n207 VSS 0.22fF $ **FLOATING
C3143 sky130_asc_pfet_01v8_lvt_60_0/GATE.t84 VSS 1.44fF
C3144 sky130_asc_pfet_01v8_lvt_60_0/GATE.n208 VSS 0.33fF $ **FLOATING
C3145 sky130_asc_pfet_01v8_lvt_60_0/GATE.n209 VSS 0.05fF $ **FLOATING
C3146 sky130_asc_pfet_01v8_lvt_60_0/GATE.n210 VSS 0.04fF $ **FLOATING
C3147 sky130_asc_pfet_01v8_lvt_60_0/GATE.n211 VSS 0.05fF $ **FLOATING
C3148 sky130_asc_pfet_01v8_lvt_60_0/GATE.n212 VSS 0.08fF $ **FLOATING
C3149 sky130_asc_pfet_01v8_lvt_60_0/GATE.t41 VSS 1.44fF
C3150 sky130_asc_pfet_01v8_lvt_60_0/GATE.n213 VSS 0.33fF $ **FLOATING
C3151 sky130_asc_pfet_01v8_lvt_60_0/GATE.n214 VSS 0.05fF $ **FLOATING
C3152 sky130_asc_pfet_01v8_lvt_60_0/GATE.n215 VSS 0.08fF $ **FLOATING
C3153 sky130_asc_pfet_01v8_lvt_60_0/GATE.n216 VSS 0.08fF $ **FLOATING
C3154 sky130_asc_pfet_01v8_lvt_60_1/GATE VSS 0.03fF $ **FLOATING
C3155 sky130_asc_pfet_01v8_lvt_60_0/GATE.n217 VSS 0.09fF $ **FLOATING
C3156 sky130_asc_pfet_01v8_lvt_60_0/GATE.t77 VSS 1.44fF
C3157 sky130_asc_pfet_01v8_lvt_60_0/GATE.n218 VSS 0.37fF $ **FLOATING
C3158 sky130_asc_pfet_01v8_lvt_60_0/GATE.n219 VSS 0.05fF $ **FLOATING
C3159 sky130_asc_pfet_01v8_lvt_60_0/GATE.n220 VSS 0.08fF $ **FLOATING
C3160 sky130_asc_pfet_01v8_lvt_60_0/GATE.t140 VSS 1.44fF
C3161 sky130_asc_pfet_01v8_lvt_60_0/GATE.n221 VSS 0.33fF $ **FLOATING
C3162 sky130_asc_pfet_01v8_lvt_60_0/GATE.n222 VSS 0.05fF $ **FLOATING
C3163 sky130_asc_pfet_01v8_lvt_60_0/GATE.n223 VSS 0.08fF $ **FLOATING
C3164 sky130_asc_pfet_01v8_lvt_60_0/GATE.t113 VSS 1.44fF
C3165 sky130_asc_pfet_01v8_lvt_60_0/GATE.n224 VSS 0.33fF $ **FLOATING
C3166 sky130_asc_pfet_01v8_lvt_60_0/GATE.n225 VSS 0.05fF $ **FLOATING
C3167 sky130_asc_pfet_01v8_lvt_60_0/GATE.n226 VSS 0.08fF $ **FLOATING
C3168 sky130_asc_pfet_01v8_lvt_60_0/GATE.t35 VSS 1.44fF
C3169 sky130_asc_pfet_01v8_lvt_60_0/GATE.n227 VSS 0.38fF $ **FLOATING
C3170 sky130_asc_pfet_01v8_lvt_60_0/GATE.n228 VSS 0.08fF $ **FLOATING
C3171 sky130_asc_pfet_01v8_lvt_60_0/GATE.t31 VSS 1.44fF
C3172 sky130_asc_pfet_01v8_lvt_60_0/GATE.n229 VSS 0.39fF $ **FLOATING
C3173 sky130_asc_pfet_01v8_lvt_60_0/GATE.n230 VSS 0.08fF $ **FLOATING
C3174 sky130_asc_pfet_01v8_lvt_60_0/GATE.t29 VSS 1.44fF
C3175 sky130_asc_pfet_01v8_lvt_60_0/GATE.n231 VSS 0.33fF $ **FLOATING
C3176 sky130_asc_pfet_01v8_lvt_60_0/GATE.n232 VSS 0.05fF $ **FLOATING
C3177 sky130_asc_pfet_01v8_lvt_60_0/GATE.n233 VSS 0.08fF $ **FLOATING
C3178 sky130_asc_pfet_01v8_lvt_60_0/GATE.n234 VSS 0.05fF $ **FLOATING
C3179 sky130_asc_pfet_01v8_lvt_60_0/GATE.n235 VSS 0.08fF $ **FLOATING
C3180 sky130_asc_pfet_01v8_lvt_60_0/GATE.t74 VSS 1.44fF
C3181 sky130_asc_pfet_01v8_lvt_60_0/GATE.n236 VSS 0.33fF $ **FLOATING
C3182 sky130_asc_pfet_01v8_lvt_60_0/GATE.n237 VSS 0.05fF $ **FLOATING
C3183 sky130_asc_pfet_01v8_lvt_60_0/GATE.n238 VSS 0.08fF $ **FLOATING
C3184 sky130_asc_pfet_01v8_lvt_60_0/GATE.t53 VSS 1.44fF
C3185 sky130_asc_pfet_01v8_lvt_60_0/GATE.n239 VSS 0.33fF $ **FLOATING
C3186 sky130_asc_pfet_01v8_lvt_60_0/GATE.n240 VSS 0.05fF $ **FLOATING
C3187 sky130_asc_pfet_01v8_lvt_60_0/GATE.n241 VSS 0.08fF $ **FLOATING
C3188 sky130_asc_pfet_01v8_lvt_60_0/GATE.t52 VSS 1.44fF
C3189 sky130_asc_pfet_01v8_lvt_60_0/GATE.n242 VSS 0.33fF $ **FLOATING
C3190 sky130_asc_pfet_01v8_lvt_60_0/GATE.n243 VSS 0.05fF $ **FLOATING
C3191 sky130_asc_pfet_01v8_lvt_60_0/GATE.n244 VSS 0.08fF $ **FLOATING
C3192 sky130_asc_pfet_01v8_lvt_60_0/GATE.t49 VSS 1.44fF
C3193 sky130_asc_pfet_01v8_lvt_60_0/GATE.n245 VSS 0.33fF $ **FLOATING
C3194 sky130_asc_pfet_01v8_lvt_60_0/GATE.n246 VSS 0.05fF $ **FLOATING
C3195 sky130_asc_pfet_01v8_lvt_60_0/GATE.n247 VSS 0.08fF $ **FLOATING
C3196 sky130_asc_pfet_01v8_lvt_60_0/GATE.t48 VSS 1.44fF
C3197 sky130_asc_pfet_01v8_lvt_60_0/GATE.n248 VSS 0.38fF $ **FLOATING
C3198 sky130_asc_pfet_01v8_lvt_60_0/GATE.n249 VSS 0.08fF $ **FLOATING
C3199 sky130_asc_pfet_01v8_lvt_60_0/GATE.t88 VSS 1.44fF
C3200 sky130_asc_pfet_01v8_lvt_60_0/GATE.n250 VSS 0.39fF $ **FLOATING
C3201 sky130_asc_pfet_01v8_lvt_60_0/GATE.n251 VSS 0.08fF $ **FLOATING
C3202 sky130_asc_pfet_01v8_lvt_60_0/GATE.t86 VSS 1.44fF
C3203 sky130_asc_pfet_01v8_lvt_60_0/GATE.n252 VSS 0.33fF $ **FLOATING
C3204 sky130_asc_pfet_01v8_lvt_60_0/GATE.n253 VSS 0.05fF $ **FLOATING
C3205 sky130_asc_pfet_01v8_lvt_60_0/GATE.n254 VSS 0.08fF $ **FLOATING
C3206 sky130_asc_pfet_01v8_lvt_60_0/GATE.n255 VSS 0.05fF $ **FLOATING
C3207 sky130_asc_pfet_01v8_lvt_60_0/GATE.n256 VSS 0.08fF $ **FLOATING
C3208 sky130_asc_pfet_01v8_lvt_60_0/GATE.t125 VSS 1.44fF
C3209 sky130_asc_pfet_01v8_lvt_60_0/GATE.n257 VSS 0.33fF $ **FLOATING
C3210 sky130_asc_pfet_01v8_lvt_60_0/GATE.n258 VSS 0.05fF $ **FLOATING
C3211 sky130_asc_pfet_01v8_lvt_60_0/GATE.n259 VSS 0.08fF $ **FLOATING
C3212 sky130_asc_pfet_01v8_lvt_60_0/GATE.t82 VSS 1.44fF
C3213 sky130_asc_pfet_01v8_lvt_60_0/GATE.n260 VSS 0.33fF $ **FLOATING
C3214 sky130_asc_pfet_01v8_lvt_60_0/GATE.n261 VSS 0.05fF $ **FLOATING
C3215 sky130_asc_pfet_01v8_lvt_60_0/GATE.n262 VSS 0.08fF $ **FLOATING
C3216 sky130_asc_pfet_01v8_lvt_60_0/GATE.t61 VSS 1.44fF
C3217 sky130_asc_pfet_01v8_lvt_60_0/GATE.n263 VSS 0.33fF $ **FLOATING
C3218 sky130_asc_pfet_01v8_lvt_60_0/GATE.n264 VSS 0.05fF $ **FLOATING
C3219 sky130_asc_pfet_01v8_lvt_60_0/GATE.n265 VSS 0.08fF $ **FLOATING
C3220 sky130_asc_pfet_01v8_lvt_60_0/GATE.t118 VSS 1.44fF
C3221 sky130_asc_pfet_01v8_lvt_60_0/GATE.n266 VSS 0.33fF $ **FLOATING
C3222 sky130_asc_pfet_01v8_lvt_60_0/GATE.n267 VSS 0.05fF $ **FLOATING
C3223 sky130_asc_pfet_01v8_lvt_60_0/GATE.n268 VSS 0.08fF $ **FLOATING
C3224 sky130_asc_pfet_01v8_lvt_60_0/GATE.t98 VSS 1.44fF
C3225 sky130_asc_pfet_01v8_lvt_60_0/GATE.n269 VSS 0.38fF $ **FLOATING
C3226 sky130_asc_pfet_01v8_lvt_60_0/GATE.n270 VSS 0.08fF $ **FLOATING
C3227 sky130_asc_pfet_01v8_lvt_60_0/GATE.t143 VSS 1.44fF
C3228 sky130_asc_pfet_01v8_lvt_60_0/GATE.n271 VSS 0.39fF $ **FLOATING
C3229 sky130_asc_pfet_01v8_lvt_60_0/GATE.n272 VSS 0.08fF $ **FLOATING
C3230 sky130_asc_pfet_01v8_lvt_60_0/GATE.t94 VSS 1.44fF
C3231 sky130_asc_pfet_01v8_lvt_60_0/GATE.n273 VSS 0.38fF $ **FLOATING
C3232 sky130_asc_pfet_01v8_lvt_60_0/GATE.n274 VSS 0.08fF $ **FLOATING
C3233 sky130_asc_pfet_01v8_lvt_60_0/GATE.n275 VSS 0.05fF $ **FLOATING
C3234 sky130_asc_pfet_01v8_lvt_60_0/GATE.n276 VSS 0.08fF $ **FLOATING
C3235 sky130_asc_pfet_01v8_lvt_60_0/GATE.t136 VSS 1.44fF
C3236 sky130_asc_pfet_01v8_lvt_60_0/GATE.n277 VSS 0.33fF $ **FLOATING
C3237 sky130_asc_pfet_01v8_lvt_60_0/GATE.n278 VSS 0.05fF $ **FLOATING
C3238 sky130_asc_pfet_01v8_lvt_60_0/GATE.n279 VSS 0.08fF $ **FLOATING
C3239 sky130_asc_pfet_01v8_lvt_60_0/GATE.t134 VSS 1.44fF
C3240 sky130_asc_pfet_01v8_lvt_60_0/GATE.n280 VSS 0.33fF $ **FLOATING
C3241 sky130_asc_pfet_01v8_lvt_60_0/GATE.n281 VSS 0.05fF $ **FLOATING
C3242 sky130_asc_pfet_01v8_lvt_60_0/GATE.n282 VSS 0.08fF $ **FLOATING
C3243 sky130_asc_pfet_01v8_lvt_60_0/GATE.t110 VSS 1.44fF
C3244 sky130_asc_pfet_01v8_lvt_60_0/GATE.n283 VSS 0.33fF $ **FLOATING
C3245 sky130_asc_pfet_01v8_lvt_60_0/GATE.n284 VSS 0.05fF $ **FLOATING
C3246 sky130_asc_pfet_01v8_lvt_60_0/GATE.n285 VSS 0.08fF $ **FLOATING
C3247 sky130_asc_pfet_01v8_lvt_60_0/GATE.t205 VSS 1.44fF
C3248 sky130_asc_pfet_01v8_lvt_60_0/GATE.n286 VSS 0.33fF $ **FLOATING
C3249 sky130_asc_pfet_01v8_lvt_60_0/GATE.n287 VSS 0.05fF $ **FLOATING
C3250 sky130_asc_pfet_01v8_lvt_60_0/GATE.n288 VSS 0.08fF $ **FLOATING
C3251 sky130_asc_pfet_01v8_lvt_60_0/GATE.t105 VSS 1.44fF
C3252 sky130_asc_pfet_01v8_lvt_60_0/GATE.n289 VSS 0.38fF $ **FLOATING
C3253 sky130_asc_pfet_01v8_lvt_60_0/GATE.n290 VSS 0.08fF $ **FLOATING
C3254 sky130_asc_pfet_01v8_lvt_60_0/GATE.t91 VSS 1.44fF
C3255 sky130_asc_pfet_01v8_lvt_60_0/GATE.n291 VSS 0.39fF $ **FLOATING
C3256 sky130_asc_pfet_01v8_lvt_60_0/GATE.n292 VSS 0.08fF $ **FLOATING
C3257 sky130_asc_pfet_01v8_lvt_60_0/GATE.t71 VSS 1.44fF
C3258 sky130_asc_pfet_01v8_lvt_60_0/GATE.n293 VSS 0.38fF $ **FLOATING
C3259 sky130_asc_pfet_01v8_lvt_60_0/GATE.n294 VSS 0.08fF $ **FLOATING
C3260 sky130_asc_pfet_01v8_lvt_60_0/GATE.t70 VSS 1.44fF
C3261 sky130_asc_pfet_01v8_lvt_60_0/GATE.n295 VSS 0.33fF $ **FLOATING
C3262 sky130_asc_pfet_01v8_lvt_60_0/GATE.n296 VSS 0.05fF $ **FLOATING
C3263 sky130_asc_pfet_01v8_lvt_60_0/GATE.n297 VSS 0.08fF $ **FLOATING
C3264 sky130_asc_pfet_01v8_lvt_60_0/GATE.n298 VSS 0.05fF $ **FLOATING
C3265 sky130_asc_pfet_01v8_lvt_60_0/GATE.n299 VSS 0.08fF $ **FLOATING
C3266 sky130_asc_pfet_01v8_lvt_60_0/GATE.t108 VSS 1.44fF
C3267 sky130_asc_pfet_01v8_lvt_60_0/GATE.n300 VSS 0.33fF $ **FLOATING
C3268 sky130_asc_pfet_01v8_lvt_60_0/GATE.n301 VSS 0.05fF $ **FLOATING
C3269 sky130_asc_pfet_01v8_lvt_60_0/GATE.n302 VSS 0.08fF $ **FLOATING
C3270 sky130_asc_pfet_01v8_lvt_60_0/GATE.t63 VSS 1.44fF
C3271 sky130_asc_pfet_01v8_lvt_60_0/GATE.n303 VSS 0.33fF $ **FLOATING
C3272 sky130_asc_pfet_01v8_lvt_60_0/GATE.n304 VSS 0.05fF $ **FLOATING
C3273 sky130_asc_pfet_01v8_lvt_60_0/GATE.n305 VSS 0.08fF $ **FLOATING
C3274 sky130_asc_pfet_01v8_lvt_60_0/GATE.t102 VSS 1.44fF
C3275 sky130_asc_pfet_01v8_lvt_60_0/GATE.n306 VSS 0.33fF $ **FLOATING
C3276 sky130_asc_pfet_01v8_lvt_60_0/GATE.n307 VSS 0.05fF $ **FLOATING
C3277 sky130_asc_pfet_01v8_lvt_60_0/GATE.n308 VSS 0.08fF $ **FLOATING
C3278 sky130_asc_pfet_01v8_lvt_60_0/GATE.t85 VSS 1.44fF
C3279 sky130_asc_pfet_01v8_lvt_60_0/GATE.n309 VSS 0.33fF $ **FLOATING
C3280 sky130_asc_pfet_01v8_lvt_60_0/GATE.n310 VSS 0.05fF $ **FLOATING
C3281 sky130_asc_pfet_01v8_lvt_60_0/GATE.n311 VSS 0.08fF $ **FLOATING
C3282 sky130_asc_pfet_01v8_lvt_60_0/GATE.t150 VSS 1.44fF
C3283 sky130_asc_pfet_01v8_lvt_60_0/GATE.n312 VSS 0.39fF $ **FLOATING
C3284 sky130_asc_pfet_01v8_lvt_60_0/GATE.n313 VSS 0.08fF $ **FLOATING
C3285 sky130_asc_pfet_01v8_lvt_60_0/GATE.t121 VSS 1.44fF
C3286 sky130_asc_pfet_01v8_lvt_60_0/GATE.n314 VSS 0.38fF $ **FLOATING
C3287 sky130_asc_pfet_01v8_lvt_60_0/GATE.n315 VSS 0.08fF $ **FLOATING
C3288 sky130_asc_pfet_01v8_lvt_60_0/GATE.t79 VSS 1.44fF
C3289 sky130_asc_pfet_01v8_lvt_60_0/GATE.n316 VSS 0.33fF $ **FLOATING
C3290 sky130_asc_pfet_01v8_lvt_60_0/GATE.n317 VSS 0.05fF $ **FLOATING
C3291 sky130_asc_pfet_01v8_lvt_60_0/GATE.n318 VSS 0.08fF $ **FLOATING
C3292 sky130_asc_pfet_01v8_lvt_60_0/GATE.n319 VSS 0.05fF $ **FLOATING
C3293 sky130_asc_pfet_01v8_lvt_60_0/GATE.n320 VSS 0.08fF $ **FLOATING
C3294 sky130_asc_pfet_01v8_lvt_60_0/GATE.t116 VSS 1.44fF
C3295 sky130_asc_pfet_01v8_lvt_60_0/GATE.n321 VSS 0.33fF $ **FLOATING
C3296 sky130_asc_pfet_01v8_lvt_60_0/GATE.n322 VSS 0.05fF $ **FLOATING
C3297 sky130_asc_pfet_01v8_lvt_60_0/GATE.n323 VSS 0.08fF $ **FLOATING
C3298 sky130_asc_pfet_01v8_lvt_60_0/GATE.t114 VSS 1.44fF
C3299 sky130_asc_pfet_01v8_lvt_60_0/GATE.n324 VSS 0.33fF $ **FLOATING
C3300 sky130_asc_pfet_01v8_lvt_60_0/GATE.n325 VSS 0.05fF $ **FLOATING
C3301 sky130_asc_pfet_01v8_lvt_60_0/GATE.n326 VSS 0.08fF $ **FLOATING
C3302 sky130_asc_pfet_01v8_lvt_60_0/GATE.t178 VSS 1.44fF
C3303 sky130_asc_pfet_01v8_lvt_60_0/GATE.n327 VSS 0.33fF $ **FLOATING
C3304 sky130_asc_pfet_01v8_lvt_60_0/GATE.n328 VSS 0.05fF $ **FLOATING
C3305 sky130_asc_pfet_01v8_lvt_60_0/GATE.n329 VSS 0.08fF $ **FLOATING
C3306 sky130_asc_pfet_01v8_lvt_60_0/GATE.t175 VSS 1.44fF
C3307 sky130_asc_pfet_01v8_lvt_60_0/GATE.n330 VSS 0.33fF $ **FLOATING
C3308 sky130_asc_pfet_01v8_lvt_60_0/GATE.n331 VSS 0.05fF $ **FLOATING
C3309 sky130_asc_pfet_01v8_lvt_60_0/GATE.n332 VSS 0.08fF $ **FLOATING
C3310 sky130_asc_pfet_01v8_lvt_60_0/GATE.t166 VSS 1.44fF
C3311 sky130_asc_pfet_01v8_lvt_60_0/GATE.n333 VSS 0.39fF $ **FLOATING
C3312 sky130_asc_pfet_01v8_lvt_60_0/GATE.n334 VSS 0.08fF $ **FLOATING
C3313 sky130_asc_pfet_01v8_lvt_60_0/GATE.t165 VSS 1.44fF
C3314 sky130_asc_pfet_01v8_lvt_60_0/GATE.n335 VSS 0.38fF $ **FLOATING
C3315 sky130_asc_pfet_01v8_lvt_60_0/GATE.n336 VSS 0.08fF $ **FLOATING
C3316 sky130_asc_pfet_01v8_lvt_60_0/GATE.t129 VSS 1.44fF
C3317 sky130_asc_pfet_01v8_lvt_60_0/GATE.n337 VSS 0.33fF $ **FLOATING
C3318 sky130_asc_pfet_01v8_lvt_60_0/GATE.n338 VSS 0.05fF $ **FLOATING
C3319 sky130_asc_pfet_01v8_lvt_60_0/GATE.n339 VSS 0.08fF $ **FLOATING
C3320 sky130_asc_pfet_01v8_lvt_60_0/GATE.n340 VSS 0.05fF $ **FLOATING
C3321 sky130_asc_pfet_01v8_lvt_60_0/GATE.n341 VSS 0.08fF $ **FLOATING
C3322 sky130_asc_pfet_01v8_lvt_60_0/GATE.t200 VSS 1.44fF
C3323 sky130_asc_pfet_01v8_lvt_60_0/GATE.n342 VSS 0.33fF $ **FLOATING
C3324 sky130_asc_pfet_01v8_lvt_60_0/GATE.n343 VSS 0.05fF $ **FLOATING
C3325 sky130_asc_pfet_01v8_lvt_60_0/GATE.n344 VSS 0.08fF $ **FLOATING
C3326 sky130_asc_pfet_01v8_lvt_60_0/GATE.t198 VSS 1.44fF
C3327 sky130_asc_pfet_01v8_lvt_60_0/GATE.n345 VSS 0.33fF $ **FLOATING
C3328 sky130_asc_pfet_01v8_lvt_60_0/GATE.n346 VSS 0.05fF $ **FLOATING
C3329 sky130_asc_pfet_01v8_lvt_60_0/GATE.n347 VSS 0.08fF $ **FLOATING
C3330 sky130_asc_pfet_01v8_lvt_60_0/GATE.t189 VSS 1.44fF
C3331 sky130_asc_pfet_01v8_lvt_60_0/GATE.n348 VSS 0.33fF $ **FLOATING
C3332 sky130_asc_pfet_01v8_lvt_60_0/GATE.n349 VSS 0.05fF $ **FLOATING
C3333 sky130_asc_pfet_01v8_lvt_60_0/GATE.n350 VSS 0.08fF $ **FLOATING
C3334 sky130_asc_pfet_01v8_lvt_60_0/GATE.t187 VSS 1.44fF
C3335 sky130_asc_pfet_01v8_lvt_60_0/GATE.n351 VSS 0.33fF $ **FLOATING
C3336 sky130_asc_pfet_01v8_lvt_60_0/GATE.n352 VSS 0.05fF $ **FLOATING
C3337 sky130_asc_pfet_01v8_lvt_60_0/GATE.n353 VSS 0.08fF $ **FLOATING
C3338 sky130_asc_pfet_01v8_lvt_60_0/GATE.t152 VSS 1.44fF
C3339 sky130_asc_pfet_01v8_lvt_60_0/GATE.n354 VSS 0.38fF $ **FLOATING
C3340 sky130_asc_pfet_01v8_lvt_60_0/GATE.n355 VSS 0.08fF $ **FLOATING
C3341 sky130_asc_pfet_01v8_lvt_60_0/GATE.t126 VSS 1.44fF
C3342 sky130_asc_pfet_01v8_lvt_60_0/GATE.n356 VSS 0.38fF $ **FLOATING
C3343 sky130_asc_pfet_01v8_lvt_60_0/GATE.n357 VSS 0.08fF $ **FLOATING
C3344 sky130_asc_pfet_01v8_lvt_60_0/GATE.t104 VSS 1.44fF
C3345 sky130_asc_pfet_01v8_lvt_60_0/GATE.n358 VSS 0.33fF $ **FLOATING
C3346 sky130_asc_pfet_01v8_lvt_60_0/GATE.n359 VSS 0.05fF $ **FLOATING
C3347 sky130_asc_pfet_01v8_lvt_60_0/GATE.n360 VSS 0.08fF $ **FLOATING
C3348 sky130_asc_pfet_01v8_lvt_60_0/GATE.n361 VSS 0.05fF $ **FLOATING
C3349 sky130_asc_pfet_01v8_lvt_60_0/GATE.n362 VSS 0.08fF $ **FLOATING
C3350 sky130_asc_pfet_01v8_lvt_60_0/GATE.t120 VSS 1.44fF
C3351 sky130_asc_pfet_01v8_lvt_60_0/GATE.n363 VSS 0.33fF $ **FLOATING
C3352 sky130_asc_pfet_01v8_lvt_60_0/GATE.n364 VSS 0.05fF $ **FLOATING
C3353 sky130_asc_pfet_01v8_lvt_60_0/GATE.n365 VSS 0.08fF $ **FLOATING
C3354 sky130_asc_pfet_01v8_lvt_60_0/GATE.t99 VSS 1.44fF
C3355 sky130_asc_pfet_01v8_lvt_60_0/GATE.n366 VSS 0.33fF $ **FLOATING
C3356 sky130_asc_pfet_01v8_lvt_60_0/GATE.n367 VSS 0.05fF $ **FLOATING
C3357 sky130_asc_pfet_01v8_lvt_60_0/GATE.n368 VSS 0.08fF $ **FLOATING
C3358 sky130_asc_pfet_01v8_lvt_60_0/GATE.t182 VSS 1.44fF
C3359 sky130_asc_pfet_01v8_lvt_60_0/GATE.n369 VSS 0.33fF $ **FLOATING
C3360 sky130_asc_pfet_01v8_lvt_60_0/GATE.n370 VSS 0.05fF $ **FLOATING
C3361 sky130_asc_pfet_01v8_lvt_60_0/GATE.n371 VSS 0.08fF $ **FLOATING
C3362 sky130_asc_pfet_01v8_lvt_60_0/GATE.t145 VSS 1.44fF
C3363 sky130_asc_pfet_01v8_lvt_60_0/GATE.n372 VSS 0.33fF $ **FLOATING
C3364 sky130_asc_pfet_01v8_lvt_60_0/GATE.n373 VSS 0.05fF $ **FLOATING
C3365 sky130_asc_pfet_01v8_lvt_60_0/GATE.n374 VSS 0.08fF $ **FLOATING
C3366 sky130_asc_pfet_01v8_lvt_60_0/GATE.t144 VSS 1.44fF
C3367 sky130_asc_pfet_01v8_lvt_60_0/GATE.n375 VSS 0.38fF $ **FLOATING
C3368 sky130_asc_pfet_01v8_lvt_60_0/GATE.n376 VSS 0.08fF $ **FLOATING
C3369 sky130_asc_pfet_01v8_lvt_60_0/GATE.t138 VSS 1.44fF
C3370 sky130_asc_pfet_01v8_lvt_60_0/GATE.n377 VSS 0.39fF $ **FLOATING
C3371 sky130_asc_pfet_01v8_lvt_60_0/GATE.n378 VSS 0.08fF $ **FLOATING
C3372 sky130_asc_pfet_01v8_lvt_60_0/GATE.t111 VSS 1.44fF
C3373 sky130_asc_pfet_01v8_lvt_60_0/GATE.n379 VSS 0.33fF $ **FLOATING
C3374 sky130_asc_pfet_01v8_lvt_60_0/GATE.n380 VSS 0.05fF $ **FLOATING
C3375 sky130_asc_pfet_01v8_lvt_60_0/GATE.n381 VSS 0.08fF $ **FLOATING
C3376 sky130_asc_pfet_01v8_lvt_60_0/GATE.n382 VSS 0.05fF $ **FLOATING
C3377 sky130_asc_pfet_01v8_lvt_60_0/GATE.n383 VSS 0.08fF $ **FLOATING
C3378 sky130_asc_pfet_01v8_lvt_60_0/GATE.t209 VSS 1.44fF
C3379 sky130_asc_pfet_01v8_lvt_60_0/GATE.n384 VSS 0.33fF $ **FLOATING
C3380 sky130_asc_pfet_01v8_lvt_60_0/GATE.n385 VSS 0.05fF $ **FLOATING
C3381 sky130_asc_pfet_01v8_lvt_60_0/GATE.n386 VSS 0.08fF $ **FLOATING
C3382 sky130_asc_pfet_01v8_lvt_60_0/GATE.t170 VSS 1.44fF
C3383 sky130_asc_pfet_01v8_lvt_60_0/GATE.n387 VSS 0.33fF $ **FLOATING
C3384 sky130_asc_pfet_01v8_lvt_60_0/GATE.n388 VSS 0.05fF $ **FLOATING
C3385 sky130_asc_pfet_01v8_lvt_60_0/GATE.n389 VSS 0.08fF $ **FLOATING
C3386 sky130_asc_pfet_01v8_lvt_60_0/GATE.t169 VSS 1.44fF
C3387 sky130_asc_pfet_01v8_lvt_60_0/GATE.n390 VSS 0.33fF $ **FLOATING
C3388 sky130_asc_pfet_01v8_lvt_60_0/GATE.n391 VSS 0.05fF $ **FLOATING
C3389 sky130_asc_pfet_01v8_lvt_60_0/GATE.n392 VSS 0.08fF $ **FLOATING
C3390 sky130_asc_pfet_01v8_lvt_60_0/GATE.t160 VSS 1.44fF
C3391 sky130_asc_pfet_01v8_lvt_60_0/GATE.n393 VSS 0.38fF $ **FLOATING
C3392 sky130_asc_pfet_01v8_lvt_60_0/GATE.n394 VSS 0.07fF $ **FLOATING
C3393 sky130_asc_pfet_01v8_lvt_60_0/GATE.n395 VSS 0.09fF $ **FLOATING
C3394 sky130_asc_pfet_01v8_lvt_60_0/GATE.t132 VSS 1.44fF
C3395 sky130_asc_pfet_01v8_lvt_60_0/GATE.n396 VSS 0.37fF $ **FLOATING
C3396 sky130_asc_pfet_01v8_lvt_60_0/GATE.n397 VSS 0.05fF $ **FLOATING
C3397 sky130_asc_pfet_01v8_lvt_60_0/GATE.n398 VSS 0.08fF $ **FLOATING
C3398 sky130_asc_pfet_01v8_lvt_60_0/GATE.t131 VSS 1.44fF
C3399 sky130_asc_pfet_01v8_lvt_60_0/GATE.n399 VSS 0.33fF $ **FLOATING
C3400 sky130_asc_pfet_01v8_lvt_60_0/GATE.n400 VSS 0.05fF $ **FLOATING
C3401 sky130_asc_pfet_01v8_lvt_60_0/GATE.n401 VSS 0.08fF $ **FLOATING
C3402 sky130_asc_pfet_01v8_lvt_60_0/GATE.t201 VSS 1.44fF
C3403 sky130_asc_pfet_01v8_lvt_60_0/GATE.n402 VSS 0.33fF $ **FLOATING
C3404 sky130_asc_pfet_01v8_lvt_60_0/GATE.n403 VSS 0.05fF $ **FLOATING
C3405 sky130_asc_pfet_01v8_lvt_60_0/GATE.n404 VSS 0.08fF $ **FLOATING
C3406 sky130_asc_pfet_01v8_lvt_60_0/GATE.t124 VSS 1.44fF
C3407 sky130_asc_pfet_01v8_lvt_60_0/GATE.n405 VSS 0.38fF $ **FLOATING
C3408 sky130_asc_pfet_01v8_lvt_60_0/GATE.n406 VSS 0.08fF $ **FLOATING
C3409 sky130_asc_pfet_01v8_lvt_60_0/GATE.t191 VSS 1.44fF
C3410 sky130_asc_pfet_01v8_lvt_60_0/GATE.n407 VSS 0.39fF $ **FLOATING
C3411 sky130_asc_pfet_01v8_lvt_60_0/GATE.n408 VSS 0.08fF $ **FLOATING
C3412 sky130_asc_pfet_01v8_lvt_60_0/GATE.t90 VSS 1.44fF
C3413 sky130_asc_pfet_01v8_lvt_60_0/GATE.n409 VSS 0.33fF $ **FLOATING
C3414 sky130_asc_pfet_01v8_lvt_60_0/GATE.n410 VSS 0.05fF $ **FLOATING
C3415 sky130_asc_pfet_01v8_lvt_60_0/GATE.n411 VSS 0.08fF $ **FLOATING
C3416 sky130_asc_pfet_01v8_lvt_60_0/GATE.n412 VSS 0.05fF $ **FLOATING
C3417 sky130_asc_pfet_01v8_lvt_60_0/GATE.n413 VSS 0.08fF $ **FLOATING
C3418 sky130_asc_pfet_01v8_lvt_60_0/GATE.t66 VSS 1.44fF
C3419 sky130_asc_pfet_01v8_lvt_60_0/GATE.n414 VSS 0.33fF $ **FLOATING
C3420 sky130_asc_pfet_01v8_lvt_60_0/GATE.n415 VSS 0.05fF $ **FLOATING
C3421 sky130_asc_pfet_01v8_lvt_60_0/GATE.n416 VSS 0.08fF $ **FLOATING
C3422 sky130_asc_pfet_01v8_lvt_60_0/GATE.t128 VSS 1.44fF
C3423 sky130_asc_pfet_01v8_lvt_60_0/GATE.n417 VSS 0.33fF $ **FLOATING
C3424 sky130_asc_pfet_01v8_lvt_60_0/GATE.n418 VSS 0.05fF $ **FLOATING
C3425 sky130_asc_pfet_01v8_lvt_60_0/GATE.n419 VSS 0.08fF $ **FLOATING
C3426 sky130_asc_pfet_01v8_lvt_60_0/GATE.t62 VSS 1.44fF
C3427 sky130_asc_pfet_01v8_lvt_60_0/GATE.n420 VSS 0.33fF $ **FLOATING
C3428 sky130_asc_pfet_01v8_lvt_60_0/GATE.n421 VSS 0.05fF $ **FLOATING
C3429 sky130_asc_pfet_01v8_lvt_60_0/GATE.n422 VSS 0.08fF $ **FLOATING
C3430 sky130_asc_pfet_01v8_lvt_60_0/GATE.t101 VSS 1.44fF
C3431 sky130_asc_pfet_01v8_lvt_60_0/GATE.n423 VSS 0.33fF $ **FLOATING
C3432 sky130_asc_pfet_01v8_lvt_60_0/GATE.n424 VSS 0.05fF $ **FLOATING
C3433 sky130_asc_pfet_01v8_lvt_60_0/GATE.n425 VSS 0.08fF $ **FLOATING
C3434 sky130_asc_pfet_01v8_lvt_60_0/GATE.t100 VSS 1.44fF
C3435 sky130_asc_pfet_01v8_lvt_60_0/GATE.n426 VSS 0.38fF $ **FLOATING
C3436 sky130_asc_pfet_01v8_lvt_60_0/GATE.n427 VSS 0.08fF $ **FLOATING
C3437 sky130_asc_pfet_01v8_lvt_60_0/GATE.t149 VSS 1.44fF
C3438 sky130_asc_pfet_01v8_lvt_60_0/GATE.n428 VSS 0.39fF $ **FLOATING
C3439 sky130_asc_pfet_01v8_lvt_60_0/GATE.n429 VSS 0.08fF $ **FLOATING
C3440 sky130_asc_pfet_01v8_lvt_60_0/GATE.t148 VSS 1.44fF
C3441 sky130_asc_pfet_01v8_lvt_60_0/GATE.n430 VSS 0.33fF $ **FLOATING
C3442 sky130_asc_pfet_01v8_lvt_60_0/GATE.n431 VSS 0.05fF $ **FLOATING
C3443 sky130_asc_pfet_01v8_lvt_60_0/GATE.n432 VSS 0.08fF $ **FLOATING
C3444 sky130_asc_pfet_01v8_lvt_60_0/GATE.n433 VSS 0.05fF $ **FLOATING
C3445 sky130_asc_pfet_01v8_lvt_60_0/GATE.n434 VSS 0.08fF $ **FLOATING
C3446 sky130_asc_pfet_01v8_lvt_60_0/GATE.t76 VSS 1.44fF
C3447 sky130_asc_pfet_01v8_lvt_60_0/GATE.n435 VSS 0.33fF $ **FLOATING
C3448 sky130_asc_pfet_01v8_lvt_60_0/GATE.n436 VSS 0.05fF $ **FLOATING
C3449 sky130_asc_pfet_01v8_lvt_60_0/GATE.n437 VSS 0.08fF $ **FLOATING
C3450 sky130_asc_pfet_01v8_lvt_60_0/GATE.t139 VSS 1.44fF
C3451 sky130_asc_pfet_01v8_lvt_60_0/GATE.n438 VSS 0.33fF $ **FLOATING
C3452 sky130_asc_pfet_01v8_lvt_60_0/GATE.n439 VSS 0.05fF $ **FLOATING
C3453 sky130_asc_pfet_01v8_lvt_60_0/GATE.n440 VSS 0.08fF $ **FLOATING
C3454 sky130_asc_pfet_01v8_lvt_60_0/GATE.t112 VSS 1.44fF
C3455 sky130_asc_pfet_01v8_lvt_60_0/GATE.n441 VSS 0.33fF $ **FLOATING
C3456 sky130_asc_pfet_01v8_lvt_60_0/GATE.n442 VSS 0.05fF $ **FLOATING
C3457 sky130_asc_pfet_01v8_lvt_60_0/GATE.n443 VSS 0.08fF $ **FLOATING
C3458 sky130_asc_pfet_01v8_lvt_60_0/GATE.t210 VSS 1.44fF
C3459 sky130_asc_pfet_01v8_lvt_60_0/GATE.n444 VSS 0.33fF $ **FLOATING
C3460 sky130_asc_pfet_01v8_lvt_60_0/GATE.n445 VSS 0.05fF $ **FLOATING
C3461 sky130_asc_pfet_01v8_lvt_60_0/GATE.n446 VSS 0.08fF $ **FLOATING
C3462 sky130_asc_pfet_01v8_lvt_60_0/GATE.t172 VSS 1.44fF
C3463 sky130_asc_pfet_01v8_lvt_60_0/GATE.n447 VSS 0.38fF $ **FLOATING
C3464 sky130_asc_pfet_01v8_lvt_60_0/GATE.n448 VSS 0.08fF $ **FLOATING
C3465 sky130_asc_pfet_01v8_lvt_60_0/GATE.t199 VSS 1.44fF
C3466 sky130_asc_pfet_01v8_lvt_60_0/GATE.n449 VSS 0.39fF $ **FLOATING
C3467 sky130_asc_pfet_01v8_lvt_60_0/GATE.n450 VSS 0.08fF $ **FLOATING
C3468 sky130_asc_pfet_01v8_lvt_60_0/GATE.t161 VSS 1.44fF
C3469 sky130_asc_pfet_01v8_lvt_60_0/GATE.n451 VSS 0.38fF $ **FLOATING
C3470 sky130_asc_pfet_01v8_lvt_60_0/GATE.n452 VSS 0.08fF $ **FLOATING
C3471 sky130_asc_pfet_01v8_lvt_60_0/GATE.n453 VSS 0.05fF $ **FLOATING
C3472 sky130_asc_pfet_01v8_lvt_60_0/GATE.n454 VSS 0.08fF $ **FLOATING
C3473 sky130_asc_pfet_01v8_lvt_60_0/GATE.t159 VSS 1.44fF
C3474 sky130_asc_pfet_01v8_lvt_60_0/GATE.n455 VSS 0.33fF $ **FLOATING
C3475 sky130_asc_pfet_01v8_lvt_60_0/GATE.n456 VSS 0.05fF $ **FLOATING
C3476 sky130_asc_pfet_01v8_lvt_60_0/GATE.n457 VSS 0.08fF $ **FLOATING
C3477 sky130_asc_pfet_01v8_lvt_60_0/GATE.t223 VSS 1.44fF
C3478 sky130_asc_pfet_01v8_lvt_60_0/GATE.n458 VSS 0.33fF $ **FLOATING
C3479 sky130_asc_pfet_01v8_lvt_60_0/GATE.n459 VSS 0.05fF $ **FLOATING
C3480 sky130_asc_pfet_01v8_lvt_60_0/GATE.n460 VSS 0.08fF $ **FLOATING
C3481 sky130_asc_pfet_01v8_lvt_60_0/GATE.t195 VSS 1.44fF
C3482 sky130_asc_pfet_01v8_lvt_60_0/GATE.n461 VSS 0.33fF $ **FLOATING
C3483 sky130_asc_pfet_01v8_lvt_60_0/GATE.n462 VSS 0.05fF $ **FLOATING
C3484 sky130_asc_pfet_01v8_lvt_60_0/GATE.n463 VSS 0.08fF $ **FLOATING
C3485 sky130_asc_pfet_01v8_lvt_60_0/GATE.t218 VSS 1.44fF
C3486 sky130_asc_pfet_01v8_lvt_60_0/GATE.n464 VSS 0.33fF $ **FLOATING
C3487 sky130_asc_pfet_01v8_lvt_60_0/GATE.n465 VSS 0.05fF $ **FLOATING
C3488 sky130_asc_pfet_01v8_lvt_60_0/GATE.n466 VSS 0.08fF $ **FLOATING
C3489 sky130_asc_pfet_01v8_lvt_60_0/GATE.t185 VSS 1.44fF
C3490 sky130_asc_pfet_01v8_lvt_60_0/GATE.n467 VSS 0.38fF $ **FLOATING
C3491 sky130_asc_pfet_01v8_lvt_60_0/GATE.n468 VSS 0.08fF $ **FLOATING
C3492 sky130_asc_pfet_01v8_lvt_60_0/GATE.t184 VSS 1.44fF
C3493 sky130_asc_pfet_01v8_lvt_60_0/GATE.n469 VSS 0.39fF $ **FLOATING
C3494 sky130_asc_pfet_01v8_lvt_60_0/GATE.n470 VSS 0.08fF $ **FLOATING
C3495 sky130_asc_pfet_01v8_lvt_60_0/GATE.t237 VSS 1.44fF
C3496 sky130_asc_pfet_01v8_lvt_60_0/GATE.n471 VSS 0.38fF $ **FLOATING
C3497 sky130_asc_pfet_01v8_lvt_60_0/GATE.n472 VSS 0.08fF $ **FLOATING
C3498 sky130_asc_pfet_01v8_lvt_60_0/GATE.t123 VSS 1.44fF
C3499 sky130_asc_pfet_01v8_lvt_60_0/GATE.n473 VSS 0.33fF $ **FLOATING
C3500 sky130_asc_pfet_01v8_lvt_60_0/GATE.n474 VSS 0.05fF $ **FLOATING
C3501 sky130_asc_pfet_01v8_lvt_60_0/GATE.n475 VSS 0.08fF $ **FLOATING
C3502 sky130_asc_pfet_01v8_lvt_60_0/GATE.n476 VSS 0.05fF $ **FLOATING
C3503 sky130_asc_pfet_01v8_lvt_60_0/GATE.n477 VSS 0.08fF $ **FLOATING
C3504 sky130_asc_pfet_01v8_lvt_60_0/GATE.t119 VSS 1.44fF
C3505 sky130_asc_pfet_01v8_lvt_60_0/GATE.n478 VSS 0.33fF $ **FLOATING
C3506 sky130_asc_pfet_01v8_lvt_60_0/GATE.n479 VSS 0.05fF $ **FLOATING
C3507 sky130_asc_pfet_01v8_lvt_60_0/GATE.n480 VSS 0.08fF $ **FLOATING
C3508 sky130_asc_pfet_01v8_lvt_60_0/GATE.t117 VSS 1.44fF
C3509 sky130_asc_pfet_01v8_lvt_60_0/GATE.n481 VSS 0.33fF $ **FLOATING
C3510 sky130_asc_pfet_01v8_lvt_60_0/GATE.n482 VSS 0.05fF $ **FLOATING
C3511 sky130_asc_pfet_01v8_lvt_60_0/GATE.n483 VSS 0.08fF $ **FLOATING
C3512 sky130_asc_pfet_01v8_lvt_60_0/GATE.t180 VSS 1.44fF
C3513 sky130_asc_pfet_01v8_lvt_60_0/GATE.n484 VSS 0.33fF $ **FLOATING
C3514 sky130_asc_pfet_01v8_lvt_60_0/GATE.n485 VSS 0.05fF $ **FLOATING
C3515 sky130_asc_pfet_01v8_lvt_60_0/GATE.n486 VSS 0.08fF $ **FLOATING
C3516 sky130_asc_pfet_01v8_lvt_60_0/GATE.t179 VSS 1.44fF
C3517 sky130_asc_pfet_01v8_lvt_60_0/GATE.n487 VSS 0.33fF $ **FLOATING
C3518 sky130_asc_pfet_01v8_lvt_60_0/GATE.n488 VSS 0.05fF $ **FLOATING
C3519 sky130_asc_pfet_01v8_lvt_60_0/GATE.n489 VSS 0.07fF $ **FLOATING
C3520 sky130_asc_pfet_01v8_lvt_60_0/GATE.n490 VSS 0.04fF $ **FLOATING
C3521 sky130_asc_pfet_01v8_lvt_60_0/GATE.t181 VSS 2.37fF
C3522 sky130_asc_pfet_01v8_lvt_60_0/GATE.n491 VSS 0.07fF $ **FLOATING
C3523 sky130_asc_pfet_01v8_lvt_60_0/GATE.t142 VSS 1.44fF
C3524 sky130_asc_pfet_01v8_lvt_60_0/GATE.n492 VSS 0.27fF $ **FLOATING
C3525 sky130_asc_pfet_01v8_lvt_60_0/GATE.n493 VSS 0.11fF $ **FLOATING
C3526 sky130_asc_pfet_01v8_lvt_60_0/GATE.n494 VSS 0.02fF $ **FLOATING
C3527 sky130_asc_pfet_01v8_lvt_60_0/GATE.n495 VSS 0.00fF $ **FLOATING
C3528 sky130_asc_pfet_01v8_lvt_60_0/GATE.n496 VSS 0.00fF $ **FLOATING
C3529 sky130_asc_pfet_01v8_lvt_60_0/GATE.n497 VSS 0.04fF $ **FLOATING
C3530 sky130_asc_pfet_01v8_lvt_60_0/GATE.t135 VSS 1.44fF
C3531 sky130_asc_pfet_01v8_lvt_60_0/GATE.n498 VSS 0.38fF $ **FLOATING
C3532 sky130_asc_pfet_01v8_lvt_60_0/GATE.n499 VSS 0.08fF $ **FLOATING
C3533 sky130_asc_pfet_01v8_lvt_60_0/GATE.t133 VSS 1.44fF
C3534 sky130_asc_pfet_01v8_lvt_60_0/GATE.n500 VSS 0.33fF $ **FLOATING
C3535 sky130_asc_pfet_01v8_lvt_60_0/GATE.n501 VSS 0.05fF $ **FLOATING
C3536 sky130_asc_pfet_01v8_lvt_60_0/GATE.n502 VSS 0.08fF $ **FLOATING
C3537 sky130_asc_pfet_01v8_lvt_60_0/GATE.n503 VSS 0.05fF $ **FLOATING
C3538 sky130_asc_pfet_01v8_lvt_60_0/GATE.n504 VSS 0.08fF $ **FLOATING
C3539 sky130_asc_pfet_01v8_lvt_60_0/GATE.t206 VSS 1.44fF
C3540 sky130_asc_pfet_01v8_lvt_60_0/GATE.n505 VSS 0.33fF $ **FLOATING
C3541 sky130_asc_pfet_01v8_lvt_60_0/GATE.n506 VSS 0.05fF $ **FLOATING
C3542 sky130_asc_pfet_01v8_lvt_60_0/GATE.n507 VSS 0.08fF $ **FLOATING
C3543 sky130_asc_pfet_01v8_lvt_60_0/GATE.t204 VSS 1.44fF
C3544 sky130_asc_pfet_01v8_lvt_60_0/GATE.n508 VSS 0.33fF $ **FLOATING
C3545 sky130_asc_pfet_01v8_lvt_60_0/GATE.n509 VSS 0.05fF $ **FLOATING
C3546 sky130_asc_pfet_01v8_lvt_60_0/GATE.n510 VSS 0.08fF $ **FLOATING
C3547 sky130_asc_pfet_01v8_lvt_60_0/GATE.t168 VSS 1.44fF
C3548 sky130_asc_pfet_01v8_lvt_60_0/GATE.n511 VSS 0.33fF $ **FLOATING
C3549 sky130_asc_pfet_01v8_lvt_60_0/GATE.n512 VSS 0.05fF $ **FLOATING
C3550 sky130_asc_pfet_01v8_lvt_60_0/GATE.n513 VSS 0.08fF $ **FLOATING
C3551 sky130_asc_pfet_01v8_lvt_60_0/GATE.t192 VSS 1.44fF
C3552 sky130_asc_pfet_01v8_lvt_60_0/GATE.n514 VSS 0.33fF $ **FLOATING
C3553 sky130_asc_pfet_01v8_lvt_60_0/GATE.n515 VSS 0.05fF $ **FLOATING
C3554 sky130_asc_pfet_01v8_lvt_60_0/GATE.n516 VSS 0.08fF $ **FLOATING
C3555 sky130_asc_pfet_01v8_lvt_60_0/GATE.t154 VSS 1.44fF
C3556 sky130_asc_pfet_01v8_lvt_60_0/GATE.n517 VSS 0.39fF $ **FLOATING
C3557 sky130_asc_pfet_01v8_lvt_60_0/GATE.n518 VSS 0.08fF $ **FLOATING
C3558 sky130_asc_pfet_01v8_lvt_60_0/GATE.t242 VSS 1.44fF
C3559 sky130_asc_pfet_01v8_lvt_60_0/GATE.n519 VSS 0.38fF $ **FLOATING
C3560 sky130_asc_pfet_01v8_lvt_60_0/GATE.n520 VSS 0.08fF $ **FLOATING
C3561 sky130_asc_pfet_01v8_lvt_60_0/GATE.t221 VSS 1.44fF
C3562 sky130_asc_pfet_01v8_lvt_60_0/GATE.n521 VSS 0.33fF $ **FLOATING
C3563 sky130_asc_pfet_01v8_lvt_60_0/GATE.n522 VSS 0.05fF $ **FLOATING
C3564 sky130_asc_pfet_01v8_lvt_60_0/GATE.n523 VSS 0.08fF $ **FLOATING
C3565 sky130_asc_pfet_01v8_lvt_60_0/GATE.n524 VSS 0.05fF $ **FLOATING
C3566 sky130_asc_pfet_01v8_lvt_60_0/GATE.n525 VSS 0.08fF $ **FLOATING
C3567 sky130_asc_pfet_01v8_lvt_60_0/GATE.t65 VSS 1.44fF
C3568 sky130_asc_pfet_01v8_lvt_60_0/GATE.n526 VSS 0.33fF $ **FLOATING
C3569 sky130_asc_pfet_01v8_lvt_60_0/GATE.n527 VSS 0.05fF $ **FLOATING
C3570 sky130_asc_pfet_01v8_lvt_60_0/GATE.n528 VSS 0.08fF $ **FLOATING
C3571 sky130_asc_pfet_01v8_lvt_60_0/GATE.t215 VSS 1.44fF
C3572 sky130_asc_pfet_01v8_lvt_60_0/GATE.n529 VSS 0.33fF $ **FLOATING
C3573 sky130_asc_pfet_01v8_lvt_60_0/GATE.n530 VSS 0.05fF $ **FLOATING
C3574 sky130_asc_pfet_01v8_lvt_60_0/GATE.n531 VSS 0.08fF $ **FLOATING
C3575 sky130_asc_pfet_01v8_lvt_60_0/GATE.t214 VSS 1.44fF
C3576 sky130_asc_pfet_01v8_lvt_60_0/GATE.n532 VSS 0.33fF $ **FLOATING
C3577 sky130_asc_pfet_01v8_lvt_60_0/GATE.n533 VSS 0.05fF $ **FLOATING
C3578 sky130_asc_pfet_01v8_lvt_60_0/GATE.n534 VSS 0.08fF $ **FLOATING
C3579 sky130_asc_pfet_01v8_lvt_60_0/GATE.t39 VSS 1.44fF
C3580 sky130_asc_pfet_01v8_lvt_60_0/GATE.n535 VSS 0.33fF $ **FLOATING
C3581 sky130_asc_pfet_01v8_lvt_60_0/GATE.n536 VSS 0.05fF $ **FLOATING
C3582 sky130_asc_pfet_01v8_lvt_60_0/GATE.n537 VSS 0.08fF $ **FLOATING
C3583 sky130_asc_pfet_01v8_lvt_60_0/GATE.t236 VSS 1.44fF
C3584 sky130_asc_pfet_01v8_lvt_60_0/GATE.n538 VSS 0.38fF $ **FLOATING
C3585 sky130_asc_pfet_01v8_lvt_60_0/GATE.n539 VSS 0.08fF $ **FLOATING
C3586 sky130_asc_pfet_01v8_lvt_60_0/GATE.t83 VSS 1.44fF
C3587 sky130_asc_pfet_01v8_lvt_60_0/GATE.n540 VSS 0.38fF $ **FLOATING
C3588 sky130_asc_pfet_01v8_lvt_60_0/GATE.n541 VSS 0.08fF $ **FLOATING
C3589 sky130_asc_pfet_01v8_lvt_60_0/GATE.t229 VSS 1.44fF
C3590 sky130_asc_pfet_01v8_lvt_60_0/GATE.n542 VSS 0.33fF $ **FLOATING
C3591 sky130_asc_pfet_01v8_lvt_60_0/GATE.n543 VSS 0.05fF $ **FLOATING
C3592 sky130_asc_pfet_01v8_lvt_60_0/GATE.n544 VSS 0.08fF $ **FLOATING
C3593 sky130_asc_pfet_01v8_lvt_60_0/GATE.n545 VSS 0.05fF $ **FLOATING
C3594 sky130_asc_pfet_01v8_lvt_60_0/GATE.n546 VSS 0.08fF $ **FLOATING
C3595 sky130_asc_pfet_01v8_lvt_60_0/GATE.t212 VSS 1.44fF
C3596 sky130_asc_pfet_01v8_lvt_60_0/GATE.n547 VSS 0.33fF $ **FLOATING
C3597 sky130_asc_pfet_01v8_lvt_60_0/GATE.n548 VSS 0.05fF $ **FLOATING
C3598 sky130_asc_pfet_01v8_lvt_60_0/GATE.n549 VSS 0.08fF $ **FLOATING
C3599 sky130_asc_pfet_01v8_lvt_60_0/GATE.t176 VSS 1.44fF
C3600 sky130_asc_pfet_01v8_lvt_60_0/GATE.n550 VSS 0.33fF $ **FLOATING
C3601 sky130_asc_pfet_01v8_lvt_60_0/GATE.n551 VSS 0.05fF $ **FLOATING
C3602 sky130_asc_pfet_01v8_lvt_60_0/GATE.n552 VSS 0.08fF $ **FLOATING
C3603 sky130_asc_pfet_01v8_lvt_60_0/GATE.t174 VSS 1.44fF
C3604 sky130_asc_pfet_01v8_lvt_60_0/GATE.n553 VSS 0.33fF $ **FLOATING
C3605 sky130_asc_pfet_01v8_lvt_60_0/GATE.n554 VSS 0.05fF $ **FLOATING
C3606 sky130_asc_pfet_01v8_lvt_60_0/GATE.n555 VSS 0.08fF $ **FLOATING
C3607 sky130_asc_pfet_01v8_lvt_60_0/GATE.t232 VSS 1.44fF
C3608 sky130_asc_pfet_01v8_lvt_60_0/GATE.n556 VSS 0.33fF $ **FLOATING
C3609 sky130_asc_pfet_01v8_lvt_60_0/GATE.n557 VSS 0.05fF $ **FLOATING
C3610 sky130_asc_pfet_01v8_lvt_60_0/GATE.n558 VSS 0.08fF $ **FLOATING
C3611 sky130_asc_pfet_01v8_lvt_60_0/GATE.t163 VSS 1.44fF
C3612 sky130_asc_pfet_01v8_lvt_60_0/GATE.n559 VSS 0.38fF $ **FLOATING
C3613 sky130_asc_pfet_01v8_lvt_60_0/GATE.n560 VSS 0.08fF $ **FLOATING
C3614 sky130_asc_pfet_01v8_lvt_60_0/GATE.t227 VSS 1.44fF
C3615 sky130_asc_pfet_01v8_lvt_60_0/GATE.n561 VSS 0.39fF $ **FLOATING
C3616 sky130_asc_pfet_01v8_lvt_60_0/GATE.n562 VSS 0.08fF $ **FLOATING
C3617 sky130_asc_pfet_01v8_lvt_60_0/GATE.t224 VSS 1.44fF
C3618 sky130_asc_pfet_01v8_lvt_60_0/GATE.n563 VSS 0.33fF $ **FLOATING
C3619 sky130_asc_pfet_01v8_lvt_60_0/GATE.n564 VSS 0.05fF $ **FLOATING
C3620 sky130_asc_pfet_01v8_lvt_60_0/GATE.n565 VSS 0.08fF $ **FLOATING
C3621 sky130_asc_pfet_01v8_lvt_60_0/GATE.n566 VSS 0.05fF $ **FLOATING
C3622 sky130_asc_pfet_01v8_lvt_60_0/GATE.n567 VSS 0.08fF $ **FLOATING
C3623 sky130_asc_pfet_01v8_lvt_60_0/GATE.t197 VSS 1.44fF
C3624 sky130_asc_pfet_01v8_lvt_60_0/GATE.n568 VSS 0.33fF $ **FLOATING
C3625 sky130_asc_pfet_01v8_lvt_60_0/GATE.n569 VSS 0.05fF $ **FLOATING
C3626 sky130_asc_pfet_01v8_lvt_60_0/GATE.n570 VSS 0.08fF $ **FLOATING
C3627 sky130_asc_pfet_01v8_lvt_60_0/GATE.t25 VSS 1.44fF
C3628 sky130_asc_pfet_01v8_lvt_60_0/GATE.n571 VSS 0.33fF $ **FLOATING
C3629 sky130_asc_pfet_01v8_lvt_60_0/GATE.n572 VSS 0.05fF $ **FLOATING
C3630 sky130_asc_pfet_01v8_lvt_60_0/GATE.n573 VSS 0.08fF $ **FLOATING
C3631 sky130_asc_pfet_01v8_lvt_60_0/GATE.t186 VSS 1.44fF
C3632 sky130_asc_pfet_01v8_lvt_60_0/GATE.n574 VSS 0.33fF $ **FLOATING
C3633 sky130_asc_pfet_01v8_lvt_60_0/GATE.n575 VSS 0.05fF $ **FLOATING
C3634 sky130_asc_pfet_01v8_lvt_60_0/GATE.n576 VSS 0.08fF $ **FLOATING
C3635 sky130_asc_pfet_01v8_lvt_60_0/GATE.t239 VSS 1.44fF
C3636 sky130_asc_pfet_01v8_lvt_60_0/GATE.n577 VSS 0.38fF $ **FLOATING
C3637 sky130_asc_pfet_01v8_lvt_60_0/GATE.n578 VSS 0.09fF $ **FLOATING
C3638 sky130_asc_pfet_01v8_lvt_60_0/GATE.t92 VSS 1.93fF
C3639 sky130_asc_pfet_01v8_lvt_60_0/GATE.n579 VSS 0.34fF $ **FLOATING
C3640 sky130_asc_pfet_01v8_lvt_60_0/GATE.t42 VSS 1.44fF
C3641 sky130_asc_pfet_01v8_lvt_60_0/GATE.n580 VSS 0.33fF $ **FLOATING
C3642 sky130_asc_pfet_01v8_lvt_60_0/GATE.n581 VSS 0.05fF $ **FLOATING
C3643 sky130_asc_pfet_01v8_lvt_60_0/GATE.t216 VSS 1.44fF
C3644 sky130_asc_pfet_01v8_lvt_60_0/GATE.n582 VSS 0.33fF $ **FLOATING
C3645 sky130_asc_pfet_01v8_lvt_60_0/GATE.n583 VSS 0.05fF $ **FLOATING
C3646 sky130_asc_pfet_01v8_lvt_60_0/GATE.n584 VSS 0.23fF $ **FLOATING
C3647 sky130_asc_pfet_01v8_lvt_60_0/GATE.t217 VSS 1.44fF
C3648 sky130_asc_pfet_01v8_lvt_60_0/GATE.n585 VSS 0.33fF $ **FLOATING
C3649 sky130_asc_pfet_01v8_lvt_60_0/GATE.n586 VSS 0.05fF $ **FLOATING
C3650 sky130_asc_pfet_01v8_lvt_60_0/GATE.n587 VSS 0.08fF $ **FLOATING
C3651 sky130_asc_pfet_01v8_lvt_60_0/GATE.n588 VSS 0.08fF $ **FLOATING
C3652 sky130_asc_pfet_01v8_lvt_60_0/GATE.n589 VSS 0.08fF $ **FLOATING
C3653 sky130_asc_pfet_01v8_lvt_60_0/GATE.t24 VSS 1.44fF
C3654 sky130_asc_pfet_01v8_lvt_60_0/GATE.n590 VSS 0.33fF $ **FLOATING
C3655 sky130_asc_pfet_01v8_lvt_60_0/GATE.n591 VSS 0.05fF $ **FLOATING
C3656 sky130_asc_pfet_01v8_lvt_60_0/GATE.n592 VSS 0.08fF $ **FLOATING
C3657 sky130_asc_pfet_01v8_lvt_60_0/GATE.n593 VSS 0.05fF $ **FLOATING
C3658 sky130_asc_pfet_01v8_lvt_60_0/GATE.n594 VSS 0.08fF $ **FLOATING
C3659 sky130_asc_pfet_01v8_lvt_60_0/GATE.t158 VSS 1.44fF
C3660 sky130_asc_pfet_01v8_lvt_60_0/GATE.n595 VSS 0.33fF $ **FLOATING
C3661 sky130_asc_pfet_01v8_lvt_60_0/GATE.n596 VSS 0.05fF $ **FLOATING
C3662 sky130_asc_pfet_01v8_lvt_60_0/GATE.n597 VSS 0.08fF $ **FLOATING
C3663 sky130_asc_pfet_01v8_lvt_60_0/GATE.t196 VSS 1.44fF
C3664 sky130_asc_pfet_01v8_lvt_60_0/GATE.n598 VSS 0.33fF $ **FLOATING
C3665 sky130_asc_pfet_01v8_lvt_60_0/GATE.n599 VSS 0.05fF $ **FLOATING
C3666 sky130_asc_pfet_01v8_lvt_60_0/GATE.n600 VSS 0.08fF $ **FLOATING
C3667 sky130_asc_pfet_01v8_lvt_60_0/GATE.t171 VSS 1.44fF
C3668 sky130_asc_pfet_01v8_lvt_60_0/GATE.n601 VSS 0.33fF $ **FLOATING
C3669 sky130_asc_pfet_01v8_lvt_60_0/GATE.n602 VSS 0.05fF $ **FLOATING
C3670 sky130_asc_pfet_01v8_lvt_60_0/GATE.n603 VSS 0.08fF $ **FLOATING
C3671 sky130_asc_pfet_01v8_lvt_60_0/GATE.t208 VSS 1.44fF
C3672 sky130_asc_pfet_01v8_lvt_60_0/GATE.n604 VSS 0.33fF $ **FLOATING
C3673 sky130_asc_pfet_01v8_lvt_60_0/GATE.n605 VSS 0.05fF $ **FLOATING
C3674 sky130_asc_pfet_01v8_lvt_60_0/GATE.n606 VSS 0.08fF $ **FLOATING
C3675 sky130_asc_pfet_01v8_lvt_60_0/GATE.n607 VSS 0.08fF $ **FLOATING
C3676 sky130_asc_pfet_01v8_lvt_60_0/GATE.n608 VSS 0.08fF $ **FLOATING
C3677 sky130_asc_pfet_01v8_lvt_60_0/GATE.t173 VSS 1.44fF
C3678 sky130_asc_pfet_01v8_lvt_60_0/GATE.n609 VSS 0.33fF $ **FLOATING
C3679 sky130_asc_pfet_01v8_lvt_60_0/GATE.n610 VSS 0.05fF $ **FLOATING
C3680 sky130_asc_pfet_01v8_lvt_60_0/GATE.n611 VSS 0.08fF $ **FLOATING
C3681 sky130_asc_pfet_01v8_lvt_60_0/GATE.n612 VSS 0.05fF $ **FLOATING
C3682 sky130_asc_pfet_01v8_lvt_60_0/GATE.n613 VSS 0.08fF $ **FLOATING
C3683 sky130_asc_pfet_01v8_lvt_60_0/GATE.t146 VSS 1.44fF
C3684 sky130_asc_pfet_01v8_lvt_60_0/GATE.n614 VSS 0.33fF $ **FLOATING
C3685 sky130_asc_pfet_01v8_lvt_60_0/GATE.n615 VSS 0.05fF $ **FLOATING
C3686 sky130_asc_pfet_01v8_lvt_60_0/GATE.n616 VSS 0.08fF $ **FLOATING
C3687 sky130_asc_pfet_01v8_lvt_60_0/GATE.t183 VSS 1.44fF
C3688 sky130_asc_pfet_01v8_lvt_60_0/GATE.n617 VSS 0.33fF $ **FLOATING
C3689 sky130_asc_pfet_01v8_lvt_60_0/GATE.n618 VSS 0.05fF $ **FLOATING
C3690 sky130_asc_pfet_01v8_lvt_60_0/GATE.n619 VSS 0.08fF $ **FLOATING
C3691 sky130_asc_pfet_01v8_lvt_60_0/GATE.t60 VSS 1.44fF
C3692 sky130_asc_pfet_01v8_lvt_60_0/GATE.n620 VSS 0.33fF $ **FLOATING
C3693 sky130_asc_pfet_01v8_lvt_60_0/GATE.n621 VSS 0.05fF $ **FLOATING
C3694 sky130_asc_pfet_01v8_lvt_60_0/GATE.n622 VSS 0.08fF $ **FLOATING
C3695 sky130_asc_pfet_01v8_lvt_60_0/GATE.t233 VSS 1.44fF
C3696 sky130_asc_pfet_01v8_lvt_60_0/GATE.n623 VSS 0.33fF $ **FLOATING
C3697 sky130_asc_pfet_01v8_lvt_60_0/GATE.n624 VSS 0.05fF $ **FLOATING
C3698 sky130_asc_pfet_01v8_lvt_60_0/GATE.n625 VSS 0.08fF $ **FLOATING
C3699 sky130_asc_pfet_01v8_lvt_60_0/GATE.n626 VSS 0.08fF $ **FLOATING
C3700 sky130_asc_pfet_01v8_lvt_60_0/GATE.n627 VSS 0.08fF $ **FLOATING
C3701 sky130_asc_pfet_01v8_lvt_60_0/GATE.n628 VSS 0.08fF $ **FLOATING
C3702 sky130_asc_pfet_01v8_lvt_60_0/GATE.n629 VSS 0.05fF $ **FLOATING
C3703 sky130_asc_pfet_01v8_lvt_60_0/GATE.n630 VSS 0.08fF $ **FLOATING
C3704 sky130_asc_pfet_01v8_lvt_60_0/GATE.n631 VSS 0.08fF $ **FLOATING
C3705 sky130_asc_pfet_01v8_lvt_60_0/GATE.t225 VSS 1.44fF
C3706 sky130_asc_pfet_01v8_lvt_60_0/GATE.n632 VSS 0.33fF $ **FLOATING
C3707 sky130_asc_pfet_01v8_lvt_60_0/GATE.n633 VSS 0.05fF $ **FLOATING
C3708 sky130_asc_pfet_01v8_lvt_60_0/GATE.t220 VSS 1.44fF
C3709 sky130_asc_pfet_01v8_lvt_60_0/GATE.n634 VSS 0.33fF $ **FLOATING
C3710 sky130_asc_pfet_01v8_lvt_60_0/GATE.t190 VSS 1.44fF
C3711 sky130_asc_pfet_01v8_lvt_60_0/GATE.t188 VSS 1.44fF
C3712 sky130_asc_pfet_01v8_lvt_60_0/GATE.n635 VSS 0.33fF $ **FLOATING
C3713 sky130_asc_pfet_01v8_lvt_60_0/GATE.n636 VSS 0.05fF $ **FLOATING
C3714 sky130_asc_pfet_01v8_lvt_60_0/GATE.n637 VSS 0.33fF $ **FLOATING
C3715 sky130_asc_pfet_01v8_lvt_60_0/GATE.n638 VSS 0.05fF $ **FLOATING
C3716 sky130_asc_pfet_01v8_lvt_60_0/GATE.n639 VSS 0.21fF $ **FLOATING
C3717 sky130_asc_pfet_01v8_lvt_60_0/GATE.n640 VSS 0.67fF $ **FLOATING
C3718 sky130_asc_pfet_01v8_lvt_60_0/GATE.t6 VSS 0.52fF
C3719 sky130_asc_pfet_01v8_lvt_60_0/GATE.n641 VSS 0.42fF $ **FLOATING
C3720 sky130_asc_pfet_01v8_lvt_60_0/GATE.n642 VSS 0.18fF $ **FLOATING
C3721 sky130_asc_pfet_01v8_lvt_60_0/GATE.n643 VSS 0.18fF $ **FLOATING
C3722 sky130_asc_pfet_01v8_lvt_60_0/GATE.n644 VSS 0.14fF $ **FLOATING
C3723 sky130_asc_pfet_01v8_lvt_6_0/DRAIN VSS 0.01fF $ **FLOATING
.ends

